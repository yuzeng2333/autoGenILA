module word_adder(clk, func, inWord, rst, clk, func, inWord, rst);
  input [0:0] clk;
  input [1:0] func;
  input [8:0] inWord;
  input [0:0] rst;
  output [8:0] result;
  reg [8:0] word;
endmodule
