module bar__DOT__i1(
__START__,
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
key,
state_in,
state_out,
__COUNTER_start__n0
);
input            __START__;
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg    [127:0] key;
output reg    [127:0] state_in;
output reg    [127:0] state_out;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire            __START__;
wire    [127:0] bv_128_0_n1;
wire      [7:0] bv_8_0_n580;
wire      [7:0] bv_8_100_n348;
wire      [7:0] bv_8_101_n49;
wire      [7:0] bv_8_102_n527;
wire      [7:0] bv_8_103_n523;
wire      [7:0] bv_8_104_n520;
wire      [7:0] bv_8_105_n148;
wire      [7:0] bv_8_106_n155;
wire      [7:0] bv_8_107_n370;
wire      [7:0] bv_8_108_n510;
wire      [7:0] bv_8_109_n9;
wire      [7:0] bv_8_10_n655;
wire      [7:0] bv_8_110_n294;
wire      [7:0] bv_8_111_n244;
wire      [7:0] bv_8_112_n482;
wire      [7:0] bv_8_113_n180;
wire      [7:0] bv_8_114_n494;
wire      [7:0] bv_8_115_n222;
wire      [7:0] bv_8_116_n345;
wire      [7:0] bv_8_117_n484;
wire      [7:0] bv_8_118_n480;
wire      [7:0] bv_8_119_n472;
wire      [7:0] bv_8_11_n379;
wire      [7:0] bv_8_120_n474;
wire      [7:0] bv_8_121_n470;
wire      [7:0] bv_8_122_n416;
wire      [7:0] bv_8_123_n17;
wire      [7:0] bv_8_124_n184;
wire      [7:0] bv_8_125_n459;
wire      [7:0] bv_8_126_n456;
wire      [7:0] bv_8_127_n453;
wire      [7:0] bv_8_128_n450;
wire      [7:0] bv_8_129_n446;
wire      [7:0] bv_8_12_n333;
wire      [7:0] bv_8_130_n33;
wire      [7:0] bv_8_131_n440;
wire      [7:0] bv_8_132_n41;
wire      [7:0] bv_8_133_n434;
wire      [7:0] bv_8_134_n431;
wire      [7:0] bv_8_135_n81;
wire      [7:0] bv_8_136_n425;
wire      [7:0] bv_8_137_n421;
wire      [7:0] bv_8_138_n418;
wire      [7:0] bv_8_139_n297;
wire      [7:0] bv_8_13_n194;
wire      [7:0] bv_8_140_n376;
wire      [7:0] bv_8_141_n410;
wire      [7:0] bv_8_142_n406;
wire      [7:0] bv_8_143_n403;
wire      [7:0] bv_8_144_n173;
wire      [7:0] bv_8_145_n397;
wire      [7:0] bv_8_146_n337;
wire      [7:0] bv_8_147_n392;
wire      [7:0] bv_8_148_n388;
wire      [7:0] bv_8_149_n384;
wire      [7:0] bv_8_14_n648;
wire      [7:0] bv_8_150_n201;
wire      [7:0] bv_8_151_n218;
wire      [7:0] bv_8_152_n374;
wire      [7:0] bv_8_153_n140;
wire      [7:0] bv_8_154_n368;
wire      [7:0] bv_8_155_n364;
wire      [7:0] bv_8_156_n279;
wire      [7:0] bv_8_157_n359;
wire      [7:0] bv_8_158_n355;
wire      [7:0] bv_8_159_n323;
wire      [7:0] bv_8_15_n190;
wire      [7:0] bv_8_160_n350;
wire      [7:0] bv_8_161_n211;
wire      [7:0] bv_8_162_n343;
wire      [7:0] bv_8_163_n339;
wire      [7:0] bv_8_164_n335;
wire      [7:0] bv_8_165_n69;
wire      [7:0] bv_8_166_n328;
wire      [7:0] bv_8_167_n325;
wire      [7:0] bv_8_168_n13;
wire      [7:0] bv_8_169_n109;
wire      [7:0] bv_8_16_n248;
wire      [7:0] bv_8_170_n77;
wire      [7:0] bv_8_171_n314;
wire      [7:0] bv_8_172_n268;
wire      [7:0] bv_8_173_n307;
wire      [7:0] bv_8_174_n152;
wire      [7:0] bv_8_175_n302;
wire      [7:0] bv_8_176_n299;
wire      [7:0] bv_8_177_n283;
wire      [7:0] bv_8_178_n292;
wire      [7:0] bv_8_179_n289;
wire      [7:0] bv_8_17_n525;
wire      [7:0] bv_8_180_n285;
wire      [7:0] bv_8_181_n281;
wire      [7:0] bv_8_182_n277;
wire      [7:0] bv_8_183_n273;
wire      [7:0] bv_8_184_n270;
wire      [7:0] bv_8_185_n266;
wire      [7:0] bv_8_186_n263;
wire      [7:0] bv_8_187_n260;
wire      [7:0] bv_8_188_n257;
wire      [7:0] bv_8_189_n254;
wire      [7:0] bv_8_18_n628;
wire      [7:0] bv_8_190_n250;
wire      [7:0] bv_8_191_n246;
wire      [7:0] bv_8_192_n242;
wire      [7:0] bv_8_193_n239;
wire      [7:0] bv_8_194_n159;
wire      [7:0] bv_8_195_n232;
wire      [7:0] bv_8_196_n228;
wire      [7:0] bv_8_197_n224;
wire      [7:0] bv_8_198_n220;
wire      [7:0] bv_8_199_n216;
wire      [7:0] bv_8_19_n588;
wire      [7:0] bv_8_1_n287;
wire      [7:0] bv_8_200_n213;
wire      [7:0] bv_8_201_n85;
wire      [7:0] bv_8_202_n207;
wire      [7:0] bv_8_203_n203;
wire      [7:0] bv_8_204_n177;
wire      [7:0] bv_8_205_n196;
wire      [7:0] bv_8_206_n192;
wire      [7:0] bv_8_207_n188;
wire      [7:0] bv_8_208_n37;
wire      [7:0] bv_8_209_n182;
wire      [7:0] bv_8_20_n341;
wire      [7:0] bv_8_210_n113;
wire      [7:0] bv_8_211_n175;
wire      [7:0] bv_8_212_n171;
wire      [7:0] bv_8_213_n167;
wire      [7:0] bv_8_214_n164;
wire      [7:0] bv_8_215_n45;
wire      [7:0] bv_8_216_n157;
wire      [7:0] bv_8_217_n128;
wire      [7:0] bv_8_218_n150;
wire      [7:0] bv_8_219_n146;
wire      [7:0] bv_8_21_n89;
wire      [7:0] bv_8_220_n142;
wire      [7:0] bv_8_221_n138;
wire      [7:0] bv_8_222_n134;
wire      [7:0] bv_8_223_n130;
wire      [7:0] bv_8_224_n126;
wire      [7:0] bv_8_225_n123;
wire      [7:0] bv_8_226_n119;
wire      [7:0] bv_8_227_n115;
wire      [7:0] bv_8_228_n111;
wire      [7:0] bv_8_229_n107;
wire      [7:0] bv_8_22_n357;
wire      [7:0] bv_8_230_n103;
wire      [7:0] bv_8_231_n99;
wire      [7:0] bv_8_232_n95;
wire      [7:0] bv_8_233_n91;
wire      [7:0] bv_8_234_n87;
wire      [7:0] bv_8_235_n83;
wire      [7:0] bv_8_236_n79;
wire      [7:0] bv_8_237_n75;
wire      [7:0] bv_8_238_n71;
wire      [7:0] bv_8_239_n67;
wire      [7:0] bv_8_23_n144;
wire      [7:0] bv_8_240_n63;
wire      [7:0] bv_8_241_n59;
wire      [7:0] bv_8_242_n55;
wire      [7:0] bv_8_243_n51;
wire      [7:0] bv_8_244_n47;
wire      [7:0] bv_8_245_n43;
wire      [7:0] bv_8_246_n39;
wire      [7:0] bv_8_247_n35;
wire      [7:0] bv_8_248_n31;
wire      [7:0] bv_8_249_n27;
wire      [7:0] bv_8_24_n448;
wire      [7:0] bv_8_250_n23;
wire      [7:0] bv_8_251_n19;
wire      [7:0] bv_8_252_n15;
wire      [7:0] bv_8_253_n11;
wire      [7:0] bv_8_254_n7;
wire      [7:0] bv_8_255_n3;
wire      [7:0] bv_8_25_n399;
wire      [7:0] bv_8_26_n53;
wire      [7:0] bv_8_27_n642;
wire      [7:0] bv_8_28_n162;
wire      [7:0] bv_8_29_n625;
wire      [7:0] bv_8_2_n751;
wire      [7:0] bv_8_30_n21;
wire      [7:0] bv_8_31_n705;
wire      [7:0] bv_8_32_n463;
wire      [7:0] bv_8_33_n486;
wire      [7:0] bv_8_34_n117;
wire      [7:0] bv_8_35_n696;
wire      [7:0] bv_8_36_n645;
wire      [7:0] bv_8_37_n506;
wire      [7:0] bv_8_38_n444;
wire      [7:0] bv_8_39_n132;
wire      [7:0] bv_8_3_n65;
wire      [7:0] bv_8_40_n366;
wire      [7:0] bv_8_41_n29;
wire      [7:0] bv_8_42_n672;
wire      [7:0] bv_8_43_n121;
wire      [7:0] bv_8_44_n5;
wire      [7:0] bv_8_45_n97;
wire      [7:0] bv_8_46_n429;
wire      [7:0] bv_8_47_n652;
wire      [7:0] bv_8_48_n660;
wire      [7:0] bv_8_49_n309;
wire      [7:0] bv_8_4_n516;
wire      [7:0] bv_8_50_n408;
wire      [7:0] bv_8_51_n101;
wire      [7:0] bv_8_52_n619;
wire      [7:0] bv_8_53_n436;
wire      [7:0] bv_8_54_n616;
wire      [7:0] bv_8_55_n650;
wire      [7:0] bv_8_56_n230;
wire      [7:0] bv_8_57_n312;
wire      [7:0] bv_8_58_n136;
wire      [7:0] bv_8_59_n382;
wire      [7:0] bv_8_5_n492;
wire      [7:0] bv_8_60_n93;
wire      [7:0] bv_8_61_n634;
wire      [7:0] bv_8_62_n205;
wire      [7:0] bv_8_63_n489;
wire      [7:0] bv_8_64_n573;
wire      [7:0] bv_8_65_n623;
wire      [7:0] bv_8_66_n466;
wire      [7:0] bv_8_67_n318;
wire      [7:0] bv_8_68_n390;
wire      [7:0] bv_8_69_n612;
wire      [7:0] bv_8_6_n169;
wire      [7:0] bv_8_70_n609;
wire      [7:0] bv_8_71_n252;
wire      [7:0] bv_8_72_n330;
wire      [7:0] bv_8_73_n275;
wire      [7:0] bv_8_74_n237;
wire      [7:0] bv_8_75_n503;
wire      [7:0] bv_8_76_n596;
wire      [7:0] bv_8_77_n593;
wire      [7:0] bv_8_78_n590;
wire      [7:0] bv_8_79_n538;
wire      [7:0] bv_8_7_n105;
wire      [7:0] bv_8_80_n73;
wire      [7:0] bv_8_81_n582;
wire      [7:0] bv_8_82_n578;
wire      [7:0] bv_8_83_n575;
wire      [7:0] bv_8_84_n386;
wire      [7:0] bv_8_85_n423;
wire      [7:0] bv_8_86_n567;
wire      [7:0] bv_8_87_n226;
wire      [7:0] bv_8_88_n562;
wire      [7:0] bv_8_89_n61;
wire      [7:0] bv_8_8_n669;
wire      [7:0] bv_8_90_n25;
wire      [7:0] bv_8_91_n555;
wire      [7:0] bv_8_92_n234;
wire      [7:0] bv_8_93_n498;
wire      [7:0] bv_8_94_n548;
wire      [7:0] bv_8_95_n545;
wire      [7:0] bv_8_96_n542;
wire      [7:0] bv_8_97_n198;
wire      [7:0] bv_8_98_n536;
wire      [7:0] bv_8_99_n476;
wire      [7:0] bv_8_9_n57;
wire            clk;
(* keep *) wire    [127:0] key_randinit;
wire      [7:0] n10;
wire            n100;
wire      [7:0] n1000;
wire      [7:0] n10000;
wire            n10001;
wire      [7:0] n10002;
wire            n10003;
wire      [7:0] n10004;
wire            n10005;
wire      [7:0] n10006;
wire            n10007;
wire      [7:0] n10008;
wire            n10009;
wire      [7:0] n1001;
wire      [7:0] n10010;
wire            n10011;
wire      [7:0] n10012;
wire            n10013;
wire      [7:0] n10014;
wire            n10015;
wire      [7:0] n10016;
wire      [7:0] n10017;
wire      [7:0] n10018;
wire      [7:0] n10019;
wire      [7:0] n1002;
wire      [7:0] n10020;
wire      [7:0] n10021;
wire      [7:0] n10022;
wire      [7:0] n10023;
wire      [7:0] n10024;
wire      [7:0] n10025;
wire      [7:0] n10026;
wire      [7:0] n10027;
wire      [7:0] n10028;
wire      [7:0] n10029;
wire      [7:0] n1003;
wire      [7:0] n10030;
wire      [7:0] n10031;
wire      [7:0] n10032;
wire      [7:0] n10033;
wire      [7:0] n10034;
wire      [7:0] n10035;
wire      [7:0] n10036;
wire      [7:0] n10037;
wire      [7:0] n10038;
wire      [7:0] n10039;
wire      [7:0] n1004;
wire      [7:0] n10040;
wire      [7:0] n10041;
wire      [7:0] n10042;
wire      [7:0] n10043;
wire      [7:0] n10044;
wire      [7:0] n10045;
wire      [7:0] n10046;
wire      [7:0] n10047;
wire      [7:0] n10048;
wire      [7:0] n10049;
wire      [7:0] n1005;
wire      [7:0] n10050;
wire      [7:0] n10051;
wire      [7:0] n10052;
wire      [7:0] n10053;
wire      [7:0] n10054;
wire      [7:0] n10055;
wire      [7:0] n10056;
wire      [7:0] n10057;
wire      [7:0] n10058;
wire      [7:0] n10059;
wire      [7:0] n1006;
wire      [7:0] n10060;
wire      [7:0] n10061;
wire      [7:0] n10062;
wire      [7:0] n10063;
wire      [7:0] n10064;
wire      [7:0] n10065;
wire      [7:0] n10066;
wire      [7:0] n10067;
wire      [7:0] n10068;
wire      [7:0] n10069;
wire      [7:0] n1007;
wire      [7:0] n10070;
wire      [7:0] n10071;
wire      [7:0] n10072;
wire      [7:0] n10073;
wire      [7:0] n10074;
wire      [7:0] n10075;
wire      [7:0] n10076;
wire      [7:0] n10077;
wire      [7:0] n10078;
wire      [7:0] n10079;
wire      [7:0] n1008;
wire      [7:0] n10080;
wire      [7:0] n10081;
wire      [7:0] n10082;
wire      [7:0] n10083;
wire      [7:0] n10084;
wire      [7:0] n10085;
wire      [7:0] n10086;
wire      [7:0] n10087;
wire      [7:0] n10088;
wire      [7:0] n10089;
wire      [7:0] n1009;
wire      [7:0] n10090;
wire      [7:0] n10091;
wire      [7:0] n10092;
wire      [7:0] n10093;
wire      [7:0] n10094;
wire      [7:0] n10095;
wire      [7:0] n10096;
wire      [7:0] n10097;
wire      [7:0] n10098;
wire      [7:0] n10099;
wire      [7:0] n1010;
wire      [7:0] n10100;
wire      [7:0] n10101;
wire      [7:0] n10102;
wire      [7:0] n10103;
wire      [7:0] n10104;
wire      [7:0] n10105;
wire      [7:0] n10106;
wire      [7:0] n10107;
wire      [7:0] n10108;
wire      [7:0] n10109;
wire      [7:0] n1011;
wire      [7:0] n10110;
wire      [7:0] n10111;
wire      [7:0] n10112;
wire      [7:0] n10113;
wire      [7:0] n10114;
wire      [7:0] n10115;
wire      [7:0] n10116;
wire      [7:0] n10117;
wire      [7:0] n10118;
wire      [7:0] n10119;
wire      [7:0] n1012;
wire      [7:0] n10120;
wire      [7:0] n10121;
wire      [7:0] n10122;
wire      [7:0] n10123;
wire      [7:0] n10124;
wire      [7:0] n10125;
wire      [7:0] n10126;
wire      [7:0] n10127;
wire      [7:0] n10128;
wire      [7:0] n10129;
wire      [7:0] n1013;
wire      [7:0] n10130;
wire      [7:0] n10131;
wire      [7:0] n10132;
wire      [7:0] n10133;
wire      [7:0] n10134;
wire      [7:0] n10135;
wire      [7:0] n10136;
wire      [7:0] n10137;
wire      [7:0] n10138;
wire      [7:0] n10139;
wire      [7:0] n1014;
wire      [7:0] n10140;
wire      [7:0] n10141;
wire      [7:0] n10142;
wire      [7:0] n10143;
wire      [7:0] n10144;
wire      [7:0] n10145;
wire      [7:0] n10146;
wire      [7:0] n10147;
wire      [7:0] n10148;
wire      [7:0] n10149;
wire      [7:0] n1015;
wire      [7:0] n10150;
wire      [7:0] n10151;
wire      [7:0] n10152;
wire      [7:0] n10153;
wire      [7:0] n10154;
wire      [7:0] n10155;
wire      [7:0] n10156;
wire      [7:0] n10157;
wire      [7:0] n10158;
wire      [7:0] n10159;
wire      [7:0] n1016;
wire      [7:0] n10160;
wire      [7:0] n10161;
wire      [7:0] n10162;
wire      [7:0] n10163;
wire      [7:0] n10164;
wire      [7:0] n10165;
wire      [7:0] n10166;
wire      [7:0] n10167;
wire      [7:0] n10168;
wire      [7:0] n10169;
wire      [7:0] n1017;
wire      [7:0] n10170;
wire      [7:0] n10171;
wire      [7:0] n10172;
wire      [7:0] n10173;
wire      [7:0] n10174;
wire      [7:0] n10175;
wire      [7:0] n10176;
wire      [7:0] n10177;
wire      [7:0] n10178;
wire      [7:0] n10179;
wire      [7:0] n1018;
wire      [7:0] n10180;
wire      [7:0] n10181;
wire      [7:0] n10182;
wire      [7:0] n10183;
wire      [7:0] n10184;
wire      [7:0] n10185;
wire      [7:0] n10186;
wire      [7:0] n10187;
wire      [7:0] n10188;
wire      [7:0] n10189;
wire      [7:0] n1019;
wire      [7:0] n10190;
wire      [7:0] n10191;
wire      [7:0] n10192;
wire      [7:0] n10193;
wire      [7:0] n10194;
wire      [7:0] n10195;
wire      [7:0] n10196;
wire      [7:0] n10197;
wire      [7:0] n10198;
wire      [7:0] n10199;
wire      [7:0] n102;
wire      [7:0] n1020;
wire      [7:0] n10200;
wire      [7:0] n10201;
wire      [7:0] n10202;
wire      [7:0] n10203;
wire      [7:0] n10204;
wire      [7:0] n10205;
wire      [7:0] n10206;
wire      [7:0] n10207;
wire      [7:0] n10208;
wire      [7:0] n10209;
wire      [7:0] n1021;
wire      [7:0] n10210;
wire      [7:0] n10211;
wire      [7:0] n10212;
wire      [7:0] n10213;
wire      [7:0] n10214;
wire      [7:0] n10215;
wire      [7:0] n10216;
wire      [7:0] n10217;
wire      [7:0] n10218;
wire      [7:0] n10219;
wire      [7:0] n1022;
wire      [7:0] n10220;
wire      [7:0] n10221;
wire      [7:0] n10222;
wire      [7:0] n10223;
wire      [7:0] n10224;
wire      [7:0] n10225;
wire      [7:0] n10226;
wire      [7:0] n10227;
wire      [7:0] n10228;
wire      [7:0] n10229;
wire      [7:0] n1023;
wire      [7:0] n10230;
wire      [7:0] n10231;
wire      [7:0] n10232;
wire      [7:0] n10233;
wire      [7:0] n10234;
wire      [7:0] n10235;
wire      [7:0] n10236;
wire      [7:0] n10237;
wire      [7:0] n10238;
wire      [7:0] n10239;
wire      [7:0] n1024;
wire      [7:0] n10240;
wire      [7:0] n10241;
wire      [7:0] n10242;
wire      [7:0] n10243;
wire      [7:0] n10244;
wire      [7:0] n10245;
wire      [7:0] n10246;
wire      [7:0] n10247;
wire      [7:0] n10248;
wire      [7:0] n10249;
wire      [7:0] n1025;
wire      [7:0] n10250;
wire      [7:0] n10251;
wire      [7:0] n10252;
wire      [7:0] n10253;
wire      [7:0] n10254;
wire      [7:0] n10255;
wire      [7:0] n10256;
wire      [7:0] n10257;
wire      [7:0] n10258;
wire      [7:0] n10259;
wire      [7:0] n1026;
wire      [7:0] n10260;
wire      [7:0] n10261;
wire      [7:0] n10262;
wire      [7:0] n10263;
wire      [7:0] n10264;
wire      [7:0] n10265;
wire      [7:0] n10266;
wire      [7:0] n10267;
wire      [7:0] n10268;
wire      [7:0] n10269;
wire            n1027;
wire      [7:0] n10270;
wire      [7:0] n10271;
wire      [7:0] n10272;
wire      [7:0] n10273;
wire      [7:0] n10274;
wire     [39:0] n10275;
wire      [7:0] n10276;
wire            n10277;
wire      [7:0] n10278;
wire            n10279;
wire      [7:0] n1028;
wire      [7:0] n10280;
wire            n10281;
wire      [7:0] n10282;
wire            n10283;
wire      [7:0] n10284;
wire            n10285;
wire      [7:0] n10286;
wire            n10287;
wire      [7:0] n10288;
wire            n10289;
wire            n1029;
wire      [7:0] n10290;
wire            n10291;
wire      [7:0] n10292;
wire            n10293;
wire      [7:0] n10294;
wire            n10295;
wire      [7:0] n10296;
wire            n10297;
wire      [7:0] n10298;
wire            n10299;
wire      [7:0] n1030;
wire      [7:0] n10300;
wire            n10301;
wire      [7:0] n10302;
wire            n10303;
wire      [7:0] n10304;
wire            n10305;
wire      [7:0] n10306;
wire            n10307;
wire      [7:0] n10308;
wire            n10309;
wire            n1031;
wire      [7:0] n10310;
wire            n10311;
wire      [7:0] n10312;
wire            n10313;
wire      [7:0] n10314;
wire            n10315;
wire      [7:0] n10316;
wire            n10317;
wire      [7:0] n10318;
wire            n10319;
wire      [7:0] n1032;
wire      [7:0] n10320;
wire            n10321;
wire      [7:0] n10322;
wire            n10323;
wire      [7:0] n10324;
wire            n10325;
wire      [7:0] n10326;
wire            n10327;
wire      [7:0] n10328;
wire            n10329;
wire            n1033;
wire      [7:0] n10330;
wire            n10331;
wire      [7:0] n10332;
wire            n10333;
wire      [7:0] n10334;
wire            n10335;
wire      [7:0] n10336;
wire            n10337;
wire      [7:0] n10338;
wire            n10339;
wire      [7:0] n1034;
wire      [7:0] n10340;
wire            n10341;
wire      [7:0] n10342;
wire            n10343;
wire      [7:0] n10344;
wire            n10345;
wire      [7:0] n10346;
wire            n10347;
wire      [7:0] n10348;
wire            n10349;
wire            n1035;
wire      [7:0] n10350;
wire            n10351;
wire      [7:0] n10352;
wire            n10353;
wire      [7:0] n10354;
wire            n10355;
wire      [7:0] n10356;
wire            n10357;
wire      [7:0] n10358;
wire            n10359;
wire      [7:0] n1036;
wire      [7:0] n10360;
wire            n10361;
wire      [7:0] n10362;
wire            n10363;
wire      [7:0] n10364;
wire            n10365;
wire      [7:0] n10366;
wire            n10367;
wire      [7:0] n10368;
wire            n10369;
wire            n1037;
wire      [7:0] n10370;
wire            n10371;
wire      [7:0] n10372;
wire            n10373;
wire      [7:0] n10374;
wire            n10375;
wire      [7:0] n10376;
wire            n10377;
wire      [7:0] n10378;
wire            n10379;
wire      [7:0] n1038;
wire      [7:0] n10380;
wire            n10381;
wire      [7:0] n10382;
wire            n10383;
wire      [7:0] n10384;
wire            n10385;
wire      [7:0] n10386;
wire            n10387;
wire      [7:0] n10388;
wire            n10389;
wire            n1039;
wire      [7:0] n10390;
wire            n10391;
wire      [7:0] n10392;
wire            n10393;
wire      [7:0] n10394;
wire            n10395;
wire      [7:0] n10396;
wire            n10397;
wire      [7:0] n10398;
wire            n10399;
wire            n104;
wire      [7:0] n1040;
wire      [7:0] n10400;
wire            n10401;
wire      [7:0] n10402;
wire            n10403;
wire      [7:0] n10404;
wire            n10405;
wire      [7:0] n10406;
wire            n10407;
wire      [7:0] n10408;
wire            n10409;
wire            n1041;
wire      [7:0] n10410;
wire            n10411;
wire      [7:0] n10412;
wire            n10413;
wire      [7:0] n10414;
wire            n10415;
wire      [7:0] n10416;
wire            n10417;
wire      [7:0] n10418;
wire            n10419;
wire      [7:0] n1042;
wire      [7:0] n10420;
wire            n10421;
wire      [7:0] n10422;
wire            n10423;
wire      [7:0] n10424;
wire            n10425;
wire      [7:0] n10426;
wire            n10427;
wire      [7:0] n10428;
wire            n10429;
wire            n1043;
wire      [7:0] n10430;
wire            n10431;
wire      [7:0] n10432;
wire            n10433;
wire      [7:0] n10434;
wire            n10435;
wire      [7:0] n10436;
wire            n10437;
wire      [7:0] n10438;
wire            n10439;
wire      [7:0] n1044;
wire      [7:0] n10440;
wire            n10441;
wire      [7:0] n10442;
wire            n10443;
wire      [7:0] n10444;
wire            n10445;
wire      [7:0] n10446;
wire            n10447;
wire      [7:0] n10448;
wire            n10449;
wire            n1045;
wire      [7:0] n10450;
wire            n10451;
wire      [7:0] n10452;
wire            n10453;
wire      [7:0] n10454;
wire            n10455;
wire      [7:0] n10456;
wire            n10457;
wire      [7:0] n10458;
wire            n10459;
wire      [7:0] n1046;
wire      [7:0] n10460;
wire            n10461;
wire      [7:0] n10462;
wire            n10463;
wire      [7:0] n10464;
wire            n10465;
wire      [7:0] n10466;
wire            n10467;
wire      [7:0] n10468;
wire            n10469;
wire            n1047;
wire      [7:0] n10470;
wire            n10471;
wire      [7:0] n10472;
wire            n10473;
wire      [7:0] n10474;
wire            n10475;
wire      [7:0] n10476;
wire            n10477;
wire      [7:0] n10478;
wire            n10479;
wire      [7:0] n1048;
wire      [7:0] n10480;
wire            n10481;
wire      [7:0] n10482;
wire            n10483;
wire      [7:0] n10484;
wire            n10485;
wire      [7:0] n10486;
wire            n10487;
wire      [7:0] n10488;
wire            n10489;
wire            n1049;
wire      [7:0] n10490;
wire            n10491;
wire      [7:0] n10492;
wire            n10493;
wire      [7:0] n10494;
wire            n10495;
wire      [7:0] n10496;
wire            n10497;
wire      [7:0] n10498;
wire            n10499;
wire      [7:0] n1050;
wire      [7:0] n10500;
wire            n10501;
wire      [7:0] n10502;
wire            n10503;
wire      [7:0] n10504;
wire            n10505;
wire      [7:0] n10506;
wire            n10507;
wire      [7:0] n10508;
wire            n10509;
wire            n1051;
wire      [7:0] n10510;
wire            n10511;
wire      [7:0] n10512;
wire            n10513;
wire      [7:0] n10514;
wire            n10515;
wire      [7:0] n10516;
wire            n10517;
wire      [7:0] n10518;
wire            n10519;
wire      [7:0] n1052;
wire      [7:0] n10520;
wire            n10521;
wire      [7:0] n10522;
wire            n10523;
wire      [7:0] n10524;
wire            n10525;
wire      [7:0] n10526;
wire            n10527;
wire      [7:0] n10528;
wire            n10529;
wire            n1053;
wire      [7:0] n10530;
wire            n10531;
wire      [7:0] n10532;
wire            n10533;
wire      [7:0] n10534;
wire            n10535;
wire      [7:0] n10536;
wire            n10537;
wire      [7:0] n10538;
wire            n10539;
wire      [7:0] n1054;
wire      [7:0] n10540;
wire            n10541;
wire      [7:0] n10542;
wire            n10543;
wire      [7:0] n10544;
wire            n10545;
wire      [7:0] n10546;
wire            n10547;
wire      [7:0] n10548;
wire            n10549;
wire            n1055;
wire      [7:0] n10550;
wire            n10551;
wire      [7:0] n10552;
wire            n10553;
wire      [7:0] n10554;
wire            n10555;
wire      [7:0] n10556;
wire            n10557;
wire      [7:0] n10558;
wire            n10559;
wire      [7:0] n1056;
wire      [7:0] n10560;
wire            n10561;
wire      [7:0] n10562;
wire            n10563;
wire      [7:0] n10564;
wire            n10565;
wire      [7:0] n10566;
wire            n10567;
wire      [7:0] n10568;
wire            n10569;
wire            n1057;
wire      [7:0] n10570;
wire            n10571;
wire      [7:0] n10572;
wire            n10573;
wire      [7:0] n10574;
wire            n10575;
wire      [7:0] n10576;
wire            n10577;
wire      [7:0] n10578;
wire            n10579;
wire      [7:0] n1058;
wire      [7:0] n10580;
wire            n10581;
wire      [7:0] n10582;
wire            n10583;
wire      [7:0] n10584;
wire            n10585;
wire      [7:0] n10586;
wire            n10587;
wire      [7:0] n10588;
wire            n10589;
wire            n1059;
wire      [7:0] n10590;
wire            n10591;
wire      [7:0] n10592;
wire            n10593;
wire      [7:0] n10594;
wire            n10595;
wire      [7:0] n10596;
wire            n10597;
wire      [7:0] n10598;
wire            n10599;
wire      [7:0] n106;
wire      [7:0] n1060;
wire      [7:0] n10600;
wire            n10601;
wire      [7:0] n10602;
wire            n10603;
wire      [7:0] n10604;
wire            n10605;
wire      [7:0] n10606;
wire            n10607;
wire      [7:0] n10608;
wire            n10609;
wire            n1061;
wire      [7:0] n10610;
wire            n10611;
wire      [7:0] n10612;
wire            n10613;
wire      [7:0] n10614;
wire            n10615;
wire      [7:0] n10616;
wire            n10617;
wire      [7:0] n10618;
wire            n10619;
wire      [7:0] n1062;
wire      [7:0] n10620;
wire            n10621;
wire      [7:0] n10622;
wire            n10623;
wire      [7:0] n10624;
wire            n10625;
wire      [7:0] n10626;
wire            n10627;
wire      [7:0] n10628;
wire            n10629;
wire            n1063;
wire      [7:0] n10630;
wire            n10631;
wire      [7:0] n10632;
wire            n10633;
wire      [7:0] n10634;
wire            n10635;
wire      [7:0] n10636;
wire            n10637;
wire      [7:0] n10638;
wire            n10639;
wire      [7:0] n1064;
wire      [7:0] n10640;
wire            n10641;
wire      [7:0] n10642;
wire            n10643;
wire      [7:0] n10644;
wire            n10645;
wire      [7:0] n10646;
wire            n10647;
wire      [7:0] n10648;
wire            n10649;
wire            n1065;
wire      [7:0] n10650;
wire            n10651;
wire      [7:0] n10652;
wire            n10653;
wire      [7:0] n10654;
wire            n10655;
wire      [7:0] n10656;
wire            n10657;
wire      [7:0] n10658;
wire            n10659;
wire      [7:0] n1066;
wire      [7:0] n10660;
wire            n10661;
wire      [7:0] n10662;
wire            n10663;
wire      [7:0] n10664;
wire            n10665;
wire      [7:0] n10666;
wire            n10667;
wire      [7:0] n10668;
wire            n10669;
wire            n1067;
wire      [7:0] n10670;
wire            n10671;
wire      [7:0] n10672;
wire            n10673;
wire      [7:0] n10674;
wire            n10675;
wire      [7:0] n10676;
wire            n10677;
wire      [7:0] n10678;
wire            n10679;
wire      [7:0] n1068;
wire      [7:0] n10680;
wire            n10681;
wire      [7:0] n10682;
wire            n10683;
wire      [7:0] n10684;
wire            n10685;
wire      [7:0] n10686;
wire            n10687;
wire      [7:0] n10688;
wire            n10689;
wire            n1069;
wire      [7:0] n10690;
wire            n10691;
wire      [7:0] n10692;
wire            n10693;
wire      [7:0] n10694;
wire            n10695;
wire      [7:0] n10696;
wire            n10697;
wire      [7:0] n10698;
wire            n10699;
wire      [7:0] n1070;
wire      [7:0] n10700;
wire            n10701;
wire      [7:0] n10702;
wire            n10703;
wire      [7:0] n10704;
wire            n10705;
wire      [7:0] n10706;
wire            n10707;
wire      [7:0] n10708;
wire            n10709;
wire            n1071;
wire      [7:0] n10710;
wire            n10711;
wire      [7:0] n10712;
wire            n10713;
wire      [7:0] n10714;
wire            n10715;
wire      [7:0] n10716;
wire            n10717;
wire      [7:0] n10718;
wire            n10719;
wire      [7:0] n1072;
wire      [7:0] n10720;
wire            n10721;
wire      [7:0] n10722;
wire            n10723;
wire      [7:0] n10724;
wire            n10725;
wire      [7:0] n10726;
wire            n10727;
wire      [7:0] n10728;
wire            n10729;
wire            n1073;
wire      [7:0] n10730;
wire            n10731;
wire      [7:0] n10732;
wire            n10733;
wire      [7:0] n10734;
wire            n10735;
wire      [7:0] n10736;
wire            n10737;
wire      [7:0] n10738;
wire            n10739;
wire      [7:0] n1074;
wire      [7:0] n10740;
wire            n10741;
wire      [7:0] n10742;
wire            n10743;
wire      [7:0] n10744;
wire            n10745;
wire      [7:0] n10746;
wire            n10747;
wire      [7:0] n10748;
wire            n10749;
wire            n1075;
wire      [7:0] n10750;
wire            n10751;
wire      [7:0] n10752;
wire            n10753;
wire      [7:0] n10754;
wire            n10755;
wire      [7:0] n10756;
wire            n10757;
wire      [7:0] n10758;
wire            n10759;
wire      [7:0] n1076;
wire      [7:0] n10760;
wire            n10761;
wire      [7:0] n10762;
wire            n10763;
wire      [7:0] n10764;
wire            n10765;
wire      [7:0] n10766;
wire            n10767;
wire      [7:0] n10768;
wire            n10769;
wire            n1077;
wire      [7:0] n10770;
wire            n10771;
wire      [7:0] n10772;
wire            n10773;
wire      [7:0] n10774;
wire            n10775;
wire      [7:0] n10776;
wire            n10777;
wire      [7:0] n10778;
wire            n10779;
wire      [7:0] n1078;
wire      [7:0] n10780;
wire            n10781;
wire      [7:0] n10782;
wire            n10783;
wire      [7:0] n10784;
wire            n10785;
wire      [7:0] n10786;
wire            n10787;
wire      [7:0] n10788;
wire      [7:0] n10789;
wire            n1079;
wire      [7:0] n10790;
wire      [7:0] n10791;
wire      [7:0] n10792;
wire      [7:0] n10793;
wire      [7:0] n10794;
wire      [7:0] n10795;
wire      [7:0] n10796;
wire      [7:0] n10797;
wire      [7:0] n10798;
wire      [7:0] n10799;
wire            n108;
wire      [7:0] n1080;
wire      [7:0] n10800;
wire      [7:0] n10801;
wire      [7:0] n10802;
wire      [7:0] n10803;
wire      [7:0] n10804;
wire      [7:0] n10805;
wire      [7:0] n10806;
wire      [7:0] n10807;
wire      [7:0] n10808;
wire      [7:0] n10809;
wire            n1081;
wire      [7:0] n10810;
wire      [7:0] n10811;
wire      [7:0] n10812;
wire      [7:0] n10813;
wire      [7:0] n10814;
wire      [7:0] n10815;
wire      [7:0] n10816;
wire      [7:0] n10817;
wire      [7:0] n10818;
wire      [7:0] n10819;
wire      [7:0] n1082;
wire      [7:0] n10820;
wire      [7:0] n10821;
wire      [7:0] n10822;
wire      [7:0] n10823;
wire      [7:0] n10824;
wire      [7:0] n10825;
wire      [7:0] n10826;
wire      [7:0] n10827;
wire      [7:0] n10828;
wire      [7:0] n10829;
wire            n1083;
wire      [7:0] n10830;
wire      [7:0] n10831;
wire      [7:0] n10832;
wire      [7:0] n10833;
wire      [7:0] n10834;
wire      [7:0] n10835;
wire      [7:0] n10836;
wire      [7:0] n10837;
wire      [7:0] n10838;
wire      [7:0] n10839;
wire      [7:0] n1084;
wire      [7:0] n10840;
wire      [7:0] n10841;
wire      [7:0] n10842;
wire      [7:0] n10843;
wire      [7:0] n10844;
wire      [7:0] n10845;
wire      [7:0] n10846;
wire      [7:0] n10847;
wire      [7:0] n10848;
wire      [7:0] n10849;
wire            n1085;
wire      [7:0] n10850;
wire      [7:0] n10851;
wire      [7:0] n10852;
wire      [7:0] n10853;
wire      [7:0] n10854;
wire      [7:0] n10855;
wire      [7:0] n10856;
wire      [7:0] n10857;
wire      [7:0] n10858;
wire      [7:0] n10859;
wire      [7:0] n1086;
wire      [7:0] n10860;
wire      [7:0] n10861;
wire      [7:0] n10862;
wire      [7:0] n10863;
wire      [7:0] n10864;
wire      [7:0] n10865;
wire      [7:0] n10866;
wire      [7:0] n10867;
wire      [7:0] n10868;
wire      [7:0] n10869;
wire            n1087;
wire      [7:0] n10870;
wire      [7:0] n10871;
wire      [7:0] n10872;
wire      [7:0] n10873;
wire      [7:0] n10874;
wire      [7:0] n10875;
wire      [7:0] n10876;
wire      [7:0] n10877;
wire      [7:0] n10878;
wire      [7:0] n10879;
wire      [7:0] n1088;
wire      [7:0] n10880;
wire      [7:0] n10881;
wire      [7:0] n10882;
wire      [7:0] n10883;
wire      [7:0] n10884;
wire      [7:0] n10885;
wire      [7:0] n10886;
wire      [7:0] n10887;
wire      [7:0] n10888;
wire      [7:0] n10889;
wire            n1089;
wire      [7:0] n10890;
wire      [7:0] n10891;
wire      [7:0] n10892;
wire      [7:0] n10893;
wire      [7:0] n10894;
wire      [7:0] n10895;
wire      [7:0] n10896;
wire      [7:0] n10897;
wire      [7:0] n10898;
wire      [7:0] n10899;
wire      [7:0] n1090;
wire      [7:0] n10900;
wire      [7:0] n10901;
wire      [7:0] n10902;
wire      [7:0] n10903;
wire      [7:0] n10904;
wire      [7:0] n10905;
wire      [7:0] n10906;
wire      [7:0] n10907;
wire      [7:0] n10908;
wire      [7:0] n10909;
wire            n1091;
wire      [7:0] n10910;
wire      [7:0] n10911;
wire      [7:0] n10912;
wire      [7:0] n10913;
wire      [7:0] n10914;
wire      [7:0] n10915;
wire      [7:0] n10916;
wire      [7:0] n10917;
wire      [7:0] n10918;
wire      [7:0] n10919;
wire      [7:0] n1092;
wire      [7:0] n10920;
wire      [7:0] n10921;
wire      [7:0] n10922;
wire      [7:0] n10923;
wire      [7:0] n10924;
wire      [7:0] n10925;
wire      [7:0] n10926;
wire      [7:0] n10927;
wire      [7:0] n10928;
wire      [7:0] n10929;
wire            n1093;
wire      [7:0] n10930;
wire      [7:0] n10931;
wire      [7:0] n10932;
wire      [7:0] n10933;
wire      [7:0] n10934;
wire      [7:0] n10935;
wire      [7:0] n10936;
wire      [7:0] n10937;
wire      [7:0] n10938;
wire      [7:0] n10939;
wire      [7:0] n1094;
wire      [7:0] n10940;
wire      [7:0] n10941;
wire      [7:0] n10942;
wire      [7:0] n10943;
wire      [7:0] n10944;
wire      [7:0] n10945;
wire      [7:0] n10946;
wire      [7:0] n10947;
wire      [7:0] n10948;
wire      [7:0] n10949;
wire            n1095;
wire      [7:0] n10950;
wire      [7:0] n10951;
wire      [7:0] n10952;
wire      [7:0] n10953;
wire      [7:0] n10954;
wire      [7:0] n10955;
wire      [7:0] n10956;
wire      [7:0] n10957;
wire      [7:0] n10958;
wire      [7:0] n10959;
wire      [7:0] n1096;
wire      [7:0] n10960;
wire      [7:0] n10961;
wire      [7:0] n10962;
wire      [7:0] n10963;
wire      [7:0] n10964;
wire      [7:0] n10965;
wire      [7:0] n10966;
wire      [7:0] n10967;
wire      [7:0] n10968;
wire      [7:0] n10969;
wire            n1097;
wire      [7:0] n10970;
wire      [7:0] n10971;
wire      [7:0] n10972;
wire      [7:0] n10973;
wire      [7:0] n10974;
wire      [7:0] n10975;
wire      [7:0] n10976;
wire      [7:0] n10977;
wire      [7:0] n10978;
wire      [7:0] n10979;
wire      [7:0] n1098;
wire      [7:0] n10980;
wire      [7:0] n10981;
wire      [7:0] n10982;
wire      [7:0] n10983;
wire      [7:0] n10984;
wire      [7:0] n10985;
wire      [7:0] n10986;
wire      [7:0] n10987;
wire      [7:0] n10988;
wire      [7:0] n10989;
wire            n1099;
wire      [7:0] n10990;
wire      [7:0] n10991;
wire      [7:0] n10992;
wire      [7:0] n10993;
wire      [7:0] n10994;
wire      [7:0] n10995;
wire      [7:0] n10996;
wire      [7:0] n10997;
wire      [7:0] n10998;
wire      [7:0] n10999;
wire      [7:0] n110;
wire      [7:0] n1100;
wire      [7:0] n11000;
wire      [7:0] n11001;
wire      [7:0] n11002;
wire      [7:0] n11003;
wire      [7:0] n11004;
wire      [7:0] n11005;
wire      [7:0] n11006;
wire      [7:0] n11007;
wire      [7:0] n11008;
wire      [7:0] n11009;
wire            n1101;
wire      [7:0] n11010;
wire      [7:0] n11011;
wire      [7:0] n11012;
wire      [7:0] n11013;
wire      [7:0] n11014;
wire      [7:0] n11015;
wire      [7:0] n11016;
wire      [7:0] n11017;
wire      [7:0] n11018;
wire      [7:0] n11019;
wire      [7:0] n1102;
wire      [7:0] n11020;
wire      [7:0] n11021;
wire      [7:0] n11022;
wire      [7:0] n11023;
wire      [7:0] n11024;
wire      [7:0] n11025;
wire      [7:0] n11026;
wire      [7:0] n11027;
wire      [7:0] n11028;
wire      [7:0] n11029;
wire            n1103;
wire      [7:0] n11030;
wire      [7:0] n11031;
wire      [7:0] n11032;
wire      [7:0] n11033;
wire      [7:0] n11034;
wire      [7:0] n11035;
wire      [7:0] n11036;
wire      [7:0] n11037;
wire      [7:0] n11038;
wire      [7:0] n11039;
wire      [7:0] n1104;
wire      [7:0] n11040;
wire      [7:0] n11041;
wire      [7:0] n11042;
wire      [7:0] n11043;
wire      [7:0] n11044;
wire      [7:0] n11045;
wire      [7:0] n11046;
wire      [7:0] n11047;
wire            n11048;
wire      [7:0] n11049;
wire            n1105;
wire            n11050;
wire      [7:0] n11051;
wire            n11052;
wire      [7:0] n11053;
wire            n11054;
wire      [7:0] n11055;
wire            n11056;
wire      [7:0] n11057;
wire            n11058;
wire      [7:0] n11059;
wire      [7:0] n1106;
wire            n11060;
wire      [7:0] n11061;
wire            n11062;
wire      [7:0] n11063;
wire            n11064;
wire      [7:0] n11065;
wire            n11066;
wire      [7:0] n11067;
wire            n11068;
wire      [7:0] n11069;
wire            n1107;
wire            n11070;
wire      [7:0] n11071;
wire            n11072;
wire      [7:0] n11073;
wire            n11074;
wire      [7:0] n11075;
wire            n11076;
wire      [7:0] n11077;
wire            n11078;
wire      [7:0] n11079;
wire      [7:0] n1108;
wire            n11080;
wire      [7:0] n11081;
wire            n11082;
wire      [7:0] n11083;
wire            n11084;
wire      [7:0] n11085;
wire            n11086;
wire      [7:0] n11087;
wire            n11088;
wire      [7:0] n11089;
wire            n1109;
wire            n11090;
wire      [7:0] n11091;
wire            n11092;
wire      [7:0] n11093;
wire            n11094;
wire      [7:0] n11095;
wire            n11096;
wire      [7:0] n11097;
wire            n11098;
wire      [7:0] n11099;
wire      [7:0] n1110;
wire            n11100;
wire      [7:0] n11101;
wire            n11102;
wire      [7:0] n11103;
wire            n11104;
wire      [7:0] n11105;
wire            n11106;
wire      [7:0] n11107;
wire            n11108;
wire      [7:0] n11109;
wire            n1111;
wire            n11110;
wire      [7:0] n11111;
wire            n11112;
wire      [7:0] n11113;
wire            n11114;
wire      [7:0] n11115;
wire            n11116;
wire      [7:0] n11117;
wire            n11118;
wire      [7:0] n11119;
wire      [7:0] n1112;
wire            n11120;
wire      [7:0] n11121;
wire            n11122;
wire      [7:0] n11123;
wire            n11124;
wire      [7:0] n11125;
wire            n11126;
wire      [7:0] n11127;
wire            n11128;
wire      [7:0] n11129;
wire            n1113;
wire            n11130;
wire      [7:0] n11131;
wire            n11132;
wire      [7:0] n11133;
wire            n11134;
wire      [7:0] n11135;
wire            n11136;
wire      [7:0] n11137;
wire            n11138;
wire      [7:0] n11139;
wire      [7:0] n1114;
wire            n11140;
wire      [7:0] n11141;
wire            n11142;
wire      [7:0] n11143;
wire            n11144;
wire      [7:0] n11145;
wire            n11146;
wire      [7:0] n11147;
wire            n11148;
wire      [7:0] n11149;
wire            n1115;
wire            n11150;
wire      [7:0] n11151;
wire            n11152;
wire      [7:0] n11153;
wire            n11154;
wire      [7:0] n11155;
wire            n11156;
wire      [7:0] n11157;
wire            n11158;
wire      [7:0] n11159;
wire      [7:0] n1116;
wire            n11160;
wire      [7:0] n11161;
wire            n11162;
wire      [7:0] n11163;
wire            n11164;
wire      [7:0] n11165;
wire            n11166;
wire      [7:0] n11167;
wire            n11168;
wire      [7:0] n11169;
wire            n1117;
wire            n11170;
wire      [7:0] n11171;
wire            n11172;
wire      [7:0] n11173;
wire            n11174;
wire      [7:0] n11175;
wire            n11176;
wire      [7:0] n11177;
wire            n11178;
wire      [7:0] n11179;
wire      [7:0] n1118;
wire            n11180;
wire      [7:0] n11181;
wire            n11182;
wire      [7:0] n11183;
wire            n11184;
wire      [7:0] n11185;
wire            n11186;
wire      [7:0] n11187;
wire            n11188;
wire      [7:0] n11189;
wire            n1119;
wire            n11190;
wire      [7:0] n11191;
wire            n11192;
wire      [7:0] n11193;
wire            n11194;
wire      [7:0] n11195;
wire            n11196;
wire      [7:0] n11197;
wire            n11198;
wire      [7:0] n11199;
wire            n112;
wire      [7:0] n1120;
wire            n11200;
wire      [7:0] n11201;
wire            n11202;
wire      [7:0] n11203;
wire            n11204;
wire      [7:0] n11205;
wire            n11206;
wire      [7:0] n11207;
wire            n11208;
wire      [7:0] n11209;
wire            n1121;
wire            n11210;
wire      [7:0] n11211;
wire            n11212;
wire      [7:0] n11213;
wire            n11214;
wire      [7:0] n11215;
wire            n11216;
wire      [7:0] n11217;
wire            n11218;
wire      [7:0] n11219;
wire      [7:0] n1122;
wire            n11220;
wire      [7:0] n11221;
wire            n11222;
wire      [7:0] n11223;
wire            n11224;
wire      [7:0] n11225;
wire            n11226;
wire      [7:0] n11227;
wire            n11228;
wire      [7:0] n11229;
wire            n1123;
wire            n11230;
wire      [7:0] n11231;
wire            n11232;
wire      [7:0] n11233;
wire            n11234;
wire      [7:0] n11235;
wire            n11236;
wire      [7:0] n11237;
wire            n11238;
wire      [7:0] n11239;
wire      [7:0] n1124;
wire            n11240;
wire      [7:0] n11241;
wire            n11242;
wire      [7:0] n11243;
wire            n11244;
wire      [7:0] n11245;
wire            n11246;
wire      [7:0] n11247;
wire            n11248;
wire      [7:0] n11249;
wire            n1125;
wire            n11250;
wire      [7:0] n11251;
wire            n11252;
wire      [7:0] n11253;
wire            n11254;
wire      [7:0] n11255;
wire            n11256;
wire      [7:0] n11257;
wire            n11258;
wire      [7:0] n11259;
wire      [7:0] n1126;
wire            n11260;
wire      [7:0] n11261;
wire            n11262;
wire      [7:0] n11263;
wire            n11264;
wire      [7:0] n11265;
wire            n11266;
wire      [7:0] n11267;
wire            n11268;
wire      [7:0] n11269;
wire            n1127;
wire            n11270;
wire      [7:0] n11271;
wire            n11272;
wire      [7:0] n11273;
wire            n11274;
wire      [7:0] n11275;
wire            n11276;
wire      [7:0] n11277;
wire            n11278;
wire      [7:0] n11279;
wire      [7:0] n1128;
wire            n11280;
wire      [7:0] n11281;
wire            n11282;
wire      [7:0] n11283;
wire            n11284;
wire      [7:0] n11285;
wire            n11286;
wire      [7:0] n11287;
wire            n11288;
wire      [7:0] n11289;
wire            n1129;
wire            n11290;
wire      [7:0] n11291;
wire            n11292;
wire      [7:0] n11293;
wire            n11294;
wire      [7:0] n11295;
wire            n11296;
wire      [7:0] n11297;
wire            n11298;
wire      [7:0] n11299;
wire      [7:0] n1130;
wire            n11300;
wire      [7:0] n11301;
wire            n11302;
wire      [7:0] n11303;
wire            n11304;
wire      [7:0] n11305;
wire            n11306;
wire      [7:0] n11307;
wire            n11308;
wire      [7:0] n11309;
wire            n1131;
wire            n11310;
wire      [7:0] n11311;
wire            n11312;
wire      [7:0] n11313;
wire            n11314;
wire      [7:0] n11315;
wire            n11316;
wire      [7:0] n11317;
wire            n11318;
wire      [7:0] n11319;
wire      [7:0] n1132;
wire            n11320;
wire      [7:0] n11321;
wire            n11322;
wire      [7:0] n11323;
wire            n11324;
wire      [7:0] n11325;
wire            n11326;
wire      [7:0] n11327;
wire            n11328;
wire      [7:0] n11329;
wire            n1133;
wire            n11330;
wire      [7:0] n11331;
wire            n11332;
wire      [7:0] n11333;
wire            n11334;
wire      [7:0] n11335;
wire            n11336;
wire      [7:0] n11337;
wire            n11338;
wire      [7:0] n11339;
wire      [7:0] n1134;
wire            n11340;
wire      [7:0] n11341;
wire            n11342;
wire      [7:0] n11343;
wire            n11344;
wire      [7:0] n11345;
wire            n11346;
wire      [7:0] n11347;
wire            n11348;
wire      [7:0] n11349;
wire            n1135;
wire            n11350;
wire      [7:0] n11351;
wire            n11352;
wire      [7:0] n11353;
wire            n11354;
wire      [7:0] n11355;
wire            n11356;
wire      [7:0] n11357;
wire            n11358;
wire      [7:0] n11359;
wire      [7:0] n1136;
wire            n11360;
wire      [7:0] n11361;
wire            n11362;
wire      [7:0] n11363;
wire            n11364;
wire      [7:0] n11365;
wire            n11366;
wire      [7:0] n11367;
wire            n11368;
wire      [7:0] n11369;
wire            n1137;
wire            n11370;
wire      [7:0] n11371;
wire            n11372;
wire      [7:0] n11373;
wire            n11374;
wire      [7:0] n11375;
wire            n11376;
wire      [7:0] n11377;
wire            n11378;
wire      [7:0] n11379;
wire      [7:0] n1138;
wire            n11380;
wire      [7:0] n11381;
wire            n11382;
wire      [7:0] n11383;
wire            n11384;
wire      [7:0] n11385;
wire            n11386;
wire      [7:0] n11387;
wire            n11388;
wire      [7:0] n11389;
wire            n1139;
wire            n11390;
wire      [7:0] n11391;
wire            n11392;
wire      [7:0] n11393;
wire            n11394;
wire      [7:0] n11395;
wire            n11396;
wire      [7:0] n11397;
wire            n11398;
wire      [7:0] n11399;
wire      [7:0] n114;
wire      [7:0] n1140;
wire            n11400;
wire      [7:0] n11401;
wire            n11402;
wire      [7:0] n11403;
wire            n11404;
wire      [7:0] n11405;
wire            n11406;
wire      [7:0] n11407;
wire            n11408;
wire      [7:0] n11409;
wire            n1141;
wire            n11410;
wire      [7:0] n11411;
wire            n11412;
wire      [7:0] n11413;
wire            n11414;
wire      [7:0] n11415;
wire            n11416;
wire      [7:0] n11417;
wire            n11418;
wire      [7:0] n11419;
wire      [7:0] n1142;
wire            n11420;
wire      [7:0] n11421;
wire            n11422;
wire      [7:0] n11423;
wire            n11424;
wire      [7:0] n11425;
wire            n11426;
wire      [7:0] n11427;
wire            n11428;
wire      [7:0] n11429;
wire            n1143;
wire            n11430;
wire      [7:0] n11431;
wire            n11432;
wire      [7:0] n11433;
wire            n11434;
wire      [7:0] n11435;
wire            n11436;
wire      [7:0] n11437;
wire            n11438;
wire      [7:0] n11439;
wire      [7:0] n1144;
wire            n11440;
wire      [7:0] n11441;
wire            n11442;
wire      [7:0] n11443;
wire            n11444;
wire      [7:0] n11445;
wire            n11446;
wire      [7:0] n11447;
wire            n11448;
wire      [7:0] n11449;
wire            n1145;
wire            n11450;
wire      [7:0] n11451;
wire            n11452;
wire      [7:0] n11453;
wire            n11454;
wire      [7:0] n11455;
wire            n11456;
wire      [7:0] n11457;
wire            n11458;
wire      [7:0] n11459;
wire      [7:0] n1146;
wire            n11460;
wire      [7:0] n11461;
wire            n11462;
wire      [7:0] n11463;
wire            n11464;
wire      [7:0] n11465;
wire            n11466;
wire      [7:0] n11467;
wire            n11468;
wire      [7:0] n11469;
wire            n1147;
wire            n11470;
wire      [7:0] n11471;
wire            n11472;
wire      [7:0] n11473;
wire            n11474;
wire      [7:0] n11475;
wire            n11476;
wire      [7:0] n11477;
wire            n11478;
wire      [7:0] n11479;
wire      [7:0] n1148;
wire            n11480;
wire      [7:0] n11481;
wire            n11482;
wire      [7:0] n11483;
wire            n11484;
wire      [7:0] n11485;
wire            n11486;
wire      [7:0] n11487;
wire            n11488;
wire      [7:0] n11489;
wire            n1149;
wire            n11490;
wire      [7:0] n11491;
wire            n11492;
wire      [7:0] n11493;
wire            n11494;
wire      [7:0] n11495;
wire            n11496;
wire      [7:0] n11497;
wire            n11498;
wire      [7:0] n11499;
wire      [7:0] n1150;
wire            n11500;
wire      [7:0] n11501;
wire            n11502;
wire      [7:0] n11503;
wire            n11504;
wire      [7:0] n11505;
wire            n11506;
wire      [7:0] n11507;
wire            n11508;
wire      [7:0] n11509;
wire            n1151;
wire            n11510;
wire      [7:0] n11511;
wire            n11512;
wire      [7:0] n11513;
wire            n11514;
wire      [7:0] n11515;
wire            n11516;
wire      [7:0] n11517;
wire            n11518;
wire      [7:0] n11519;
wire      [7:0] n1152;
wire            n11520;
wire      [7:0] n11521;
wire            n11522;
wire      [7:0] n11523;
wire            n11524;
wire      [7:0] n11525;
wire            n11526;
wire      [7:0] n11527;
wire            n11528;
wire      [7:0] n11529;
wire            n1153;
wire            n11530;
wire      [7:0] n11531;
wire            n11532;
wire      [7:0] n11533;
wire            n11534;
wire      [7:0] n11535;
wire            n11536;
wire      [7:0] n11537;
wire            n11538;
wire      [7:0] n11539;
wire      [7:0] n1154;
wire            n11540;
wire      [7:0] n11541;
wire            n11542;
wire      [7:0] n11543;
wire            n11544;
wire      [7:0] n11545;
wire            n11546;
wire      [7:0] n11547;
wire            n11548;
wire      [7:0] n11549;
wire            n1155;
wire            n11550;
wire      [7:0] n11551;
wire            n11552;
wire      [7:0] n11553;
wire            n11554;
wire      [7:0] n11555;
wire            n11556;
wire      [7:0] n11557;
wire            n11558;
wire      [7:0] n11559;
wire      [7:0] n1156;
wire      [7:0] n11560;
wire      [7:0] n11561;
wire      [7:0] n11562;
wire      [7:0] n11563;
wire      [7:0] n11564;
wire      [7:0] n11565;
wire      [7:0] n11566;
wire      [7:0] n11567;
wire      [7:0] n11568;
wire      [7:0] n11569;
wire            n1157;
wire      [7:0] n11570;
wire      [7:0] n11571;
wire      [7:0] n11572;
wire      [7:0] n11573;
wire      [7:0] n11574;
wire      [7:0] n11575;
wire      [7:0] n11576;
wire      [7:0] n11577;
wire      [7:0] n11578;
wire      [7:0] n11579;
wire      [7:0] n1158;
wire      [7:0] n11580;
wire      [7:0] n11581;
wire      [7:0] n11582;
wire      [7:0] n11583;
wire      [7:0] n11584;
wire      [7:0] n11585;
wire      [7:0] n11586;
wire      [7:0] n11587;
wire      [7:0] n11588;
wire      [7:0] n11589;
wire            n1159;
wire      [7:0] n11590;
wire      [7:0] n11591;
wire      [7:0] n11592;
wire      [7:0] n11593;
wire      [7:0] n11594;
wire      [7:0] n11595;
wire      [7:0] n11596;
wire      [7:0] n11597;
wire      [7:0] n11598;
wire      [7:0] n11599;
wire            n116;
wire      [7:0] n1160;
wire      [7:0] n11600;
wire      [7:0] n11601;
wire      [7:0] n11602;
wire      [7:0] n11603;
wire      [7:0] n11604;
wire      [7:0] n11605;
wire      [7:0] n11606;
wire      [7:0] n11607;
wire      [7:0] n11608;
wire      [7:0] n11609;
wire            n1161;
wire      [7:0] n11610;
wire      [7:0] n11611;
wire      [7:0] n11612;
wire      [7:0] n11613;
wire      [7:0] n11614;
wire      [7:0] n11615;
wire      [7:0] n11616;
wire      [7:0] n11617;
wire      [7:0] n11618;
wire      [7:0] n11619;
wire      [7:0] n1162;
wire      [7:0] n11620;
wire      [7:0] n11621;
wire      [7:0] n11622;
wire      [7:0] n11623;
wire      [7:0] n11624;
wire      [7:0] n11625;
wire      [7:0] n11626;
wire      [7:0] n11627;
wire      [7:0] n11628;
wire      [7:0] n11629;
wire            n1163;
wire      [7:0] n11630;
wire      [7:0] n11631;
wire      [7:0] n11632;
wire      [7:0] n11633;
wire      [7:0] n11634;
wire      [7:0] n11635;
wire      [7:0] n11636;
wire      [7:0] n11637;
wire      [7:0] n11638;
wire      [7:0] n11639;
wire      [7:0] n1164;
wire      [7:0] n11640;
wire      [7:0] n11641;
wire      [7:0] n11642;
wire      [7:0] n11643;
wire      [7:0] n11644;
wire      [7:0] n11645;
wire      [7:0] n11646;
wire      [7:0] n11647;
wire      [7:0] n11648;
wire      [7:0] n11649;
wire            n1165;
wire      [7:0] n11650;
wire      [7:0] n11651;
wire      [7:0] n11652;
wire      [7:0] n11653;
wire      [7:0] n11654;
wire      [7:0] n11655;
wire      [7:0] n11656;
wire      [7:0] n11657;
wire      [7:0] n11658;
wire      [7:0] n11659;
wire      [7:0] n1166;
wire      [7:0] n11660;
wire      [7:0] n11661;
wire      [7:0] n11662;
wire      [7:0] n11663;
wire      [7:0] n11664;
wire      [7:0] n11665;
wire      [7:0] n11666;
wire      [7:0] n11667;
wire      [7:0] n11668;
wire      [7:0] n11669;
wire            n1167;
wire      [7:0] n11670;
wire      [7:0] n11671;
wire      [7:0] n11672;
wire      [7:0] n11673;
wire      [7:0] n11674;
wire      [7:0] n11675;
wire      [7:0] n11676;
wire      [7:0] n11677;
wire      [7:0] n11678;
wire      [7:0] n11679;
wire      [7:0] n1168;
wire      [7:0] n11680;
wire      [7:0] n11681;
wire      [7:0] n11682;
wire      [7:0] n11683;
wire      [7:0] n11684;
wire      [7:0] n11685;
wire      [7:0] n11686;
wire      [7:0] n11687;
wire      [7:0] n11688;
wire      [7:0] n11689;
wire            n1169;
wire      [7:0] n11690;
wire      [7:0] n11691;
wire      [7:0] n11692;
wire      [7:0] n11693;
wire      [7:0] n11694;
wire      [7:0] n11695;
wire      [7:0] n11696;
wire      [7:0] n11697;
wire      [7:0] n11698;
wire      [7:0] n11699;
wire      [7:0] n1170;
wire      [7:0] n11700;
wire      [7:0] n11701;
wire      [7:0] n11702;
wire      [7:0] n11703;
wire      [7:0] n11704;
wire      [7:0] n11705;
wire      [7:0] n11706;
wire      [7:0] n11707;
wire      [7:0] n11708;
wire      [7:0] n11709;
wire            n1171;
wire      [7:0] n11710;
wire      [7:0] n11711;
wire      [7:0] n11712;
wire      [7:0] n11713;
wire      [7:0] n11714;
wire      [7:0] n11715;
wire      [7:0] n11716;
wire      [7:0] n11717;
wire      [7:0] n11718;
wire      [7:0] n11719;
wire      [7:0] n1172;
wire      [7:0] n11720;
wire      [7:0] n11721;
wire      [7:0] n11722;
wire      [7:0] n11723;
wire      [7:0] n11724;
wire      [7:0] n11725;
wire      [7:0] n11726;
wire      [7:0] n11727;
wire      [7:0] n11728;
wire      [7:0] n11729;
wire            n1173;
wire      [7:0] n11730;
wire      [7:0] n11731;
wire      [7:0] n11732;
wire      [7:0] n11733;
wire      [7:0] n11734;
wire      [7:0] n11735;
wire      [7:0] n11736;
wire      [7:0] n11737;
wire      [7:0] n11738;
wire      [7:0] n11739;
wire      [7:0] n1174;
wire      [7:0] n11740;
wire      [7:0] n11741;
wire      [7:0] n11742;
wire      [7:0] n11743;
wire      [7:0] n11744;
wire      [7:0] n11745;
wire      [7:0] n11746;
wire      [7:0] n11747;
wire      [7:0] n11748;
wire      [7:0] n11749;
wire            n1175;
wire      [7:0] n11750;
wire      [7:0] n11751;
wire      [7:0] n11752;
wire      [7:0] n11753;
wire      [7:0] n11754;
wire      [7:0] n11755;
wire      [7:0] n11756;
wire      [7:0] n11757;
wire      [7:0] n11758;
wire      [7:0] n11759;
wire      [7:0] n1176;
wire      [7:0] n11760;
wire      [7:0] n11761;
wire      [7:0] n11762;
wire      [7:0] n11763;
wire      [7:0] n11764;
wire      [7:0] n11765;
wire      [7:0] n11766;
wire      [7:0] n11767;
wire      [7:0] n11768;
wire      [7:0] n11769;
wire            n1177;
wire      [7:0] n11770;
wire      [7:0] n11771;
wire      [7:0] n11772;
wire      [7:0] n11773;
wire      [7:0] n11774;
wire      [7:0] n11775;
wire      [7:0] n11776;
wire      [7:0] n11777;
wire      [7:0] n11778;
wire      [7:0] n11779;
wire      [7:0] n1178;
wire      [7:0] n11780;
wire      [7:0] n11781;
wire      [7:0] n11782;
wire      [7:0] n11783;
wire      [7:0] n11784;
wire      [7:0] n11785;
wire      [7:0] n11786;
wire      [7:0] n11787;
wire      [7:0] n11788;
wire      [7:0] n11789;
wire            n1179;
wire      [7:0] n11790;
wire      [7:0] n11791;
wire      [7:0] n11792;
wire      [7:0] n11793;
wire      [7:0] n11794;
wire      [7:0] n11795;
wire      [7:0] n11796;
wire      [7:0] n11797;
wire      [7:0] n11798;
wire      [7:0] n11799;
wire      [7:0] n118;
wire      [7:0] n1180;
wire      [7:0] n11800;
wire      [7:0] n11801;
wire      [7:0] n11802;
wire      [7:0] n11803;
wire      [7:0] n11804;
wire      [7:0] n11805;
wire      [7:0] n11806;
wire      [7:0] n11807;
wire      [7:0] n11808;
wire      [7:0] n11809;
wire            n1181;
wire      [7:0] n11810;
wire      [7:0] n11811;
wire      [7:0] n11812;
wire      [7:0] n11813;
wire      [7:0] n11814;
wire      [7:0] n11815;
wire      [7:0] n11816;
wire      [7:0] n11817;
wire     [47:0] n11818;
wire      [7:0] n11819;
wire      [7:0] n1182;
wire            n11820;
wire      [7:0] n11821;
wire            n11822;
wire      [7:0] n11823;
wire            n11824;
wire      [7:0] n11825;
wire            n11826;
wire      [7:0] n11827;
wire            n11828;
wire      [7:0] n11829;
wire            n1183;
wire            n11830;
wire      [7:0] n11831;
wire            n11832;
wire      [7:0] n11833;
wire            n11834;
wire      [7:0] n11835;
wire            n11836;
wire      [7:0] n11837;
wire            n11838;
wire      [7:0] n11839;
wire      [7:0] n1184;
wire            n11840;
wire      [7:0] n11841;
wire            n11842;
wire      [7:0] n11843;
wire            n11844;
wire      [7:0] n11845;
wire            n11846;
wire      [7:0] n11847;
wire            n11848;
wire      [7:0] n11849;
wire            n1185;
wire            n11850;
wire      [7:0] n11851;
wire            n11852;
wire      [7:0] n11853;
wire            n11854;
wire      [7:0] n11855;
wire            n11856;
wire      [7:0] n11857;
wire            n11858;
wire      [7:0] n11859;
wire      [7:0] n1186;
wire            n11860;
wire      [7:0] n11861;
wire            n11862;
wire      [7:0] n11863;
wire            n11864;
wire      [7:0] n11865;
wire            n11866;
wire      [7:0] n11867;
wire            n11868;
wire      [7:0] n11869;
wire            n1187;
wire            n11870;
wire      [7:0] n11871;
wire            n11872;
wire      [7:0] n11873;
wire            n11874;
wire      [7:0] n11875;
wire            n11876;
wire      [7:0] n11877;
wire            n11878;
wire      [7:0] n11879;
wire      [7:0] n1188;
wire            n11880;
wire      [7:0] n11881;
wire            n11882;
wire      [7:0] n11883;
wire            n11884;
wire      [7:0] n11885;
wire            n11886;
wire      [7:0] n11887;
wire            n11888;
wire      [7:0] n11889;
wire            n1189;
wire            n11890;
wire      [7:0] n11891;
wire            n11892;
wire      [7:0] n11893;
wire            n11894;
wire      [7:0] n11895;
wire            n11896;
wire      [7:0] n11897;
wire            n11898;
wire      [7:0] n11899;
wire      [7:0] n1190;
wire            n11900;
wire      [7:0] n11901;
wire            n11902;
wire      [7:0] n11903;
wire            n11904;
wire      [7:0] n11905;
wire            n11906;
wire      [7:0] n11907;
wire            n11908;
wire      [7:0] n11909;
wire            n1191;
wire            n11910;
wire      [7:0] n11911;
wire            n11912;
wire      [7:0] n11913;
wire            n11914;
wire      [7:0] n11915;
wire            n11916;
wire      [7:0] n11917;
wire            n11918;
wire      [7:0] n11919;
wire      [7:0] n1192;
wire            n11920;
wire      [7:0] n11921;
wire            n11922;
wire      [7:0] n11923;
wire            n11924;
wire      [7:0] n11925;
wire            n11926;
wire      [7:0] n11927;
wire            n11928;
wire      [7:0] n11929;
wire            n1193;
wire            n11930;
wire      [7:0] n11931;
wire            n11932;
wire      [7:0] n11933;
wire            n11934;
wire      [7:0] n11935;
wire            n11936;
wire      [7:0] n11937;
wire            n11938;
wire      [7:0] n11939;
wire      [7:0] n1194;
wire            n11940;
wire      [7:0] n11941;
wire            n11942;
wire      [7:0] n11943;
wire            n11944;
wire      [7:0] n11945;
wire            n11946;
wire      [7:0] n11947;
wire            n11948;
wire      [7:0] n11949;
wire            n1195;
wire            n11950;
wire      [7:0] n11951;
wire            n11952;
wire      [7:0] n11953;
wire            n11954;
wire      [7:0] n11955;
wire            n11956;
wire      [7:0] n11957;
wire            n11958;
wire      [7:0] n11959;
wire      [7:0] n1196;
wire            n11960;
wire      [7:0] n11961;
wire            n11962;
wire      [7:0] n11963;
wire            n11964;
wire      [7:0] n11965;
wire            n11966;
wire      [7:0] n11967;
wire            n11968;
wire      [7:0] n11969;
wire            n1197;
wire            n11970;
wire      [7:0] n11971;
wire            n11972;
wire      [7:0] n11973;
wire            n11974;
wire      [7:0] n11975;
wire            n11976;
wire      [7:0] n11977;
wire            n11978;
wire      [7:0] n11979;
wire      [7:0] n1198;
wire            n11980;
wire      [7:0] n11981;
wire            n11982;
wire      [7:0] n11983;
wire            n11984;
wire      [7:0] n11985;
wire            n11986;
wire      [7:0] n11987;
wire            n11988;
wire      [7:0] n11989;
wire            n1199;
wire            n11990;
wire      [7:0] n11991;
wire            n11992;
wire      [7:0] n11993;
wire            n11994;
wire      [7:0] n11995;
wire            n11996;
wire      [7:0] n11997;
wire            n11998;
wire      [7:0] n11999;
wire            n12;
wire            n120;
wire      [7:0] n1200;
wire            n12000;
wire      [7:0] n12001;
wire            n12002;
wire      [7:0] n12003;
wire            n12004;
wire      [7:0] n12005;
wire            n12006;
wire      [7:0] n12007;
wire            n12008;
wire      [7:0] n12009;
wire            n1201;
wire            n12010;
wire      [7:0] n12011;
wire            n12012;
wire      [7:0] n12013;
wire            n12014;
wire      [7:0] n12015;
wire            n12016;
wire      [7:0] n12017;
wire            n12018;
wire      [7:0] n12019;
wire      [7:0] n1202;
wire            n12020;
wire      [7:0] n12021;
wire            n12022;
wire      [7:0] n12023;
wire            n12024;
wire      [7:0] n12025;
wire            n12026;
wire      [7:0] n12027;
wire            n12028;
wire      [7:0] n12029;
wire            n1203;
wire            n12030;
wire      [7:0] n12031;
wire            n12032;
wire      [7:0] n12033;
wire            n12034;
wire      [7:0] n12035;
wire            n12036;
wire      [7:0] n12037;
wire            n12038;
wire      [7:0] n12039;
wire      [7:0] n1204;
wire            n12040;
wire      [7:0] n12041;
wire            n12042;
wire      [7:0] n12043;
wire            n12044;
wire      [7:0] n12045;
wire            n12046;
wire      [7:0] n12047;
wire            n12048;
wire      [7:0] n12049;
wire            n1205;
wire            n12050;
wire      [7:0] n12051;
wire            n12052;
wire      [7:0] n12053;
wire            n12054;
wire      [7:0] n12055;
wire            n12056;
wire      [7:0] n12057;
wire            n12058;
wire      [7:0] n12059;
wire      [7:0] n1206;
wire            n12060;
wire      [7:0] n12061;
wire            n12062;
wire      [7:0] n12063;
wire            n12064;
wire      [7:0] n12065;
wire            n12066;
wire      [7:0] n12067;
wire            n12068;
wire      [7:0] n12069;
wire            n1207;
wire            n12070;
wire      [7:0] n12071;
wire            n12072;
wire      [7:0] n12073;
wire            n12074;
wire      [7:0] n12075;
wire            n12076;
wire      [7:0] n12077;
wire            n12078;
wire      [7:0] n12079;
wire      [7:0] n1208;
wire            n12080;
wire      [7:0] n12081;
wire            n12082;
wire      [7:0] n12083;
wire            n12084;
wire      [7:0] n12085;
wire            n12086;
wire      [7:0] n12087;
wire            n12088;
wire      [7:0] n12089;
wire            n1209;
wire            n12090;
wire      [7:0] n12091;
wire            n12092;
wire      [7:0] n12093;
wire            n12094;
wire      [7:0] n12095;
wire            n12096;
wire      [7:0] n12097;
wire            n12098;
wire      [7:0] n12099;
wire      [7:0] n1210;
wire            n12100;
wire      [7:0] n12101;
wire            n12102;
wire      [7:0] n12103;
wire            n12104;
wire      [7:0] n12105;
wire            n12106;
wire      [7:0] n12107;
wire            n12108;
wire      [7:0] n12109;
wire            n1211;
wire            n12110;
wire      [7:0] n12111;
wire            n12112;
wire      [7:0] n12113;
wire            n12114;
wire      [7:0] n12115;
wire            n12116;
wire      [7:0] n12117;
wire            n12118;
wire      [7:0] n12119;
wire      [7:0] n1212;
wire            n12120;
wire      [7:0] n12121;
wire            n12122;
wire      [7:0] n12123;
wire            n12124;
wire      [7:0] n12125;
wire            n12126;
wire      [7:0] n12127;
wire            n12128;
wire      [7:0] n12129;
wire            n1213;
wire            n12130;
wire      [7:0] n12131;
wire            n12132;
wire      [7:0] n12133;
wire            n12134;
wire      [7:0] n12135;
wire            n12136;
wire      [7:0] n12137;
wire            n12138;
wire      [7:0] n12139;
wire      [7:0] n1214;
wire            n12140;
wire      [7:0] n12141;
wire            n12142;
wire      [7:0] n12143;
wire            n12144;
wire      [7:0] n12145;
wire            n12146;
wire      [7:0] n12147;
wire            n12148;
wire      [7:0] n12149;
wire            n1215;
wire            n12150;
wire      [7:0] n12151;
wire            n12152;
wire      [7:0] n12153;
wire            n12154;
wire      [7:0] n12155;
wire            n12156;
wire      [7:0] n12157;
wire            n12158;
wire      [7:0] n12159;
wire      [7:0] n1216;
wire            n12160;
wire      [7:0] n12161;
wire            n12162;
wire      [7:0] n12163;
wire            n12164;
wire      [7:0] n12165;
wire            n12166;
wire      [7:0] n12167;
wire            n12168;
wire      [7:0] n12169;
wire            n1217;
wire            n12170;
wire      [7:0] n12171;
wire            n12172;
wire      [7:0] n12173;
wire            n12174;
wire      [7:0] n12175;
wire            n12176;
wire      [7:0] n12177;
wire            n12178;
wire      [7:0] n12179;
wire      [7:0] n1218;
wire            n12180;
wire      [7:0] n12181;
wire            n12182;
wire      [7:0] n12183;
wire            n12184;
wire      [7:0] n12185;
wire            n12186;
wire      [7:0] n12187;
wire            n12188;
wire      [7:0] n12189;
wire            n1219;
wire            n12190;
wire      [7:0] n12191;
wire            n12192;
wire      [7:0] n12193;
wire            n12194;
wire      [7:0] n12195;
wire            n12196;
wire      [7:0] n12197;
wire            n12198;
wire      [7:0] n12199;
wire      [7:0] n122;
wire      [7:0] n1220;
wire            n12200;
wire      [7:0] n12201;
wire            n12202;
wire      [7:0] n12203;
wire            n12204;
wire      [7:0] n12205;
wire            n12206;
wire      [7:0] n12207;
wire            n12208;
wire      [7:0] n12209;
wire            n1221;
wire            n12210;
wire      [7:0] n12211;
wire            n12212;
wire      [7:0] n12213;
wire            n12214;
wire      [7:0] n12215;
wire            n12216;
wire      [7:0] n12217;
wire            n12218;
wire      [7:0] n12219;
wire      [7:0] n1222;
wire            n12220;
wire      [7:0] n12221;
wire            n12222;
wire      [7:0] n12223;
wire            n12224;
wire      [7:0] n12225;
wire            n12226;
wire      [7:0] n12227;
wire            n12228;
wire      [7:0] n12229;
wire            n1223;
wire            n12230;
wire      [7:0] n12231;
wire            n12232;
wire      [7:0] n12233;
wire            n12234;
wire      [7:0] n12235;
wire            n12236;
wire      [7:0] n12237;
wire            n12238;
wire      [7:0] n12239;
wire      [7:0] n1224;
wire            n12240;
wire      [7:0] n12241;
wire            n12242;
wire      [7:0] n12243;
wire            n12244;
wire      [7:0] n12245;
wire            n12246;
wire      [7:0] n12247;
wire            n12248;
wire      [7:0] n12249;
wire            n1225;
wire            n12250;
wire      [7:0] n12251;
wire            n12252;
wire      [7:0] n12253;
wire            n12254;
wire      [7:0] n12255;
wire            n12256;
wire      [7:0] n12257;
wire            n12258;
wire      [7:0] n12259;
wire      [7:0] n1226;
wire            n12260;
wire      [7:0] n12261;
wire            n12262;
wire      [7:0] n12263;
wire            n12264;
wire      [7:0] n12265;
wire            n12266;
wire      [7:0] n12267;
wire            n12268;
wire      [7:0] n12269;
wire            n1227;
wire            n12270;
wire      [7:0] n12271;
wire            n12272;
wire      [7:0] n12273;
wire            n12274;
wire      [7:0] n12275;
wire            n12276;
wire      [7:0] n12277;
wire            n12278;
wire      [7:0] n12279;
wire      [7:0] n1228;
wire            n12280;
wire      [7:0] n12281;
wire            n12282;
wire      [7:0] n12283;
wire            n12284;
wire      [7:0] n12285;
wire            n12286;
wire      [7:0] n12287;
wire            n12288;
wire      [7:0] n12289;
wire            n1229;
wire            n12290;
wire      [7:0] n12291;
wire            n12292;
wire      [7:0] n12293;
wire            n12294;
wire      [7:0] n12295;
wire            n12296;
wire      [7:0] n12297;
wire            n12298;
wire      [7:0] n12299;
wire      [7:0] n1230;
wire            n12300;
wire      [7:0] n12301;
wire            n12302;
wire      [7:0] n12303;
wire            n12304;
wire      [7:0] n12305;
wire            n12306;
wire      [7:0] n12307;
wire            n12308;
wire      [7:0] n12309;
wire            n1231;
wire            n12310;
wire      [7:0] n12311;
wire            n12312;
wire      [7:0] n12313;
wire            n12314;
wire      [7:0] n12315;
wire            n12316;
wire      [7:0] n12317;
wire            n12318;
wire      [7:0] n12319;
wire      [7:0] n1232;
wire            n12320;
wire      [7:0] n12321;
wire            n12322;
wire      [7:0] n12323;
wire            n12324;
wire      [7:0] n12325;
wire            n12326;
wire      [7:0] n12327;
wire            n12328;
wire      [7:0] n12329;
wire            n1233;
wire            n12330;
wire      [7:0] n12331;
wire      [7:0] n12332;
wire      [7:0] n12333;
wire      [7:0] n12334;
wire      [7:0] n12335;
wire      [7:0] n12336;
wire      [7:0] n12337;
wire      [7:0] n12338;
wire      [7:0] n12339;
wire      [7:0] n1234;
wire      [7:0] n12340;
wire      [7:0] n12341;
wire      [7:0] n12342;
wire      [7:0] n12343;
wire      [7:0] n12344;
wire      [7:0] n12345;
wire      [7:0] n12346;
wire      [7:0] n12347;
wire      [7:0] n12348;
wire      [7:0] n12349;
wire            n1235;
wire      [7:0] n12350;
wire      [7:0] n12351;
wire      [7:0] n12352;
wire      [7:0] n12353;
wire      [7:0] n12354;
wire      [7:0] n12355;
wire      [7:0] n12356;
wire      [7:0] n12357;
wire      [7:0] n12358;
wire      [7:0] n12359;
wire      [7:0] n1236;
wire      [7:0] n12360;
wire      [7:0] n12361;
wire      [7:0] n12362;
wire      [7:0] n12363;
wire      [7:0] n12364;
wire      [7:0] n12365;
wire      [7:0] n12366;
wire      [7:0] n12367;
wire      [7:0] n12368;
wire      [7:0] n12369;
wire            n1237;
wire      [7:0] n12370;
wire      [7:0] n12371;
wire      [7:0] n12372;
wire      [7:0] n12373;
wire      [7:0] n12374;
wire      [7:0] n12375;
wire      [7:0] n12376;
wire      [7:0] n12377;
wire      [7:0] n12378;
wire      [7:0] n12379;
wire      [7:0] n1238;
wire      [7:0] n12380;
wire      [7:0] n12381;
wire      [7:0] n12382;
wire      [7:0] n12383;
wire      [7:0] n12384;
wire      [7:0] n12385;
wire      [7:0] n12386;
wire      [7:0] n12387;
wire      [7:0] n12388;
wire      [7:0] n12389;
wire            n1239;
wire      [7:0] n12390;
wire      [7:0] n12391;
wire      [7:0] n12392;
wire      [7:0] n12393;
wire      [7:0] n12394;
wire      [7:0] n12395;
wire      [7:0] n12396;
wire      [7:0] n12397;
wire      [7:0] n12398;
wire      [7:0] n12399;
wire            n124;
wire      [7:0] n1240;
wire      [7:0] n12400;
wire      [7:0] n12401;
wire      [7:0] n12402;
wire      [7:0] n12403;
wire      [7:0] n12404;
wire      [7:0] n12405;
wire      [7:0] n12406;
wire      [7:0] n12407;
wire      [7:0] n12408;
wire      [7:0] n12409;
wire            n1241;
wire      [7:0] n12410;
wire      [7:0] n12411;
wire      [7:0] n12412;
wire      [7:0] n12413;
wire      [7:0] n12414;
wire      [7:0] n12415;
wire      [7:0] n12416;
wire      [7:0] n12417;
wire      [7:0] n12418;
wire      [7:0] n12419;
wire      [7:0] n1242;
wire      [7:0] n12420;
wire      [7:0] n12421;
wire      [7:0] n12422;
wire      [7:0] n12423;
wire      [7:0] n12424;
wire      [7:0] n12425;
wire      [7:0] n12426;
wire      [7:0] n12427;
wire      [7:0] n12428;
wire      [7:0] n12429;
wire            n1243;
wire      [7:0] n12430;
wire      [7:0] n12431;
wire      [7:0] n12432;
wire      [7:0] n12433;
wire      [7:0] n12434;
wire      [7:0] n12435;
wire      [7:0] n12436;
wire      [7:0] n12437;
wire      [7:0] n12438;
wire      [7:0] n12439;
wire      [7:0] n1244;
wire      [7:0] n12440;
wire      [7:0] n12441;
wire      [7:0] n12442;
wire      [7:0] n12443;
wire      [7:0] n12444;
wire      [7:0] n12445;
wire      [7:0] n12446;
wire      [7:0] n12447;
wire      [7:0] n12448;
wire      [7:0] n12449;
wire            n1245;
wire      [7:0] n12450;
wire      [7:0] n12451;
wire      [7:0] n12452;
wire      [7:0] n12453;
wire      [7:0] n12454;
wire      [7:0] n12455;
wire      [7:0] n12456;
wire      [7:0] n12457;
wire      [7:0] n12458;
wire      [7:0] n12459;
wire      [7:0] n1246;
wire      [7:0] n12460;
wire      [7:0] n12461;
wire      [7:0] n12462;
wire      [7:0] n12463;
wire      [7:0] n12464;
wire      [7:0] n12465;
wire      [7:0] n12466;
wire      [7:0] n12467;
wire      [7:0] n12468;
wire      [7:0] n12469;
wire            n1247;
wire      [7:0] n12470;
wire      [7:0] n12471;
wire      [7:0] n12472;
wire      [7:0] n12473;
wire      [7:0] n12474;
wire      [7:0] n12475;
wire      [7:0] n12476;
wire      [7:0] n12477;
wire      [7:0] n12478;
wire      [7:0] n12479;
wire      [7:0] n1248;
wire      [7:0] n12480;
wire      [7:0] n12481;
wire      [7:0] n12482;
wire      [7:0] n12483;
wire      [7:0] n12484;
wire      [7:0] n12485;
wire      [7:0] n12486;
wire      [7:0] n12487;
wire      [7:0] n12488;
wire      [7:0] n12489;
wire            n1249;
wire      [7:0] n12490;
wire      [7:0] n12491;
wire      [7:0] n12492;
wire      [7:0] n12493;
wire      [7:0] n12494;
wire      [7:0] n12495;
wire      [7:0] n12496;
wire      [7:0] n12497;
wire      [7:0] n12498;
wire      [7:0] n12499;
wire      [7:0] n125;
wire      [7:0] n1250;
wire      [7:0] n12500;
wire      [7:0] n12501;
wire      [7:0] n12502;
wire      [7:0] n12503;
wire      [7:0] n12504;
wire      [7:0] n12505;
wire      [7:0] n12506;
wire      [7:0] n12507;
wire      [7:0] n12508;
wire      [7:0] n12509;
wire            n1251;
wire      [7:0] n12510;
wire      [7:0] n12511;
wire      [7:0] n12512;
wire      [7:0] n12513;
wire      [7:0] n12514;
wire      [7:0] n12515;
wire      [7:0] n12516;
wire      [7:0] n12517;
wire      [7:0] n12518;
wire      [7:0] n12519;
wire      [7:0] n1252;
wire      [7:0] n12520;
wire      [7:0] n12521;
wire      [7:0] n12522;
wire      [7:0] n12523;
wire      [7:0] n12524;
wire      [7:0] n12525;
wire      [7:0] n12526;
wire      [7:0] n12527;
wire      [7:0] n12528;
wire      [7:0] n12529;
wire            n1253;
wire      [7:0] n12530;
wire      [7:0] n12531;
wire      [7:0] n12532;
wire      [7:0] n12533;
wire      [7:0] n12534;
wire      [7:0] n12535;
wire      [7:0] n12536;
wire      [7:0] n12537;
wire      [7:0] n12538;
wire      [7:0] n12539;
wire      [7:0] n1254;
wire      [7:0] n12540;
wire      [7:0] n12541;
wire      [7:0] n12542;
wire      [7:0] n12543;
wire      [7:0] n12544;
wire      [7:0] n12545;
wire      [7:0] n12546;
wire      [7:0] n12547;
wire      [7:0] n12548;
wire      [7:0] n12549;
wire            n1255;
wire      [7:0] n12550;
wire      [7:0] n12551;
wire      [7:0] n12552;
wire      [7:0] n12553;
wire      [7:0] n12554;
wire      [7:0] n12555;
wire      [7:0] n12556;
wire      [7:0] n12557;
wire      [7:0] n12558;
wire      [7:0] n12559;
wire      [7:0] n1256;
wire      [7:0] n12560;
wire      [7:0] n12561;
wire      [7:0] n12562;
wire      [7:0] n12563;
wire      [7:0] n12564;
wire      [7:0] n12565;
wire      [7:0] n12566;
wire      [7:0] n12567;
wire      [7:0] n12568;
wire      [7:0] n12569;
wire            n1257;
wire      [7:0] n12570;
wire      [7:0] n12571;
wire      [7:0] n12572;
wire      [7:0] n12573;
wire      [7:0] n12574;
wire      [7:0] n12575;
wire      [7:0] n12576;
wire      [7:0] n12577;
wire      [7:0] n12578;
wire      [7:0] n12579;
wire      [7:0] n1258;
wire      [7:0] n12580;
wire      [7:0] n12581;
wire      [7:0] n12582;
wire      [7:0] n12583;
wire      [7:0] n12584;
wire      [7:0] n12585;
wire      [7:0] n12586;
wire      [7:0] n12587;
wire      [7:0] n12588;
wire      [7:0] n12589;
wire            n1259;
wire      [7:0] n12590;
wire      [7:0] n12591;
wire      [7:0] n12592;
wire     [55:0] n12593;
wire      [7:0] n12594;
wire      [7:0] n12595;
wire      [7:0] n12596;
wire      [7:0] n12597;
wire      [7:0] n12598;
wire      [7:0] n12599;
wire      [7:0] n1260;
wire     [63:0] n12600;
wire      [7:0] n12601;
wire            n12602;
wire      [7:0] n12603;
wire            n12604;
wire      [7:0] n12605;
wire            n12606;
wire      [7:0] n12607;
wire            n12608;
wire      [7:0] n12609;
wire            n1261;
wire            n12610;
wire      [7:0] n12611;
wire            n12612;
wire      [7:0] n12613;
wire            n12614;
wire      [7:0] n12615;
wire            n12616;
wire      [7:0] n12617;
wire            n12618;
wire      [7:0] n12619;
wire      [7:0] n1262;
wire            n12620;
wire      [7:0] n12621;
wire            n12622;
wire      [7:0] n12623;
wire            n12624;
wire      [7:0] n12625;
wire            n12626;
wire      [7:0] n12627;
wire            n12628;
wire      [7:0] n12629;
wire            n1263;
wire            n12630;
wire      [7:0] n12631;
wire            n12632;
wire      [7:0] n12633;
wire            n12634;
wire      [7:0] n12635;
wire            n12636;
wire      [7:0] n12637;
wire            n12638;
wire      [7:0] n12639;
wire      [7:0] n1264;
wire            n12640;
wire      [7:0] n12641;
wire            n12642;
wire      [7:0] n12643;
wire            n12644;
wire      [7:0] n12645;
wire            n12646;
wire      [7:0] n12647;
wire            n12648;
wire      [7:0] n12649;
wire            n1265;
wire            n12650;
wire      [7:0] n12651;
wire            n12652;
wire      [7:0] n12653;
wire            n12654;
wire      [7:0] n12655;
wire            n12656;
wire      [7:0] n12657;
wire            n12658;
wire      [7:0] n12659;
wire      [7:0] n1266;
wire            n12660;
wire      [7:0] n12661;
wire            n12662;
wire      [7:0] n12663;
wire            n12664;
wire      [7:0] n12665;
wire            n12666;
wire      [7:0] n12667;
wire            n12668;
wire      [7:0] n12669;
wire            n1267;
wire            n12670;
wire      [7:0] n12671;
wire            n12672;
wire      [7:0] n12673;
wire            n12674;
wire      [7:0] n12675;
wire            n12676;
wire      [7:0] n12677;
wire            n12678;
wire      [7:0] n12679;
wire      [7:0] n1268;
wire            n12680;
wire      [7:0] n12681;
wire            n12682;
wire      [7:0] n12683;
wire            n12684;
wire      [7:0] n12685;
wire            n12686;
wire      [7:0] n12687;
wire            n12688;
wire      [7:0] n12689;
wire            n1269;
wire            n12690;
wire      [7:0] n12691;
wire            n12692;
wire      [7:0] n12693;
wire            n12694;
wire      [7:0] n12695;
wire            n12696;
wire      [7:0] n12697;
wire            n12698;
wire      [7:0] n12699;
wire            n127;
wire      [7:0] n1270;
wire            n12700;
wire      [7:0] n12701;
wire            n12702;
wire      [7:0] n12703;
wire            n12704;
wire      [7:0] n12705;
wire            n12706;
wire      [7:0] n12707;
wire            n12708;
wire      [7:0] n12709;
wire            n1271;
wire            n12710;
wire      [7:0] n12711;
wire            n12712;
wire      [7:0] n12713;
wire            n12714;
wire      [7:0] n12715;
wire            n12716;
wire      [7:0] n12717;
wire            n12718;
wire      [7:0] n12719;
wire      [7:0] n1272;
wire            n12720;
wire      [7:0] n12721;
wire            n12722;
wire      [7:0] n12723;
wire            n12724;
wire      [7:0] n12725;
wire            n12726;
wire      [7:0] n12727;
wire            n12728;
wire      [7:0] n12729;
wire            n1273;
wire            n12730;
wire      [7:0] n12731;
wire            n12732;
wire      [7:0] n12733;
wire            n12734;
wire      [7:0] n12735;
wire            n12736;
wire      [7:0] n12737;
wire            n12738;
wire      [7:0] n12739;
wire      [7:0] n1274;
wire            n12740;
wire      [7:0] n12741;
wire            n12742;
wire      [7:0] n12743;
wire            n12744;
wire      [7:0] n12745;
wire            n12746;
wire      [7:0] n12747;
wire            n12748;
wire      [7:0] n12749;
wire            n1275;
wire            n12750;
wire      [7:0] n12751;
wire            n12752;
wire      [7:0] n12753;
wire            n12754;
wire      [7:0] n12755;
wire            n12756;
wire      [7:0] n12757;
wire            n12758;
wire      [7:0] n12759;
wire      [7:0] n1276;
wire            n12760;
wire      [7:0] n12761;
wire            n12762;
wire      [7:0] n12763;
wire            n12764;
wire      [7:0] n12765;
wire            n12766;
wire      [7:0] n12767;
wire            n12768;
wire      [7:0] n12769;
wire            n1277;
wire            n12770;
wire      [7:0] n12771;
wire            n12772;
wire      [7:0] n12773;
wire            n12774;
wire      [7:0] n12775;
wire            n12776;
wire      [7:0] n12777;
wire            n12778;
wire      [7:0] n12779;
wire      [7:0] n1278;
wire            n12780;
wire      [7:0] n12781;
wire            n12782;
wire      [7:0] n12783;
wire            n12784;
wire      [7:0] n12785;
wire            n12786;
wire      [7:0] n12787;
wire            n12788;
wire      [7:0] n12789;
wire            n1279;
wire            n12790;
wire      [7:0] n12791;
wire            n12792;
wire      [7:0] n12793;
wire            n12794;
wire      [7:0] n12795;
wire            n12796;
wire      [7:0] n12797;
wire            n12798;
wire      [7:0] n12799;
wire      [7:0] n1280;
wire            n12800;
wire      [7:0] n12801;
wire            n12802;
wire      [7:0] n12803;
wire            n12804;
wire      [7:0] n12805;
wire            n12806;
wire      [7:0] n12807;
wire            n12808;
wire      [7:0] n12809;
wire            n1281;
wire            n12810;
wire      [7:0] n12811;
wire            n12812;
wire      [7:0] n12813;
wire            n12814;
wire      [7:0] n12815;
wire            n12816;
wire      [7:0] n12817;
wire            n12818;
wire      [7:0] n12819;
wire      [7:0] n1282;
wire            n12820;
wire      [7:0] n12821;
wire            n12822;
wire      [7:0] n12823;
wire            n12824;
wire      [7:0] n12825;
wire            n12826;
wire      [7:0] n12827;
wire            n12828;
wire      [7:0] n12829;
wire            n1283;
wire            n12830;
wire      [7:0] n12831;
wire            n12832;
wire      [7:0] n12833;
wire            n12834;
wire      [7:0] n12835;
wire            n12836;
wire      [7:0] n12837;
wire            n12838;
wire      [7:0] n12839;
wire      [7:0] n1284;
wire            n12840;
wire      [7:0] n12841;
wire            n12842;
wire      [7:0] n12843;
wire            n12844;
wire      [7:0] n12845;
wire            n12846;
wire      [7:0] n12847;
wire            n12848;
wire      [7:0] n12849;
wire            n1285;
wire            n12850;
wire      [7:0] n12851;
wire            n12852;
wire      [7:0] n12853;
wire            n12854;
wire      [7:0] n12855;
wire            n12856;
wire      [7:0] n12857;
wire            n12858;
wire      [7:0] n12859;
wire      [7:0] n1286;
wire            n12860;
wire      [7:0] n12861;
wire            n12862;
wire      [7:0] n12863;
wire            n12864;
wire      [7:0] n12865;
wire            n12866;
wire      [7:0] n12867;
wire            n12868;
wire      [7:0] n12869;
wire            n1287;
wire            n12870;
wire      [7:0] n12871;
wire            n12872;
wire      [7:0] n12873;
wire            n12874;
wire      [7:0] n12875;
wire            n12876;
wire      [7:0] n12877;
wire            n12878;
wire      [7:0] n12879;
wire      [7:0] n1288;
wire            n12880;
wire      [7:0] n12881;
wire            n12882;
wire      [7:0] n12883;
wire            n12884;
wire      [7:0] n12885;
wire            n12886;
wire      [7:0] n12887;
wire            n12888;
wire      [7:0] n12889;
wire            n1289;
wire            n12890;
wire      [7:0] n12891;
wire            n12892;
wire      [7:0] n12893;
wire            n12894;
wire      [7:0] n12895;
wire            n12896;
wire      [7:0] n12897;
wire            n12898;
wire      [7:0] n12899;
wire      [7:0] n129;
wire      [7:0] n1290;
wire            n12900;
wire      [7:0] n12901;
wire            n12902;
wire      [7:0] n12903;
wire            n12904;
wire      [7:0] n12905;
wire            n12906;
wire      [7:0] n12907;
wire            n12908;
wire      [7:0] n12909;
wire            n1291;
wire            n12910;
wire      [7:0] n12911;
wire            n12912;
wire      [7:0] n12913;
wire            n12914;
wire      [7:0] n12915;
wire            n12916;
wire      [7:0] n12917;
wire            n12918;
wire      [7:0] n12919;
wire      [7:0] n1292;
wire            n12920;
wire      [7:0] n12921;
wire            n12922;
wire      [7:0] n12923;
wire            n12924;
wire      [7:0] n12925;
wire            n12926;
wire      [7:0] n12927;
wire            n12928;
wire      [7:0] n12929;
wire            n1293;
wire            n12930;
wire      [7:0] n12931;
wire            n12932;
wire      [7:0] n12933;
wire            n12934;
wire      [7:0] n12935;
wire            n12936;
wire      [7:0] n12937;
wire            n12938;
wire      [7:0] n12939;
wire      [7:0] n1294;
wire            n12940;
wire      [7:0] n12941;
wire            n12942;
wire      [7:0] n12943;
wire            n12944;
wire      [7:0] n12945;
wire            n12946;
wire      [7:0] n12947;
wire            n12948;
wire      [7:0] n12949;
wire            n1295;
wire            n12950;
wire      [7:0] n12951;
wire            n12952;
wire      [7:0] n12953;
wire            n12954;
wire      [7:0] n12955;
wire            n12956;
wire      [7:0] n12957;
wire            n12958;
wire      [7:0] n12959;
wire      [7:0] n1296;
wire            n12960;
wire      [7:0] n12961;
wire            n12962;
wire      [7:0] n12963;
wire            n12964;
wire      [7:0] n12965;
wire            n12966;
wire      [7:0] n12967;
wire            n12968;
wire      [7:0] n12969;
wire            n1297;
wire            n12970;
wire      [7:0] n12971;
wire            n12972;
wire      [7:0] n12973;
wire            n12974;
wire      [7:0] n12975;
wire            n12976;
wire      [7:0] n12977;
wire            n12978;
wire      [7:0] n12979;
wire      [7:0] n1298;
wire            n12980;
wire      [7:0] n12981;
wire            n12982;
wire      [7:0] n12983;
wire            n12984;
wire      [7:0] n12985;
wire            n12986;
wire      [7:0] n12987;
wire            n12988;
wire      [7:0] n12989;
wire            n1299;
wire            n12990;
wire      [7:0] n12991;
wire            n12992;
wire      [7:0] n12993;
wire            n12994;
wire      [7:0] n12995;
wire            n12996;
wire      [7:0] n12997;
wire            n12998;
wire      [7:0] n12999;
wire      [7:0] n1300;
wire            n13000;
wire      [7:0] n13001;
wire            n13002;
wire      [7:0] n13003;
wire            n13004;
wire      [7:0] n13005;
wire            n13006;
wire      [7:0] n13007;
wire            n13008;
wire      [7:0] n13009;
wire            n1301;
wire            n13010;
wire      [7:0] n13011;
wire            n13012;
wire      [7:0] n13013;
wire            n13014;
wire      [7:0] n13015;
wire            n13016;
wire      [7:0] n13017;
wire            n13018;
wire      [7:0] n13019;
wire      [7:0] n1302;
wire            n13020;
wire      [7:0] n13021;
wire            n13022;
wire      [7:0] n13023;
wire            n13024;
wire      [7:0] n13025;
wire            n13026;
wire      [7:0] n13027;
wire            n13028;
wire      [7:0] n13029;
wire            n1303;
wire            n13030;
wire      [7:0] n13031;
wire            n13032;
wire      [7:0] n13033;
wire            n13034;
wire      [7:0] n13035;
wire            n13036;
wire      [7:0] n13037;
wire            n13038;
wire      [7:0] n13039;
wire      [7:0] n1304;
wire            n13040;
wire      [7:0] n13041;
wire            n13042;
wire      [7:0] n13043;
wire            n13044;
wire      [7:0] n13045;
wire            n13046;
wire      [7:0] n13047;
wire            n13048;
wire      [7:0] n13049;
wire            n1305;
wire            n13050;
wire      [7:0] n13051;
wire            n13052;
wire      [7:0] n13053;
wire            n13054;
wire      [7:0] n13055;
wire            n13056;
wire      [7:0] n13057;
wire            n13058;
wire      [7:0] n13059;
wire      [7:0] n1306;
wire            n13060;
wire      [7:0] n13061;
wire            n13062;
wire      [7:0] n13063;
wire            n13064;
wire      [7:0] n13065;
wire            n13066;
wire      [7:0] n13067;
wire            n13068;
wire      [7:0] n13069;
wire            n1307;
wire            n13070;
wire      [7:0] n13071;
wire            n13072;
wire      [7:0] n13073;
wire            n13074;
wire      [7:0] n13075;
wire            n13076;
wire      [7:0] n13077;
wire            n13078;
wire      [7:0] n13079;
wire      [7:0] n1308;
wire            n13080;
wire      [7:0] n13081;
wire            n13082;
wire      [7:0] n13083;
wire            n13084;
wire      [7:0] n13085;
wire            n13086;
wire      [7:0] n13087;
wire            n13088;
wire      [7:0] n13089;
wire            n1309;
wire            n13090;
wire      [7:0] n13091;
wire            n13092;
wire      [7:0] n13093;
wire            n13094;
wire      [7:0] n13095;
wire            n13096;
wire      [7:0] n13097;
wire            n13098;
wire      [7:0] n13099;
wire            n131;
wire      [7:0] n1310;
wire            n13100;
wire      [7:0] n13101;
wire            n13102;
wire      [7:0] n13103;
wire            n13104;
wire      [7:0] n13105;
wire            n13106;
wire      [7:0] n13107;
wire            n13108;
wire      [7:0] n13109;
wire            n1311;
wire            n13110;
wire      [7:0] n13111;
wire            n13112;
wire      [7:0] n13113;
wire      [7:0] n13114;
wire      [7:0] n13115;
wire      [7:0] n13116;
wire      [7:0] n13117;
wire      [7:0] n13118;
wire      [7:0] n13119;
wire      [7:0] n1312;
wire      [7:0] n13120;
wire      [7:0] n13121;
wire      [7:0] n13122;
wire      [7:0] n13123;
wire      [7:0] n13124;
wire      [7:0] n13125;
wire      [7:0] n13126;
wire      [7:0] n13127;
wire      [7:0] n13128;
wire      [7:0] n13129;
wire            n1313;
wire      [7:0] n13130;
wire      [7:0] n13131;
wire      [7:0] n13132;
wire      [7:0] n13133;
wire      [7:0] n13134;
wire      [7:0] n13135;
wire      [7:0] n13136;
wire      [7:0] n13137;
wire      [7:0] n13138;
wire      [7:0] n13139;
wire      [7:0] n1314;
wire      [7:0] n13140;
wire      [7:0] n13141;
wire      [7:0] n13142;
wire      [7:0] n13143;
wire      [7:0] n13144;
wire      [7:0] n13145;
wire      [7:0] n13146;
wire      [7:0] n13147;
wire      [7:0] n13148;
wire      [7:0] n13149;
wire            n1315;
wire      [7:0] n13150;
wire      [7:0] n13151;
wire      [7:0] n13152;
wire      [7:0] n13153;
wire      [7:0] n13154;
wire      [7:0] n13155;
wire      [7:0] n13156;
wire      [7:0] n13157;
wire      [7:0] n13158;
wire      [7:0] n13159;
wire      [7:0] n1316;
wire      [7:0] n13160;
wire      [7:0] n13161;
wire      [7:0] n13162;
wire      [7:0] n13163;
wire      [7:0] n13164;
wire      [7:0] n13165;
wire      [7:0] n13166;
wire      [7:0] n13167;
wire      [7:0] n13168;
wire      [7:0] n13169;
wire            n1317;
wire      [7:0] n13170;
wire      [7:0] n13171;
wire      [7:0] n13172;
wire      [7:0] n13173;
wire      [7:0] n13174;
wire      [7:0] n13175;
wire      [7:0] n13176;
wire      [7:0] n13177;
wire      [7:0] n13178;
wire      [7:0] n13179;
wire      [7:0] n1318;
wire      [7:0] n13180;
wire      [7:0] n13181;
wire      [7:0] n13182;
wire      [7:0] n13183;
wire      [7:0] n13184;
wire      [7:0] n13185;
wire      [7:0] n13186;
wire      [7:0] n13187;
wire      [7:0] n13188;
wire      [7:0] n13189;
wire            n1319;
wire      [7:0] n13190;
wire      [7:0] n13191;
wire      [7:0] n13192;
wire      [7:0] n13193;
wire      [7:0] n13194;
wire      [7:0] n13195;
wire      [7:0] n13196;
wire      [7:0] n13197;
wire      [7:0] n13198;
wire      [7:0] n13199;
wire      [7:0] n1320;
wire      [7:0] n13200;
wire      [7:0] n13201;
wire      [7:0] n13202;
wire      [7:0] n13203;
wire      [7:0] n13204;
wire      [7:0] n13205;
wire      [7:0] n13206;
wire      [7:0] n13207;
wire      [7:0] n13208;
wire      [7:0] n13209;
wire            n1321;
wire      [7:0] n13210;
wire      [7:0] n13211;
wire      [7:0] n13212;
wire      [7:0] n13213;
wire      [7:0] n13214;
wire      [7:0] n13215;
wire      [7:0] n13216;
wire      [7:0] n13217;
wire      [7:0] n13218;
wire      [7:0] n13219;
wire      [7:0] n1322;
wire      [7:0] n13220;
wire      [7:0] n13221;
wire      [7:0] n13222;
wire      [7:0] n13223;
wire      [7:0] n13224;
wire      [7:0] n13225;
wire      [7:0] n13226;
wire      [7:0] n13227;
wire      [7:0] n13228;
wire      [7:0] n13229;
wire            n1323;
wire      [7:0] n13230;
wire      [7:0] n13231;
wire      [7:0] n13232;
wire      [7:0] n13233;
wire      [7:0] n13234;
wire      [7:0] n13235;
wire      [7:0] n13236;
wire      [7:0] n13237;
wire      [7:0] n13238;
wire      [7:0] n13239;
wire      [7:0] n1324;
wire      [7:0] n13240;
wire      [7:0] n13241;
wire      [7:0] n13242;
wire      [7:0] n13243;
wire      [7:0] n13244;
wire      [7:0] n13245;
wire      [7:0] n13246;
wire      [7:0] n13247;
wire      [7:0] n13248;
wire      [7:0] n13249;
wire            n1325;
wire      [7:0] n13250;
wire      [7:0] n13251;
wire      [7:0] n13252;
wire      [7:0] n13253;
wire      [7:0] n13254;
wire      [7:0] n13255;
wire      [7:0] n13256;
wire      [7:0] n13257;
wire      [7:0] n13258;
wire      [7:0] n13259;
wire      [7:0] n1326;
wire      [7:0] n13260;
wire      [7:0] n13261;
wire      [7:0] n13262;
wire      [7:0] n13263;
wire      [7:0] n13264;
wire      [7:0] n13265;
wire      [7:0] n13266;
wire      [7:0] n13267;
wire      [7:0] n13268;
wire      [7:0] n13269;
wire            n1327;
wire      [7:0] n13270;
wire      [7:0] n13271;
wire      [7:0] n13272;
wire      [7:0] n13273;
wire      [7:0] n13274;
wire      [7:0] n13275;
wire      [7:0] n13276;
wire      [7:0] n13277;
wire      [7:0] n13278;
wire      [7:0] n13279;
wire      [7:0] n1328;
wire      [7:0] n13280;
wire      [7:0] n13281;
wire      [7:0] n13282;
wire      [7:0] n13283;
wire      [7:0] n13284;
wire      [7:0] n13285;
wire      [7:0] n13286;
wire      [7:0] n13287;
wire      [7:0] n13288;
wire      [7:0] n13289;
wire            n1329;
wire      [7:0] n13290;
wire      [7:0] n13291;
wire      [7:0] n13292;
wire      [7:0] n13293;
wire      [7:0] n13294;
wire      [7:0] n13295;
wire      [7:0] n13296;
wire      [7:0] n13297;
wire      [7:0] n13298;
wire      [7:0] n13299;
wire      [7:0] n133;
wire      [7:0] n1330;
wire      [7:0] n13300;
wire      [7:0] n13301;
wire      [7:0] n13302;
wire      [7:0] n13303;
wire      [7:0] n13304;
wire      [7:0] n13305;
wire      [7:0] n13306;
wire      [7:0] n13307;
wire      [7:0] n13308;
wire      [7:0] n13309;
wire            n1331;
wire      [7:0] n13310;
wire      [7:0] n13311;
wire      [7:0] n13312;
wire      [7:0] n13313;
wire      [7:0] n13314;
wire      [7:0] n13315;
wire      [7:0] n13316;
wire      [7:0] n13317;
wire      [7:0] n13318;
wire      [7:0] n13319;
wire      [7:0] n1332;
wire      [7:0] n13320;
wire      [7:0] n13321;
wire      [7:0] n13322;
wire      [7:0] n13323;
wire      [7:0] n13324;
wire      [7:0] n13325;
wire      [7:0] n13326;
wire      [7:0] n13327;
wire      [7:0] n13328;
wire      [7:0] n13329;
wire            n1333;
wire      [7:0] n13330;
wire      [7:0] n13331;
wire      [7:0] n13332;
wire      [7:0] n13333;
wire      [7:0] n13334;
wire      [7:0] n13335;
wire      [7:0] n13336;
wire      [7:0] n13337;
wire      [7:0] n13338;
wire      [7:0] n13339;
wire      [7:0] n1334;
wire      [7:0] n13340;
wire      [7:0] n13341;
wire      [7:0] n13342;
wire      [7:0] n13343;
wire      [7:0] n13344;
wire      [7:0] n13345;
wire      [7:0] n13346;
wire      [7:0] n13347;
wire      [7:0] n13348;
wire      [7:0] n13349;
wire            n1335;
wire      [7:0] n13350;
wire      [7:0] n13351;
wire      [7:0] n13352;
wire      [7:0] n13353;
wire      [7:0] n13354;
wire      [7:0] n13355;
wire      [7:0] n13356;
wire      [7:0] n13357;
wire      [7:0] n13358;
wire      [7:0] n13359;
wire      [7:0] n1336;
wire      [7:0] n13360;
wire      [7:0] n13361;
wire      [7:0] n13362;
wire      [7:0] n13363;
wire      [7:0] n13364;
wire      [7:0] n13365;
wire      [7:0] n13366;
wire      [7:0] n13367;
wire      [7:0] n13368;
wire      [7:0] n13369;
wire            n1337;
wire            n13370;
wire      [7:0] n13371;
wire            n13372;
wire      [7:0] n13373;
wire            n13374;
wire      [7:0] n13375;
wire            n13376;
wire      [7:0] n13377;
wire            n13378;
wire      [7:0] n13379;
wire      [7:0] n1338;
wire            n13380;
wire      [7:0] n13381;
wire            n13382;
wire      [7:0] n13383;
wire            n13384;
wire      [7:0] n13385;
wire            n13386;
wire      [7:0] n13387;
wire            n13388;
wire      [7:0] n13389;
wire            n1339;
wire            n13390;
wire      [7:0] n13391;
wire            n13392;
wire      [7:0] n13393;
wire            n13394;
wire      [7:0] n13395;
wire            n13396;
wire      [7:0] n13397;
wire            n13398;
wire      [7:0] n13399;
wire      [7:0] n1340;
wire            n13400;
wire      [7:0] n13401;
wire            n13402;
wire      [7:0] n13403;
wire            n13404;
wire      [7:0] n13405;
wire            n13406;
wire      [7:0] n13407;
wire            n13408;
wire      [7:0] n13409;
wire            n1341;
wire            n13410;
wire      [7:0] n13411;
wire            n13412;
wire      [7:0] n13413;
wire            n13414;
wire      [7:0] n13415;
wire            n13416;
wire      [7:0] n13417;
wire            n13418;
wire      [7:0] n13419;
wire      [7:0] n1342;
wire            n13420;
wire      [7:0] n13421;
wire            n13422;
wire      [7:0] n13423;
wire            n13424;
wire      [7:0] n13425;
wire            n13426;
wire      [7:0] n13427;
wire            n13428;
wire      [7:0] n13429;
wire            n1343;
wire            n13430;
wire      [7:0] n13431;
wire            n13432;
wire      [7:0] n13433;
wire            n13434;
wire      [7:0] n13435;
wire            n13436;
wire      [7:0] n13437;
wire            n13438;
wire      [7:0] n13439;
wire      [7:0] n1344;
wire            n13440;
wire      [7:0] n13441;
wire            n13442;
wire      [7:0] n13443;
wire            n13444;
wire      [7:0] n13445;
wire            n13446;
wire      [7:0] n13447;
wire            n13448;
wire      [7:0] n13449;
wire            n1345;
wire            n13450;
wire      [7:0] n13451;
wire            n13452;
wire      [7:0] n13453;
wire            n13454;
wire      [7:0] n13455;
wire            n13456;
wire      [7:0] n13457;
wire            n13458;
wire      [7:0] n13459;
wire      [7:0] n1346;
wire            n13460;
wire      [7:0] n13461;
wire            n13462;
wire      [7:0] n13463;
wire            n13464;
wire      [7:0] n13465;
wire            n13466;
wire      [7:0] n13467;
wire            n13468;
wire      [7:0] n13469;
wire            n1347;
wire            n13470;
wire      [7:0] n13471;
wire            n13472;
wire      [7:0] n13473;
wire            n13474;
wire      [7:0] n13475;
wire            n13476;
wire      [7:0] n13477;
wire            n13478;
wire      [7:0] n13479;
wire      [7:0] n1348;
wire            n13480;
wire      [7:0] n13481;
wire            n13482;
wire      [7:0] n13483;
wire            n13484;
wire      [7:0] n13485;
wire            n13486;
wire      [7:0] n13487;
wire            n13488;
wire      [7:0] n13489;
wire            n1349;
wire            n13490;
wire      [7:0] n13491;
wire            n13492;
wire      [7:0] n13493;
wire            n13494;
wire      [7:0] n13495;
wire            n13496;
wire      [7:0] n13497;
wire            n13498;
wire      [7:0] n13499;
wire            n135;
wire      [7:0] n1350;
wire            n13500;
wire      [7:0] n13501;
wire            n13502;
wire      [7:0] n13503;
wire            n13504;
wire      [7:0] n13505;
wire            n13506;
wire      [7:0] n13507;
wire            n13508;
wire      [7:0] n13509;
wire            n1351;
wire            n13510;
wire      [7:0] n13511;
wire            n13512;
wire      [7:0] n13513;
wire            n13514;
wire      [7:0] n13515;
wire            n13516;
wire      [7:0] n13517;
wire            n13518;
wire      [7:0] n13519;
wire      [7:0] n1352;
wire            n13520;
wire      [7:0] n13521;
wire            n13522;
wire      [7:0] n13523;
wire            n13524;
wire      [7:0] n13525;
wire            n13526;
wire      [7:0] n13527;
wire            n13528;
wire      [7:0] n13529;
wire            n1353;
wire            n13530;
wire      [7:0] n13531;
wire            n13532;
wire      [7:0] n13533;
wire            n13534;
wire      [7:0] n13535;
wire            n13536;
wire      [7:0] n13537;
wire            n13538;
wire      [7:0] n13539;
wire      [7:0] n1354;
wire            n13540;
wire      [7:0] n13541;
wire            n13542;
wire      [7:0] n13543;
wire            n13544;
wire      [7:0] n13545;
wire            n13546;
wire      [7:0] n13547;
wire            n13548;
wire      [7:0] n13549;
wire            n1355;
wire            n13550;
wire      [7:0] n13551;
wire            n13552;
wire      [7:0] n13553;
wire            n13554;
wire      [7:0] n13555;
wire            n13556;
wire      [7:0] n13557;
wire            n13558;
wire      [7:0] n13559;
wire      [7:0] n1356;
wire            n13560;
wire      [7:0] n13561;
wire            n13562;
wire      [7:0] n13563;
wire            n13564;
wire      [7:0] n13565;
wire            n13566;
wire      [7:0] n13567;
wire            n13568;
wire      [7:0] n13569;
wire            n1357;
wire            n13570;
wire      [7:0] n13571;
wire            n13572;
wire      [7:0] n13573;
wire            n13574;
wire      [7:0] n13575;
wire            n13576;
wire      [7:0] n13577;
wire            n13578;
wire      [7:0] n13579;
wire      [7:0] n1358;
wire            n13580;
wire      [7:0] n13581;
wire            n13582;
wire      [7:0] n13583;
wire            n13584;
wire      [7:0] n13585;
wire            n13586;
wire      [7:0] n13587;
wire            n13588;
wire      [7:0] n13589;
wire            n1359;
wire            n13590;
wire      [7:0] n13591;
wire            n13592;
wire      [7:0] n13593;
wire            n13594;
wire      [7:0] n13595;
wire            n13596;
wire      [7:0] n13597;
wire            n13598;
wire      [7:0] n13599;
wire      [7:0] n1360;
wire            n13600;
wire      [7:0] n13601;
wire            n13602;
wire      [7:0] n13603;
wire            n13604;
wire      [7:0] n13605;
wire            n13606;
wire      [7:0] n13607;
wire            n13608;
wire      [7:0] n13609;
wire            n1361;
wire            n13610;
wire      [7:0] n13611;
wire            n13612;
wire      [7:0] n13613;
wire            n13614;
wire      [7:0] n13615;
wire            n13616;
wire      [7:0] n13617;
wire            n13618;
wire      [7:0] n13619;
wire      [7:0] n1362;
wire            n13620;
wire      [7:0] n13621;
wire            n13622;
wire      [7:0] n13623;
wire            n13624;
wire      [7:0] n13625;
wire            n13626;
wire      [7:0] n13627;
wire            n13628;
wire      [7:0] n13629;
wire            n1363;
wire            n13630;
wire      [7:0] n13631;
wire            n13632;
wire      [7:0] n13633;
wire            n13634;
wire      [7:0] n13635;
wire            n13636;
wire      [7:0] n13637;
wire            n13638;
wire      [7:0] n13639;
wire      [7:0] n1364;
wire            n13640;
wire      [7:0] n13641;
wire            n13642;
wire      [7:0] n13643;
wire            n13644;
wire      [7:0] n13645;
wire            n13646;
wire      [7:0] n13647;
wire            n13648;
wire      [7:0] n13649;
wire            n1365;
wire            n13650;
wire      [7:0] n13651;
wire            n13652;
wire      [7:0] n13653;
wire            n13654;
wire      [7:0] n13655;
wire            n13656;
wire      [7:0] n13657;
wire            n13658;
wire      [7:0] n13659;
wire      [7:0] n1366;
wire            n13660;
wire      [7:0] n13661;
wire            n13662;
wire      [7:0] n13663;
wire            n13664;
wire      [7:0] n13665;
wire            n13666;
wire      [7:0] n13667;
wire            n13668;
wire      [7:0] n13669;
wire            n1367;
wire            n13670;
wire      [7:0] n13671;
wire            n13672;
wire      [7:0] n13673;
wire            n13674;
wire      [7:0] n13675;
wire            n13676;
wire      [7:0] n13677;
wire            n13678;
wire      [7:0] n13679;
wire      [7:0] n1368;
wire            n13680;
wire      [7:0] n13681;
wire            n13682;
wire      [7:0] n13683;
wire            n13684;
wire      [7:0] n13685;
wire            n13686;
wire      [7:0] n13687;
wire            n13688;
wire      [7:0] n13689;
wire            n1369;
wire            n13690;
wire      [7:0] n13691;
wire            n13692;
wire      [7:0] n13693;
wire            n13694;
wire      [7:0] n13695;
wire            n13696;
wire      [7:0] n13697;
wire            n13698;
wire      [7:0] n13699;
wire      [7:0] n137;
wire      [7:0] n1370;
wire            n13700;
wire      [7:0] n13701;
wire            n13702;
wire      [7:0] n13703;
wire            n13704;
wire      [7:0] n13705;
wire            n13706;
wire      [7:0] n13707;
wire            n13708;
wire      [7:0] n13709;
wire            n1371;
wire            n13710;
wire      [7:0] n13711;
wire            n13712;
wire      [7:0] n13713;
wire            n13714;
wire      [7:0] n13715;
wire            n13716;
wire      [7:0] n13717;
wire            n13718;
wire      [7:0] n13719;
wire      [7:0] n1372;
wire            n13720;
wire      [7:0] n13721;
wire            n13722;
wire      [7:0] n13723;
wire            n13724;
wire      [7:0] n13725;
wire            n13726;
wire      [7:0] n13727;
wire            n13728;
wire      [7:0] n13729;
wire            n1373;
wire            n13730;
wire      [7:0] n13731;
wire            n13732;
wire      [7:0] n13733;
wire            n13734;
wire      [7:0] n13735;
wire            n13736;
wire      [7:0] n13737;
wire            n13738;
wire      [7:0] n13739;
wire      [7:0] n1374;
wire            n13740;
wire      [7:0] n13741;
wire            n13742;
wire      [7:0] n13743;
wire            n13744;
wire      [7:0] n13745;
wire            n13746;
wire      [7:0] n13747;
wire            n13748;
wire      [7:0] n13749;
wire            n1375;
wire            n13750;
wire      [7:0] n13751;
wire            n13752;
wire      [7:0] n13753;
wire            n13754;
wire      [7:0] n13755;
wire            n13756;
wire      [7:0] n13757;
wire            n13758;
wire      [7:0] n13759;
wire      [7:0] n1376;
wire            n13760;
wire      [7:0] n13761;
wire            n13762;
wire      [7:0] n13763;
wire            n13764;
wire      [7:0] n13765;
wire            n13766;
wire      [7:0] n13767;
wire            n13768;
wire      [7:0] n13769;
wire            n1377;
wire            n13770;
wire      [7:0] n13771;
wire            n13772;
wire      [7:0] n13773;
wire            n13774;
wire      [7:0] n13775;
wire            n13776;
wire      [7:0] n13777;
wire            n13778;
wire      [7:0] n13779;
wire      [7:0] n1378;
wire            n13780;
wire      [7:0] n13781;
wire            n13782;
wire      [7:0] n13783;
wire            n13784;
wire      [7:0] n13785;
wire            n13786;
wire      [7:0] n13787;
wire            n13788;
wire      [7:0] n13789;
wire            n1379;
wire            n13790;
wire      [7:0] n13791;
wire            n13792;
wire      [7:0] n13793;
wire            n13794;
wire      [7:0] n13795;
wire            n13796;
wire      [7:0] n13797;
wire            n13798;
wire      [7:0] n13799;
wire      [7:0] n1380;
wire            n13800;
wire      [7:0] n13801;
wire            n13802;
wire      [7:0] n13803;
wire            n13804;
wire      [7:0] n13805;
wire            n13806;
wire      [7:0] n13807;
wire            n13808;
wire      [7:0] n13809;
wire            n1381;
wire            n13810;
wire      [7:0] n13811;
wire            n13812;
wire      [7:0] n13813;
wire            n13814;
wire      [7:0] n13815;
wire            n13816;
wire      [7:0] n13817;
wire            n13818;
wire      [7:0] n13819;
wire      [7:0] n1382;
wire            n13820;
wire      [7:0] n13821;
wire            n13822;
wire      [7:0] n13823;
wire            n13824;
wire      [7:0] n13825;
wire            n13826;
wire      [7:0] n13827;
wire            n13828;
wire      [7:0] n13829;
wire            n1383;
wire            n13830;
wire      [7:0] n13831;
wire            n13832;
wire      [7:0] n13833;
wire            n13834;
wire      [7:0] n13835;
wire            n13836;
wire      [7:0] n13837;
wire            n13838;
wire      [7:0] n13839;
wire      [7:0] n1384;
wire            n13840;
wire      [7:0] n13841;
wire            n13842;
wire      [7:0] n13843;
wire            n13844;
wire      [7:0] n13845;
wire            n13846;
wire      [7:0] n13847;
wire            n13848;
wire      [7:0] n13849;
wire            n1385;
wire            n13850;
wire      [7:0] n13851;
wire            n13852;
wire      [7:0] n13853;
wire            n13854;
wire      [7:0] n13855;
wire            n13856;
wire      [7:0] n13857;
wire            n13858;
wire      [7:0] n13859;
wire      [7:0] n1386;
wire            n13860;
wire      [7:0] n13861;
wire            n13862;
wire      [7:0] n13863;
wire            n13864;
wire      [7:0] n13865;
wire            n13866;
wire      [7:0] n13867;
wire            n13868;
wire      [7:0] n13869;
wire            n1387;
wire            n13870;
wire      [7:0] n13871;
wire            n13872;
wire      [7:0] n13873;
wire            n13874;
wire      [7:0] n13875;
wire            n13876;
wire      [7:0] n13877;
wire            n13878;
wire      [7:0] n13879;
wire      [7:0] n1388;
wire            n13880;
wire      [7:0] n13881;
wire      [7:0] n13882;
wire      [7:0] n13883;
wire      [7:0] n13884;
wire      [7:0] n13885;
wire      [7:0] n13886;
wire      [7:0] n13887;
wire      [7:0] n13888;
wire      [7:0] n13889;
wire            n1389;
wire      [7:0] n13890;
wire      [7:0] n13891;
wire      [7:0] n13892;
wire      [7:0] n13893;
wire      [7:0] n13894;
wire      [7:0] n13895;
wire      [7:0] n13896;
wire      [7:0] n13897;
wire      [7:0] n13898;
wire      [7:0] n13899;
wire            n139;
wire      [7:0] n1390;
wire      [7:0] n13900;
wire      [7:0] n13901;
wire      [7:0] n13902;
wire      [7:0] n13903;
wire      [7:0] n13904;
wire      [7:0] n13905;
wire      [7:0] n13906;
wire      [7:0] n13907;
wire      [7:0] n13908;
wire      [7:0] n13909;
wire            n1391;
wire      [7:0] n13910;
wire      [7:0] n13911;
wire      [7:0] n13912;
wire      [7:0] n13913;
wire      [7:0] n13914;
wire      [7:0] n13915;
wire      [7:0] n13916;
wire      [7:0] n13917;
wire      [7:0] n13918;
wire      [7:0] n13919;
wire      [7:0] n1392;
wire      [7:0] n13920;
wire      [7:0] n13921;
wire      [7:0] n13922;
wire      [7:0] n13923;
wire      [7:0] n13924;
wire      [7:0] n13925;
wire      [7:0] n13926;
wire      [7:0] n13927;
wire      [7:0] n13928;
wire      [7:0] n13929;
wire            n1393;
wire      [7:0] n13930;
wire      [7:0] n13931;
wire      [7:0] n13932;
wire      [7:0] n13933;
wire      [7:0] n13934;
wire      [7:0] n13935;
wire      [7:0] n13936;
wire      [7:0] n13937;
wire      [7:0] n13938;
wire      [7:0] n13939;
wire      [7:0] n1394;
wire      [7:0] n13940;
wire      [7:0] n13941;
wire      [7:0] n13942;
wire      [7:0] n13943;
wire      [7:0] n13944;
wire      [7:0] n13945;
wire      [7:0] n13946;
wire      [7:0] n13947;
wire      [7:0] n13948;
wire      [7:0] n13949;
wire            n1395;
wire      [7:0] n13950;
wire      [7:0] n13951;
wire      [7:0] n13952;
wire      [7:0] n13953;
wire      [7:0] n13954;
wire      [7:0] n13955;
wire      [7:0] n13956;
wire      [7:0] n13957;
wire      [7:0] n13958;
wire      [7:0] n13959;
wire      [7:0] n1396;
wire      [7:0] n13960;
wire      [7:0] n13961;
wire      [7:0] n13962;
wire      [7:0] n13963;
wire      [7:0] n13964;
wire      [7:0] n13965;
wire      [7:0] n13966;
wire      [7:0] n13967;
wire      [7:0] n13968;
wire      [7:0] n13969;
wire            n1397;
wire      [7:0] n13970;
wire      [7:0] n13971;
wire      [7:0] n13972;
wire      [7:0] n13973;
wire      [7:0] n13974;
wire      [7:0] n13975;
wire      [7:0] n13976;
wire      [7:0] n13977;
wire      [7:0] n13978;
wire      [7:0] n13979;
wire      [7:0] n1398;
wire      [7:0] n13980;
wire      [7:0] n13981;
wire      [7:0] n13982;
wire      [7:0] n13983;
wire      [7:0] n13984;
wire      [7:0] n13985;
wire      [7:0] n13986;
wire      [7:0] n13987;
wire      [7:0] n13988;
wire      [7:0] n13989;
wire            n1399;
wire      [7:0] n13990;
wire      [7:0] n13991;
wire      [7:0] n13992;
wire      [7:0] n13993;
wire      [7:0] n13994;
wire      [7:0] n13995;
wire      [7:0] n13996;
wire      [7:0] n13997;
wire      [7:0] n13998;
wire      [7:0] n13999;
wire      [7:0] n14;
wire      [7:0] n1400;
wire      [7:0] n14000;
wire      [7:0] n14001;
wire      [7:0] n14002;
wire      [7:0] n14003;
wire      [7:0] n14004;
wire      [7:0] n14005;
wire      [7:0] n14006;
wire      [7:0] n14007;
wire      [7:0] n14008;
wire      [7:0] n14009;
wire            n1401;
wire      [7:0] n14010;
wire      [7:0] n14011;
wire      [7:0] n14012;
wire      [7:0] n14013;
wire      [7:0] n14014;
wire      [7:0] n14015;
wire      [7:0] n14016;
wire      [7:0] n14017;
wire      [7:0] n14018;
wire      [7:0] n14019;
wire      [7:0] n1402;
wire      [7:0] n14020;
wire      [7:0] n14021;
wire      [7:0] n14022;
wire      [7:0] n14023;
wire      [7:0] n14024;
wire      [7:0] n14025;
wire      [7:0] n14026;
wire      [7:0] n14027;
wire      [7:0] n14028;
wire      [7:0] n14029;
wire            n1403;
wire      [7:0] n14030;
wire      [7:0] n14031;
wire      [7:0] n14032;
wire      [7:0] n14033;
wire      [7:0] n14034;
wire      [7:0] n14035;
wire      [7:0] n14036;
wire      [7:0] n14037;
wire      [7:0] n14038;
wire      [7:0] n14039;
wire      [7:0] n1404;
wire      [7:0] n14040;
wire      [7:0] n14041;
wire      [7:0] n14042;
wire      [7:0] n14043;
wire      [7:0] n14044;
wire      [7:0] n14045;
wire      [7:0] n14046;
wire      [7:0] n14047;
wire      [7:0] n14048;
wire      [7:0] n14049;
wire            n1405;
wire      [7:0] n14050;
wire      [7:0] n14051;
wire      [7:0] n14052;
wire      [7:0] n14053;
wire      [7:0] n14054;
wire      [7:0] n14055;
wire      [7:0] n14056;
wire      [7:0] n14057;
wire      [7:0] n14058;
wire      [7:0] n14059;
wire      [7:0] n1406;
wire      [7:0] n14060;
wire      [7:0] n14061;
wire      [7:0] n14062;
wire      [7:0] n14063;
wire      [7:0] n14064;
wire      [7:0] n14065;
wire      [7:0] n14066;
wire      [7:0] n14067;
wire      [7:0] n14068;
wire      [7:0] n14069;
wire            n1407;
wire      [7:0] n14070;
wire      [7:0] n14071;
wire      [7:0] n14072;
wire      [7:0] n14073;
wire      [7:0] n14074;
wire      [7:0] n14075;
wire      [7:0] n14076;
wire      [7:0] n14077;
wire      [7:0] n14078;
wire      [7:0] n14079;
wire      [7:0] n1408;
wire      [7:0] n14080;
wire      [7:0] n14081;
wire      [7:0] n14082;
wire      [7:0] n14083;
wire      [7:0] n14084;
wire      [7:0] n14085;
wire      [7:0] n14086;
wire      [7:0] n14087;
wire      [7:0] n14088;
wire      [7:0] n14089;
wire            n1409;
wire      [7:0] n14090;
wire      [7:0] n14091;
wire      [7:0] n14092;
wire      [7:0] n14093;
wire      [7:0] n14094;
wire      [7:0] n14095;
wire      [7:0] n14096;
wire      [7:0] n14097;
wire      [7:0] n14098;
wire      [7:0] n14099;
wire      [7:0] n141;
wire      [7:0] n1410;
wire      [7:0] n14100;
wire      [7:0] n14101;
wire      [7:0] n14102;
wire      [7:0] n14103;
wire      [7:0] n14104;
wire      [7:0] n14105;
wire      [7:0] n14106;
wire      [7:0] n14107;
wire      [7:0] n14108;
wire      [7:0] n14109;
wire            n1411;
wire      [7:0] n14110;
wire      [7:0] n14111;
wire      [7:0] n14112;
wire      [7:0] n14113;
wire      [7:0] n14114;
wire      [7:0] n14115;
wire      [7:0] n14116;
wire      [7:0] n14117;
wire      [7:0] n14118;
wire      [7:0] n14119;
wire      [7:0] n1412;
wire      [7:0] n14120;
wire      [7:0] n14121;
wire      [7:0] n14122;
wire      [7:0] n14123;
wire      [7:0] n14124;
wire      [7:0] n14125;
wire      [7:0] n14126;
wire      [7:0] n14127;
wire      [7:0] n14128;
wire      [7:0] n14129;
wire            n1413;
wire      [7:0] n14130;
wire      [7:0] n14131;
wire      [7:0] n14132;
wire      [7:0] n14133;
wire      [7:0] n14134;
wire      [7:0] n14135;
wire      [7:0] n14136;
wire      [7:0] n14137;
wire      [7:0] n14138;
wire            n14139;
wire      [7:0] n1414;
wire      [7:0] n14140;
wire            n14141;
wire      [7:0] n14142;
wire            n14143;
wire      [7:0] n14144;
wire            n14145;
wire      [7:0] n14146;
wire            n14147;
wire      [7:0] n14148;
wire            n14149;
wire            n1415;
wire      [7:0] n14150;
wire            n14151;
wire      [7:0] n14152;
wire            n14153;
wire      [7:0] n14154;
wire            n14155;
wire      [7:0] n14156;
wire            n14157;
wire      [7:0] n14158;
wire            n14159;
wire      [7:0] n1416;
wire      [7:0] n14160;
wire            n14161;
wire      [7:0] n14162;
wire            n14163;
wire      [7:0] n14164;
wire            n14165;
wire      [7:0] n14166;
wire            n14167;
wire      [7:0] n14168;
wire            n14169;
wire            n1417;
wire      [7:0] n14170;
wire            n14171;
wire      [7:0] n14172;
wire            n14173;
wire      [7:0] n14174;
wire            n14175;
wire      [7:0] n14176;
wire            n14177;
wire      [7:0] n14178;
wire            n14179;
wire      [7:0] n1418;
wire      [7:0] n14180;
wire            n14181;
wire      [7:0] n14182;
wire            n14183;
wire      [7:0] n14184;
wire            n14185;
wire      [7:0] n14186;
wire            n14187;
wire      [7:0] n14188;
wire            n14189;
wire            n1419;
wire      [7:0] n14190;
wire            n14191;
wire      [7:0] n14192;
wire            n14193;
wire      [7:0] n14194;
wire            n14195;
wire      [7:0] n14196;
wire            n14197;
wire      [7:0] n14198;
wire            n14199;
wire      [7:0] n1420;
wire      [7:0] n14200;
wire            n14201;
wire      [7:0] n14202;
wire            n14203;
wire      [7:0] n14204;
wire            n14205;
wire      [7:0] n14206;
wire            n14207;
wire      [7:0] n14208;
wire            n14209;
wire            n1421;
wire      [7:0] n14210;
wire            n14211;
wire      [7:0] n14212;
wire            n14213;
wire      [7:0] n14214;
wire            n14215;
wire      [7:0] n14216;
wire            n14217;
wire      [7:0] n14218;
wire            n14219;
wire      [7:0] n1422;
wire      [7:0] n14220;
wire            n14221;
wire      [7:0] n14222;
wire            n14223;
wire      [7:0] n14224;
wire            n14225;
wire      [7:0] n14226;
wire            n14227;
wire      [7:0] n14228;
wire            n14229;
wire            n1423;
wire      [7:0] n14230;
wire            n14231;
wire      [7:0] n14232;
wire            n14233;
wire      [7:0] n14234;
wire            n14235;
wire      [7:0] n14236;
wire            n14237;
wire      [7:0] n14238;
wire            n14239;
wire      [7:0] n1424;
wire      [7:0] n14240;
wire            n14241;
wire      [7:0] n14242;
wire            n14243;
wire      [7:0] n14244;
wire            n14245;
wire      [7:0] n14246;
wire            n14247;
wire      [7:0] n14248;
wire            n14249;
wire            n1425;
wire      [7:0] n14250;
wire            n14251;
wire      [7:0] n14252;
wire            n14253;
wire      [7:0] n14254;
wire            n14255;
wire      [7:0] n14256;
wire            n14257;
wire      [7:0] n14258;
wire            n14259;
wire      [7:0] n1426;
wire      [7:0] n14260;
wire            n14261;
wire      [7:0] n14262;
wire            n14263;
wire      [7:0] n14264;
wire            n14265;
wire      [7:0] n14266;
wire            n14267;
wire      [7:0] n14268;
wire            n14269;
wire            n1427;
wire      [7:0] n14270;
wire            n14271;
wire      [7:0] n14272;
wire            n14273;
wire      [7:0] n14274;
wire            n14275;
wire      [7:0] n14276;
wire            n14277;
wire      [7:0] n14278;
wire            n14279;
wire      [7:0] n1428;
wire      [7:0] n14280;
wire            n14281;
wire      [7:0] n14282;
wire            n14283;
wire      [7:0] n14284;
wire            n14285;
wire      [7:0] n14286;
wire            n14287;
wire      [7:0] n14288;
wire            n14289;
wire            n1429;
wire      [7:0] n14290;
wire            n14291;
wire      [7:0] n14292;
wire            n14293;
wire      [7:0] n14294;
wire            n14295;
wire      [7:0] n14296;
wire            n14297;
wire      [7:0] n14298;
wire            n14299;
wire            n143;
wire      [7:0] n1430;
wire      [7:0] n14300;
wire            n14301;
wire      [7:0] n14302;
wire            n14303;
wire      [7:0] n14304;
wire            n14305;
wire      [7:0] n14306;
wire            n14307;
wire      [7:0] n14308;
wire            n14309;
wire            n1431;
wire      [7:0] n14310;
wire            n14311;
wire      [7:0] n14312;
wire            n14313;
wire      [7:0] n14314;
wire            n14315;
wire      [7:0] n14316;
wire            n14317;
wire      [7:0] n14318;
wire            n14319;
wire      [7:0] n1432;
wire      [7:0] n14320;
wire            n14321;
wire      [7:0] n14322;
wire            n14323;
wire      [7:0] n14324;
wire            n14325;
wire      [7:0] n14326;
wire            n14327;
wire      [7:0] n14328;
wire            n14329;
wire            n1433;
wire      [7:0] n14330;
wire            n14331;
wire      [7:0] n14332;
wire            n14333;
wire      [7:0] n14334;
wire            n14335;
wire      [7:0] n14336;
wire            n14337;
wire      [7:0] n14338;
wire            n14339;
wire      [7:0] n1434;
wire      [7:0] n14340;
wire            n14341;
wire      [7:0] n14342;
wire            n14343;
wire      [7:0] n14344;
wire            n14345;
wire      [7:0] n14346;
wire            n14347;
wire      [7:0] n14348;
wire            n14349;
wire            n1435;
wire      [7:0] n14350;
wire            n14351;
wire      [7:0] n14352;
wire            n14353;
wire      [7:0] n14354;
wire            n14355;
wire      [7:0] n14356;
wire            n14357;
wire      [7:0] n14358;
wire            n14359;
wire      [7:0] n1436;
wire      [7:0] n14360;
wire            n14361;
wire      [7:0] n14362;
wire            n14363;
wire      [7:0] n14364;
wire            n14365;
wire      [7:0] n14366;
wire            n14367;
wire      [7:0] n14368;
wire            n14369;
wire            n1437;
wire      [7:0] n14370;
wire            n14371;
wire      [7:0] n14372;
wire            n14373;
wire      [7:0] n14374;
wire            n14375;
wire      [7:0] n14376;
wire            n14377;
wire      [7:0] n14378;
wire            n14379;
wire      [7:0] n1438;
wire      [7:0] n14380;
wire            n14381;
wire      [7:0] n14382;
wire            n14383;
wire      [7:0] n14384;
wire            n14385;
wire      [7:0] n14386;
wire            n14387;
wire      [7:0] n14388;
wire            n14389;
wire            n1439;
wire      [7:0] n14390;
wire            n14391;
wire      [7:0] n14392;
wire            n14393;
wire      [7:0] n14394;
wire            n14395;
wire      [7:0] n14396;
wire            n14397;
wire      [7:0] n14398;
wire            n14399;
wire      [7:0] n1440;
wire      [7:0] n14400;
wire            n14401;
wire      [7:0] n14402;
wire            n14403;
wire      [7:0] n14404;
wire            n14405;
wire      [7:0] n14406;
wire            n14407;
wire      [7:0] n14408;
wire            n14409;
wire            n1441;
wire      [7:0] n14410;
wire            n14411;
wire      [7:0] n14412;
wire            n14413;
wire      [7:0] n14414;
wire            n14415;
wire      [7:0] n14416;
wire            n14417;
wire      [7:0] n14418;
wire            n14419;
wire      [7:0] n1442;
wire      [7:0] n14420;
wire            n14421;
wire      [7:0] n14422;
wire            n14423;
wire      [7:0] n14424;
wire            n14425;
wire      [7:0] n14426;
wire            n14427;
wire      [7:0] n14428;
wire            n14429;
wire            n1443;
wire      [7:0] n14430;
wire            n14431;
wire      [7:0] n14432;
wire            n14433;
wire      [7:0] n14434;
wire            n14435;
wire      [7:0] n14436;
wire            n14437;
wire      [7:0] n14438;
wire            n14439;
wire      [7:0] n1444;
wire      [7:0] n14440;
wire            n14441;
wire      [7:0] n14442;
wire            n14443;
wire      [7:0] n14444;
wire            n14445;
wire      [7:0] n14446;
wire            n14447;
wire      [7:0] n14448;
wire            n14449;
wire            n1445;
wire      [7:0] n14450;
wire            n14451;
wire      [7:0] n14452;
wire            n14453;
wire      [7:0] n14454;
wire            n14455;
wire      [7:0] n14456;
wire            n14457;
wire      [7:0] n14458;
wire            n14459;
wire      [7:0] n1446;
wire      [7:0] n14460;
wire            n14461;
wire      [7:0] n14462;
wire            n14463;
wire      [7:0] n14464;
wire            n14465;
wire      [7:0] n14466;
wire            n14467;
wire      [7:0] n14468;
wire            n14469;
wire            n1447;
wire      [7:0] n14470;
wire            n14471;
wire      [7:0] n14472;
wire            n14473;
wire      [7:0] n14474;
wire            n14475;
wire      [7:0] n14476;
wire            n14477;
wire      [7:0] n14478;
wire            n14479;
wire      [7:0] n1448;
wire      [7:0] n14480;
wire            n14481;
wire      [7:0] n14482;
wire            n14483;
wire      [7:0] n14484;
wire            n14485;
wire      [7:0] n14486;
wire            n14487;
wire      [7:0] n14488;
wire            n14489;
wire            n1449;
wire      [7:0] n14490;
wire            n14491;
wire      [7:0] n14492;
wire            n14493;
wire      [7:0] n14494;
wire            n14495;
wire      [7:0] n14496;
wire            n14497;
wire      [7:0] n14498;
wire            n14499;
wire      [7:0] n145;
wire      [7:0] n1450;
wire      [7:0] n14500;
wire            n14501;
wire      [7:0] n14502;
wire            n14503;
wire      [7:0] n14504;
wire            n14505;
wire      [7:0] n14506;
wire            n14507;
wire      [7:0] n14508;
wire            n14509;
wire            n1451;
wire      [7:0] n14510;
wire            n14511;
wire      [7:0] n14512;
wire            n14513;
wire      [7:0] n14514;
wire            n14515;
wire      [7:0] n14516;
wire            n14517;
wire      [7:0] n14518;
wire            n14519;
wire      [7:0] n1452;
wire      [7:0] n14520;
wire            n14521;
wire      [7:0] n14522;
wire            n14523;
wire      [7:0] n14524;
wire            n14525;
wire      [7:0] n14526;
wire            n14527;
wire      [7:0] n14528;
wire            n14529;
wire            n1453;
wire      [7:0] n14530;
wire            n14531;
wire      [7:0] n14532;
wire            n14533;
wire      [7:0] n14534;
wire            n14535;
wire      [7:0] n14536;
wire            n14537;
wire      [7:0] n14538;
wire            n14539;
wire      [7:0] n1454;
wire      [7:0] n14540;
wire            n14541;
wire      [7:0] n14542;
wire            n14543;
wire      [7:0] n14544;
wire            n14545;
wire      [7:0] n14546;
wire            n14547;
wire      [7:0] n14548;
wire            n14549;
wire            n1455;
wire      [7:0] n14550;
wire            n14551;
wire      [7:0] n14552;
wire            n14553;
wire      [7:0] n14554;
wire            n14555;
wire      [7:0] n14556;
wire            n14557;
wire      [7:0] n14558;
wire            n14559;
wire      [7:0] n1456;
wire      [7:0] n14560;
wire            n14561;
wire      [7:0] n14562;
wire            n14563;
wire      [7:0] n14564;
wire            n14565;
wire      [7:0] n14566;
wire            n14567;
wire      [7:0] n14568;
wire            n14569;
wire            n1457;
wire      [7:0] n14570;
wire            n14571;
wire      [7:0] n14572;
wire            n14573;
wire      [7:0] n14574;
wire            n14575;
wire      [7:0] n14576;
wire            n14577;
wire      [7:0] n14578;
wire            n14579;
wire      [7:0] n1458;
wire      [7:0] n14580;
wire            n14581;
wire      [7:0] n14582;
wire            n14583;
wire      [7:0] n14584;
wire            n14585;
wire      [7:0] n14586;
wire            n14587;
wire      [7:0] n14588;
wire            n14589;
wire            n1459;
wire      [7:0] n14590;
wire            n14591;
wire      [7:0] n14592;
wire            n14593;
wire      [7:0] n14594;
wire            n14595;
wire      [7:0] n14596;
wire            n14597;
wire      [7:0] n14598;
wire            n14599;
wire      [7:0] n1460;
wire      [7:0] n14600;
wire            n14601;
wire      [7:0] n14602;
wire            n14603;
wire      [7:0] n14604;
wire            n14605;
wire      [7:0] n14606;
wire            n14607;
wire      [7:0] n14608;
wire            n14609;
wire            n1461;
wire      [7:0] n14610;
wire            n14611;
wire      [7:0] n14612;
wire            n14613;
wire      [7:0] n14614;
wire            n14615;
wire      [7:0] n14616;
wire            n14617;
wire      [7:0] n14618;
wire            n14619;
wire      [7:0] n1462;
wire      [7:0] n14620;
wire            n14621;
wire      [7:0] n14622;
wire            n14623;
wire      [7:0] n14624;
wire            n14625;
wire      [7:0] n14626;
wire            n14627;
wire      [7:0] n14628;
wire            n14629;
wire            n1463;
wire      [7:0] n14630;
wire            n14631;
wire      [7:0] n14632;
wire            n14633;
wire      [7:0] n14634;
wire            n14635;
wire      [7:0] n14636;
wire            n14637;
wire      [7:0] n14638;
wire            n14639;
wire      [7:0] n1464;
wire      [7:0] n14640;
wire            n14641;
wire      [7:0] n14642;
wire            n14643;
wire      [7:0] n14644;
wire            n14645;
wire      [7:0] n14646;
wire            n14647;
wire      [7:0] n14648;
wire            n14649;
wire            n1465;
wire      [7:0] n14650;
wire      [7:0] n14651;
wire      [7:0] n14652;
wire      [7:0] n14653;
wire      [7:0] n14654;
wire      [7:0] n14655;
wire      [7:0] n14656;
wire      [7:0] n14657;
wire      [7:0] n14658;
wire      [7:0] n14659;
wire      [7:0] n1466;
wire      [7:0] n14660;
wire      [7:0] n14661;
wire      [7:0] n14662;
wire      [7:0] n14663;
wire      [7:0] n14664;
wire      [7:0] n14665;
wire      [7:0] n14666;
wire      [7:0] n14667;
wire      [7:0] n14668;
wire      [7:0] n14669;
wire            n1467;
wire      [7:0] n14670;
wire      [7:0] n14671;
wire      [7:0] n14672;
wire      [7:0] n14673;
wire      [7:0] n14674;
wire      [7:0] n14675;
wire      [7:0] n14676;
wire      [7:0] n14677;
wire      [7:0] n14678;
wire      [7:0] n14679;
wire      [7:0] n1468;
wire      [7:0] n14680;
wire      [7:0] n14681;
wire      [7:0] n14682;
wire      [7:0] n14683;
wire      [7:0] n14684;
wire      [7:0] n14685;
wire      [7:0] n14686;
wire      [7:0] n14687;
wire      [7:0] n14688;
wire      [7:0] n14689;
wire            n1469;
wire      [7:0] n14690;
wire      [7:0] n14691;
wire      [7:0] n14692;
wire      [7:0] n14693;
wire      [7:0] n14694;
wire      [7:0] n14695;
wire      [7:0] n14696;
wire      [7:0] n14697;
wire      [7:0] n14698;
wire      [7:0] n14699;
wire            n147;
wire      [7:0] n1470;
wire      [7:0] n14700;
wire      [7:0] n14701;
wire      [7:0] n14702;
wire      [7:0] n14703;
wire      [7:0] n14704;
wire      [7:0] n14705;
wire      [7:0] n14706;
wire      [7:0] n14707;
wire      [7:0] n14708;
wire      [7:0] n14709;
wire            n1471;
wire      [7:0] n14710;
wire      [7:0] n14711;
wire      [7:0] n14712;
wire      [7:0] n14713;
wire      [7:0] n14714;
wire      [7:0] n14715;
wire      [7:0] n14716;
wire      [7:0] n14717;
wire      [7:0] n14718;
wire      [7:0] n14719;
wire      [7:0] n1472;
wire      [7:0] n14720;
wire      [7:0] n14721;
wire      [7:0] n14722;
wire      [7:0] n14723;
wire      [7:0] n14724;
wire      [7:0] n14725;
wire      [7:0] n14726;
wire      [7:0] n14727;
wire      [7:0] n14728;
wire      [7:0] n14729;
wire            n1473;
wire      [7:0] n14730;
wire      [7:0] n14731;
wire      [7:0] n14732;
wire      [7:0] n14733;
wire      [7:0] n14734;
wire      [7:0] n14735;
wire      [7:0] n14736;
wire      [7:0] n14737;
wire      [7:0] n14738;
wire      [7:0] n14739;
wire      [7:0] n1474;
wire      [7:0] n14740;
wire      [7:0] n14741;
wire      [7:0] n14742;
wire      [7:0] n14743;
wire      [7:0] n14744;
wire      [7:0] n14745;
wire      [7:0] n14746;
wire      [7:0] n14747;
wire      [7:0] n14748;
wire      [7:0] n14749;
wire            n1475;
wire      [7:0] n14750;
wire      [7:0] n14751;
wire      [7:0] n14752;
wire      [7:0] n14753;
wire      [7:0] n14754;
wire      [7:0] n14755;
wire      [7:0] n14756;
wire      [7:0] n14757;
wire      [7:0] n14758;
wire      [7:0] n14759;
wire      [7:0] n1476;
wire      [7:0] n14760;
wire      [7:0] n14761;
wire      [7:0] n14762;
wire      [7:0] n14763;
wire      [7:0] n14764;
wire      [7:0] n14765;
wire      [7:0] n14766;
wire      [7:0] n14767;
wire      [7:0] n14768;
wire      [7:0] n14769;
wire            n1477;
wire      [7:0] n14770;
wire      [7:0] n14771;
wire      [7:0] n14772;
wire      [7:0] n14773;
wire      [7:0] n14774;
wire      [7:0] n14775;
wire      [7:0] n14776;
wire      [7:0] n14777;
wire      [7:0] n14778;
wire      [7:0] n14779;
wire      [7:0] n1478;
wire      [7:0] n14780;
wire      [7:0] n14781;
wire      [7:0] n14782;
wire      [7:0] n14783;
wire      [7:0] n14784;
wire      [7:0] n14785;
wire      [7:0] n14786;
wire      [7:0] n14787;
wire      [7:0] n14788;
wire      [7:0] n14789;
wire            n1479;
wire      [7:0] n14790;
wire      [7:0] n14791;
wire      [7:0] n14792;
wire      [7:0] n14793;
wire      [7:0] n14794;
wire      [7:0] n14795;
wire      [7:0] n14796;
wire      [7:0] n14797;
wire      [7:0] n14798;
wire      [7:0] n14799;
wire      [7:0] n1480;
wire      [7:0] n14800;
wire      [7:0] n14801;
wire      [7:0] n14802;
wire      [7:0] n14803;
wire      [7:0] n14804;
wire      [7:0] n14805;
wire      [7:0] n14806;
wire      [7:0] n14807;
wire      [7:0] n14808;
wire      [7:0] n14809;
wire            n1481;
wire      [7:0] n14810;
wire      [7:0] n14811;
wire      [7:0] n14812;
wire      [7:0] n14813;
wire      [7:0] n14814;
wire      [7:0] n14815;
wire      [7:0] n14816;
wire      [7:0] n14817;
wire      [7:0] n14818;
wire      [7:0] n14819;
wire      [7:0] n1482;
wire      [7:0] n14820;
wire      [7:0] n14821;
wire      [7:0] n14822;
wire      [7:0] n14823;
wire      [7:0] n14824;
wire      [7:0] n14825;
wire      [7:0] n14826;
wire      [7:0] n14827;
wire      [7:0] n14828;
wire      [7:0] n14829;
wire            n1483;
wire      [7:0] n14830;
wire      [7:0] n14831;
wire      [7:0] n14832;
wire      [7:0] n14833;
wire      [7:0] n14834;
wire      [7:0] n14835;
wire      [7:0] n14836;
wire      [7:0] n14837;
wire      [7:0] n14838;
wire      [7:0] n14839;
wire      [7:0] n1484;
wire      [7:0] n14840;
wire      [7:0] n14841;
wire      [7:0] n14842;
wire      [7:0] n14843;
wire      [7:0] n14844;
wire      [7:0] n14845;
wire      [7:0] n14846;
wire      [7:0] n14847;
wire      [7:0] n14848;
wire      [7:0] n14849;
wire            n1485;
wire      [7:0] n14850;
wire      [7:0] n14851;
wire      [7:0] n14852;
wire      [7:0] n14853;
wire      [7:0] n14854;
wire      [7:0] n14855;
wire      [7:0] n14856;
wire      [7:0] n14857;
wire      [7:0] n14858;
wire      [7:0] n14859;
wire      [7:0] n1486;
wire      [7:0] n14860;
wire      [7:0] n14861;
wire      [7:0] n14862;
wire      [7:0] n14863;
wire      [7:0] n14864;
wire      [7:0] n14865;
wire      [7:0] n14866;
wire      [7:0] n14867;
wire      [7:0] n14868;
wire      [7:0] n14869;
wire            n1487;
wire      [7:0] n14870;
wire      [7:0] n14871;
wire      [7:0] n14872;
wire      [7:0] n14873;
wire      [7:0] n14874;
wire      [7:0] n14875;
wire      [7:0] n14876;
wire      [7:0] n14877;
wire      [7:0] n14878;
wire      [7:0] n14879;
wire      [7:0] n1488;
wire      [7:0] n14880;
wire      [7:0] n14881;
wire      [7:0] n14882;
wire      [7:0] n14883;
wire      [7:0] n14884;
wire      [7:0] n14885;
wire      [7:0] n14886;
wire      [7:0] n14887;
wire      [7:0] n14888;
wire      [7:0] n14889;
wire            n1489;
wire      [7:0] n14890;
wire      [7:0] n14891;
wire      [7:0] n14892;
wire      [7:0] n14893;
wire      [7:0] n14894;
wire      [7:0] n14895;
wire      [7:0] n14896;
wire      [7:0] n14897;
wire      [7:0] n14898;
wire      [7:0] n14899;
wire      [7:0] n149;
wire      [7:0] n1490;
wire      [7:0] n14900;
wire      [7:0] n14901;
wire      [7:0] n14902;
wire      [7:0] n14903;
wire      [7:0] n14904;
wire      [7:0] n14905;
wire      [7:0] n14906;
wire      [7:0] n14907;
wire            n14908;
wire      [7:0] n14909;
wire            n1491;
wire            n14910;
wire      [7:0] n14911;
wire            n14912;
wire      [7:0] n14913;
wire            n14914;
wire      [7:0] n14915;
wire            n14916;
wire      [7:0] n14917;
wire            n14918;
wire      [7:0] n14919;
wire      [7:0] n1492;
wire            n14920;
wire      [7:0] n14921;
wire            n14922;
wire      [7:0] n14923;
wire            n14924;
wire      [7:0] n14925;
wire            n14926;
wire      [7:0] n14927;
wire            n14928;
wire      [7:0] n14929;
wire            n1493;
wire            n14930;
wire      [7:0] n14931;
wire            n14932;
wire      [7:0] n14933;
wire            n14934;
wire      [7:0] n14935;
wire            n14936;
wire      [7:0] n14937;
wire            n14938;
wire      [7:0] n14939;
wire      [7:0] n1494;
wire            n14940;
wire      [7:0] n14941;
wire            n14942;
wire      [7:0] n14943;
wire            n14944;
wire      [7:0] n14945;
wire            n14946;
wire      [7:0] n14947;
wire            n14948;
wire      [7:0] n14949;
wire            n1495;
wire            n14950;
wire      [7:0] n14951;
wire            n14952;
wire      [7:0] n14953;
wire            n14954;
wire      [7:0] n14955;
wire            n14956;
wire      [7:0] n14957;
wire            n14958;
wire      [7:0] n14959;
wire      [7:0] n1496;
wire            n14960;
wire      [7:0] n14961;
wire            n14962;
wire      [7:0] n14963;
wire            n14964;
wire      [7:0] n14965;
wire            n14966;
wire      [7:0] n14967;
wire            n14968;
wire      [7:0] n14969;
wire            n1497;
wire            n14970;
wire      [7:0] n14971;
wire            n14972;
wire      [7:0] n14973;
wire            n14974;
wire      [7:0] n14975;
wire            n14976;
wire      [7:0] n14977;
wire            n14978;
wire      [7:0] n14979;
wire      [7:0] n1498;
wire            n14980;
wire      [7:0] n14981;
wire            n14982;
wire      [7:0] n14983;
wire            n14984;
wire      [7:0] n14985;
wire            n14986;
wire      [7:0] n14987;
wire            n14988;
wire      [7:0] n14989;
wire            n1499;
wire            n14990;
wire      [7:0] n14991;
wire            n14992;
wire      [7:0] n14993;
wire            n14994;
wire      [7:0] n14995;
wire            n14996;
wire      [7:0] n14997;
wire            n14998;
wire      [7:0] n14999;
wire      [7:0] n1500;
wire            n15000;
wire      [7:0] n15001;
wire            n15002;
wire      [7:0] n15003;
wire            n15004;
wire      [7:0] n15005;
wire            n15006;
wire      [7:0] n15007;
wire            n15008;
wire      [7:0] n15009;
wire            n1501;
wire            n15010;
wire      [7:0] n15011;
wire            n15012;
wire      [7:0] n15013;
wire            n15014;
wire      [7:0] n15015;
wire            n15016;
wire      [7:0] n15017;
wire            n15018;
wire      [7:0] n15019;
wire      [7:0] n1502;
wire            n15020;
wire      [7:0] n15021;
wire            n15022;
wire      [7:0] n15023;
wire            n15024;
wire      [7:0] n15025;
wire            n15026;
wire      [7:0] n15027;
wire            n15028;
wire      [7:0] n15029;
wire            n1503;
wire            n15030;
wire      [7:0] n15031;
wire            n15032;
wire      [7:0] n15033;
wire            n15034;
wire      [7:0] n15035;
wire            n15036;
wire      [7:0] n15037;
wire            n15038;
wire      [7:0] n15039;
wire      [7:0] n1504;
wire            n15040;
wire      [7:0] n15041;
wire            n15042;
wire      [7:0] n15043;
wire            n15044;
wire      [7:0] n15045;
wire            n15046;
wire      [7:0] n15047;
wire            n15048;
wire      [7:0] n15049;
wire            n1505;
wire            n15050;
wire      [7:0] n15051;
wire            n15052;
wire      [7:0] n15053;
wire            n15054;
wire      [7:0] n15055;
wire            n15056;
wire      [7:0] n15057;
wire            n15058;
wire      [7:0] n15059;
wire      [7:0] n1506;
wire            n15060;
wire      [7:0] n15061;
wire            n15062;
wire      [7:0] n15063;
wire            n15064;
wire      [7:0] n15065;
wire            n15066;
wire      [7:0] n15067;
wire            n15068;
wire      [7:0] n15069;
wire            n1507;
wire            n15070;
wire      [7:0] n15071;
wire            n15072;
wire      [7:0] n15073;
wire            n15074;
wire      [7:0] n15075;
wire            n15076;
wire      [7:0] n15077;
wire            n15078;
wire      [7:0] n15079;
wire      [7:0] n1508;
wire            n15080;
wire      [7:0] n15081;
wire            n15082;
wire      [7:0] n15083;
wire            n15084;
wire      [7:0] n15085;
wire            n15086;
wire      [7:0] n15087;
wire            n15088;
wire      [7:0] n15089;
wire            n1509;
wire            n15090;
wire      [7:0] n15091;
wire            n15092;
wire      [7:0] n15093;
wire            n15094;
wire      [7:0] n15095;
wire            n15096;
wire      [7:0] n15097;
wire            n15098;
wire      [7:0] n15099;
wire            n151;
wire      [7:0] n1510;
wire            n15100;
wire      [7:0] n15101;
wire            n15102;
wire      [7:0] n15103;
wire            n15104;
wire      [7:0] n15105;
wire            n15106;
wire      [7:0] n15107;
wire            n15108;
wire      [7:0] n15109;
wire            n1511;
wire            n15110;
wire      [7:0] n15111;
wire            n15112;
wire      [7:0] n15113;
wire            n15114;
wire      [7:0] n15115;
wire            n15116;
wire      [7:0] n15117;
wire            n15118;
wire      [7:0] n15119;
wire      [7:0] n1512;
wire            n15120;
wire      [7:0] n15121;
wire            n15122;
wire      [7:0] n15123;
wire            n15124;
wire      [7:0] n15125;
wire            n15126;
wire      [7:0] n15127;
wire            n15128;
wire      [7:0] n15129;
wire            n1513;
wire            n15130;
wire      [7:0] n15131;
wire            n15132;
wire      [7:0] n15133;
wire            n15134;
wire      [7:0] n15135;
wire            n15136;
wire      [7:0] n15137;
wire            n15138;
wire      [7:0] n15139;
wire      [7:0] n1514;
wire            n15140;
wire      [7:0] n15141;
wire            n15142;
wire      [7:0] n15143;
wire            n15144;
wire      [7:0] n15145;
wire            n15146;
wire      [7:0] n15147;
wire            n15148;
wire      [7:0] n15149;
wire            n1515;
wire            n15150;
wire      [7:0] n15151;
wire            n15152;
wire      [7:0] n15153;
wire            n15154;
wire      [7:0] n15155;
wire            n15156;
wire      [7:0] n15157;
wire            n15158;
wire      [7:0] n15159;
wire      [7:0] n1516;
wire            n15160;
wire      [7:0] n15161;
wire            n15162;
wire      [7:0] n15163;
wire            n15164;
wire      [7:0] n15165;
wire            n15166;
wire      [7:0] n15167;
wire            n15168;
wire      [7:0] n15169;
wire            n1517;
wire            n15170;
wire      [7:0] n15171;
wire            n15172;
wire      [7:0] n15173;
wire            n15174;
wire      [7:0] n15175;
wire            n15176;
wire      [7:0] n15177;
wire            n15178;
wire      [7:0] n15179;
wire      [7:0] n1518;
wire            n15180;
wire      [7:0] n15181;
wire            n15182;
wire      [7:0] n15183;
wire            n15184;
wire      [7:0] n15185;
wire            n15186;
wire      [7:0] n15187;
wire            n15188;
wire      [7:0] n15189;
wire            n1519;
wire            n15190;
wire      [7:0] n15191;
wire            n15192;
wire      [7:0] n15193;
wire            n15194;
wire      [7:0] n15195;
wire            n15196;
wire      [7:0] n15197;
wire            n15198;
wire      [7:0] n15199;
wire      [7:0] n1520;
wire            n15200;
wire      [7:0] n15201;
wire            n15202;
wire      [7:0] n15203;
wire            n15204;
wire      [7:0] n15205;
wire            n15206;
wire      [7:0] n15207;
wire            n15208;
wire      [7:0] n15209;
wire            n1521;
wire            n15210;
wire      [7:0] n15211;
wire            n15212;
wire      [7:0] n15213;
wire            n15214;
wire      [7:0] n15215;
wire            n15216;
wire      [7:0] n15217;
wire            n15218;
wire      [7:0] n15219;
wire      [7:0] n1522;
wire            n15220;
wire      [7:0] n15221;
wire            n15222;
wire      [7:0] n15223;
wire            n15224;
wire      [7:0] n15225;
wire            n15226;
wire      [7:0] n15227;
wire            n15228;
wire      [7:0] n15229;
wire            n1523;
wire            n15230;
wire      [7:0] n15231;
wire            n15232;
wire      [7:0] n15233;
wire            n15234;
wire      [7:0] n15235;
wire            n15236;
wire      [7:0] n15237;
wire            n15238;
wire      [7:0] n15239;
wire      [7:0] n1524;
wire            n15240;
wire      [7:0] n15241;
wire            n15242;
wire      [7:0] n15243;
wire            n15244;
wire      [7:0] n15245;
wire            n15246;
wire      [7:0] n15247;
wire            n15248;
wire      [7:0] n15249;
wire            n1525;
wire            n15250;
wire      [7:0] n15251;
wire            n15252;
wire      [7:0] n15253;
wire            n15254;
wire      [7:0] n15255;
wire            n15256;
wire      [7:0] n15257;
wire            n15258;
wire      [7:0] n15259;
wire      [7:0] n1526;
wire            n15260;
wire      [7:0] n15261;
wire            n15262;
wire      [7:0] n15263;
wire            n15264;
wire      [7:0] n15265;
wire            n15266;
wire      [7:0] n15267;
wire            n15268;
wire      [7:0] n15269;
wire            n1527;
wire            n15270;
wire      [7:0] n15271;
wire            n15272;
wire      [7:0] n15273;
wire            n15274;
wire      [7:0] n15275;
wire            n15276;
wire      [7:0] n15277;
wire            n15278;
wire      [7:0] n15279;
wire      [7:0] n1528;
wire            n15280;
wire      [7:0] n15281;
wire            n15282;
wire      [7:0] n15283;
wire            n15284;
wire      [7:0] n15285;
wire            n15286;
wire      [7:0] n15287;
wire            n15288;
wire      [7:0] n15289;
wire            n1529;
wire            n15290;
wire      [7:0] n15291;
wire            n15292;
wire      [7:0] n15293;
wire            n15294;
wire      [7:0] n15295;
wire            n15296;
wire      [7:0] n15297;
wire            n15298;
wire      [7:0] n15299;
wire      [7:0] n153;
wire      [7:0] n1530;
wire            n15300;
wire      [7:0] n15301;
wire            n15302;
wire      [7:0] n15303;
wire            n15304;
wire      [7:0] n15305;
wire            n15306;
wire      [7:0] n15307;
wire            n15308;
wire      [7:0] n15309;
wire            n1531;
wire            n15310;
wire      [7:0] n15311;
wire            n15312;
wire      [7:0] n15313;
wire            n15314;
wire      [7:0] n15315;
wire            n15316;
wire      [7:0] n15317;
wire            n15318;
wire      [7:0] n15319;
wire      [7:0] n1532;
wire            n15320;
wire      [7:0] n15321;
wire            n15322;
wire      [7:0] n15323;
wire            n15324;
wire      [7:0] n15325;
wire            n15326;
wire      [7:0] n15327;
wire            n15328;
wire      [7:0] n15329;
wire            n1533;
wire            n15330;
wire      [7:0] n15331;
wire            n15332;
wire      [7:0] n15333;
wire            n15334;
wire      [7:0] n15335;
wire            n15336;
wire      [7:0] n15337;
wire            n15338;
wire      [7:0] n15339;
wire      [7:0] n1534;
wire            n15340;
wire      [7:0] n15341;
wire            n15342;
wire      [7:0] n15343;
wire            n15344;
wire      [7:0] n15345;
wire            n15346;
wire      [7:0] n15347;
wire            n15348;
wire      [7:0] n15349;
wire            n1535;
wire            n15350;
wire      [7:0] n15351;
wire            n15352;
wire      [7:0] n15353;
wire            n15354;
wire      [7:0] n15355;
wire            n15356;
wire      [7:0] n15357;
wire            n15358;
wire      [7:0] n15359;
wire      [7:0] n1536;
wire            n15360;
wire      [7:0] n15361;
wire            n15362;
wire      [7:0] n15363;
wire            n15364;
wire      [7:0] n15365;
wire            n15366;
wire      [7:0] n15367;
wire            n15368;
wire      [7:0] n15369;
wire            n1537;
wire            n15370;
wire      [7:0] n15371;
wire            n15372;
wire      [7:0] n15373;
wire            n15374;
wire      [7:0] n15375;
wire            n15376;
wire      [7:0] n15377;
wire            n15378;
wire      [7:0] n15379;
wire      [7:0] n1538;
wire            n15380;
wire      [7:0] n15381;
wire            n15382;
wire      [7:0] n15383;
wire            n15384;
wire      [7:0] n15385;
wire            n15386;
wire      [7:0] n15387;
wire            n15388;
wire      [7:0] n15389;
wire      [7:0] n1539;
wire            n15390;
wire      [7:0] n15391;
wire            n15392;
wire      [7:0] n15393;
wire            n15394;
wire      [7:0] n15395;
wire            n15396;
wire      [7:0] n15397;
wire            n15398;
wire      [7:0] n15399;
wire            n154;
wire      [7:0] n1540;
wire            n15400;
wire      [7:0] n15401;
wire            n15402;
wire      [7:0] n15403;
wire            n15404;
wire      [7:0] n15405;
wire            n15406;
wire      [7:0] n15407;
wire            n15408;
wire      [7:0] n15409;
wire      [7:0] n1541;
wire            n15410;
wire      [7:0] n15411;
wire            n15412;
wire      [7:0] n15413;
wire            n15414;
wire      [7:0] n15415;
wire            n15416;
wire      [7:0] n15417;
wire            n15418;
wire      [7:0] n15419;
wire      [7:0] n1542;
wire      [7:0] n15420;
wire      [7:0] n15421;
wire      [7:0] n15422;
wire      [7:0] n15423;
wire      [7:0] n15424;
wire      [7:0] n15425;
wire      [7:0] n15426;
wire      [7:0] n15427;
wire      [7:0] n15428;
wire      [7:0] n15429;
wire      [7:0] n1543;
wire      [7:0] n15430;
wire      [7:0] n15431;
wire      [7:0] n15432;
wire      [7:0] n15433;
wire      [7:0] n15434;
wire      [7:0] n15435;
wire      [7:0] n15436;
wire      [7:0] n15437;
wire      [7:0] n15438;
wire      [7:0] n15439;
wire      [7:0] n1544;
wire      [7:0] n15440;
wire      [7:0] n15441;
wire      [7:0] n15442;
wire      [7:0] n15443;
wire      [7:0] n15444;
wire      [7:0] n15445;
wire      [7:0] n15446;
wire      [7:0] n15447;
wire      [7:0] n15448;
wire      [7:0] n15449;
wire      [7:0] n1545;
wire      [7:0] n15450;
wire      [7:0] n15451;
wire      [7:0] n15452;
wire      [7:0] n15453;
wire      [7:0] n15454;
wire      [7:0] n15455;
wire      [7:0] n15456;
wire      [7:0] n15457;
wire      [7:0] n15458;
wire      [7:0] n15459;
wire      [7:0] n1546;
wire      [7:0] n15460;
wire      [7:0] n15461;
wire      [7:0] n15462;
wire      [7:0] n15463;
wire      [7:0] n15464;
wire      [7:0] n15465;
wire      [7:0] n15466;
wire      [7:0] n15467;
wire      [7:0] n15468;
wire      [7:0] n15469;
wire      [7:0] n1547;
wire      [7:0] n15470;
wire      [7:0] n15471;
wire      [7:0] n15472;
wire      [7:0] n15473;
wire      [7:0] n15474;
wire      [7:0] n15475;
wire      [7:0] n15476;
wire      [7:0] n15477;
wire      [7:0] n15478;
wire      [7:0] n15479;
wire      [7:0] n1548;
wire      [7:0] n15480;
wire      [7:0] n15481;
wire      [7:0] n15482;
wire      [7:0] n15483;
wire      [7:0] n15484;
wire      [7:0] n15485;
wire      [7:0] n15486;
wire      [7:0] n15487;
wire      [7:0] n15488;
wire      [7:0] n15489;
wire      [7:0] n1549;
wire      [7:0] n15490;
wire      [7:0] n15491;
wire      [7:0] n15492;
wire      [7:0] n15493;
wire      [7:0] n15494;
wire      [7:0] n15495;
wire      [7:0] n15496;
wire      [7:0] n15497;
wire      [7:0] n15498;
wire      [7:0] n15499;
wire      [7:0] n1550;
wire      [7:0] n15500;
wire      [7:0] n15501;
wire      [7:0] n15502;
wire      [7:0] n15503;
wire      [7:0] n15504;
wire      [7:0] n15505;
wire      [7:0] n15506;
wire      [7:0] n15507;
wire      [7:0] n15508;
wire      [7:0] n15509;
wire      [7:0] n1551;
wire      [7:0] n15510;
wire      [7:0] n15511;
wire      [7:0] n15512;
wire      [7:0] n15513;
wire      [7:0] n15514;
wire      [7:0] n15515;
wire      [7:0] n15516;
wire      [7:0] n15517;
wire      [7:0] n15518;
wire      [7:0] n15519;
wire      [7:0] n1552;
wire      [7:0] n15520;
wire      [7:0] n15521;
wire      [7:0] n15522;
wire      [7:0] n15523;
wire      [7:0] n15524;
wire      [7:0] n15525;
wire      [7:0] n15526;
wire      [7:0] n15527;
wire      [7:0] n15528;
wire      [7:0] n15529;
wire      [7:0] n1553;
wire      [7:0] n15530;
wire      [7:0] n15531;
wire      [7:0] n15532;
wire      [7:0] n15533;
wire      [7:0] n15534;
wire      [7:0] n15535;
wire      [7:0] n15536;
wire      [7:0] n15537;
wire      [7:0] n15538;
wire      [7:0] n15539;
wire      [7:0] n1554;
wire      [7:0] n15540;
wire      [7:0] n15541;
wire      [7:0] n15542;
wire      [7:0] n15543;
wire      [7:0] n15544;
wire      [7:0] n15545;
wire      [7:0] n15546;
wire      [7:0] n15547;
wire      [7:0] n15548;
wire      [7:0] n15549;
wire      [7:0] n1555;
wire      [7:0] n15550;
wire      [7:0] n15551;
wire      [7:0] n15552;
wire      [7:0] n15553;
wire      [7:0] n15554;
wire      [7:0] n15555;
wire      [7:0] n15556;
wire      [7:0] n15557;
wire      [7:0] n15558;
wire      [7:0] n15559;
wire      [7:0] n1556;
wire      [7:0] n15560;
wire      [7:0] n15561;
wire      [7:0] n15562;
wire      [7:0] n15563;
wire      [7:0] n15564;
wire      [7:0] n15565;
wire      [7:0] n15566;
wire      [7:0] n15567;
wire      [7:0] n15568;
wire      [7:0] n15569;
wire      [7:0] n1557;
wire      [7:0] n15570;
wire      [7:0] n15571;
wire      [7:0] n15572;
wire      [7:0] n15573;
wire      [7:0] n15574;
wire      [7:0] n15575;
wire      [7:0] n15576;
wire      [7:0] n15577;
wire      [7:0] n15578;
wire      [7:0] n15579;
wire      [7:0] n1558;
wire      [7:0] n15580;
wire      [7:0] n15581;
wire      [7:0] n15582;
wire      [7:0] n15583;
wire      [7:0] n15584;
wire      [7:0] n15585;
wire      [7:0] n15586;
wire      [7:0] n15587;
wire      [7:0] n15588;
wire      [7:0] n15589;
wire      [7:0] n1559;
wire      [7:0] n15590;
wire      [7:0] n15591;
wire      [7:0] n15592;
wire      [7:0] n15593;
wire      [7:0] n15594;
wire      [7:0] n15595;
wire      [7:0] n15596;
wire      [7:0] n15597;
wire      [7:0] n15598;
wire      [7:0] n15599;
wire      [7:0] n156;
wire      [7:0] n1560;
wire      [7:0] n15600;
wire      [7:0] n15601;
wire      [7:0] n15602;
wire      [7:0] n15603;
wire      [7:0] n15604;
wire      [7:0] n15605;
wire      [7:0] n15606;
wire      [7:0] n15607;
wire      [7:0] n15608;
wire      [7:0] n15609;
wire      [7:0] n1561;
wire      [7:0] n15610;
wire      [7:0] n15611;
wire      [7:0] n15612;
wire      [7:0] n15613;
wire      [7:0] n15614;
wire      [7:0] n15615;
wire      [7:0] n15616;
wire      [7:0] n15617;
wire      [7:0] n15618;
wire      [7:0] n15619;
wire      [7:0] n1562;
wire      [7:0] n15620;
wire      [7:0] n15621;
wire      [7:0] n15622;
wire      [7:0] n15623;
wire      [7:0] n15624;
wire      [7:0] n15625;
wire      [7:0] n15626;
wire      [7:0] n15627;
wire      [7:0] n15628;
wire      [7:0] n15629;
wire      [7:0] n1563;
wire      [7:0] n15630;
wire      [7:0] n15631;
wire      [7:0] n15632;
wire      [7:0] n15633;
wire      [7:0] n15634;
wire      [7:0] n15635;
wire      [7:0] n15636;
wire      [7:0] n15637;
wire      [7:0] n15638;
wire      [7:0] n15639;
wire      [7:0] n1564;
wire      [7:0] n15640;
wire      [7:0] n15641;
wire      [7:0] n15642;
wire      [7:0] n15643;
wire      [7:0] n15644;
wire      [7:0] n15645;
wire      [7:0] n15646;
wire      [7:0] n15647;
wire      [7:0] n15648;
wire      [7:0] n15649;
wire      [7:0] n1565;
wire      [7:0] n15650;
wire      [7:0] n15651;
wire      [7:0] n15652;
wire      [7:0] n15653;
wire      [7:0] n15654;
wire      [7:0] n15655;
wire      [7:0] n15656;
wire      [7:0] n15657;
wire      [7:0] n15658;
wire      [7:0] n15659;
wire      [7:0] n1566;
wire      [7:0] n15660;
wire      [7:0] n15661;
wire      [7:0] n15662;
wire      [7:0] n15663;
wire      [7:0] n15664;
wire      [7:0] n15665;
wire      [7:0] n15666;
wire      [7:0] n15667;
wire      [7:0] n15668;
wire      [7:0] n15669;
wire      [7:0] n1567;
wire      [7:0] n15670;
wire      [7:0] n15671;
wire      [7:0] n15672;
wire      [7:0] n15673;
wire      [7:0] n15674;
wire      [7:0] n15675;
wire      [7:0] n15676;
wire            n15677;
wire      [7:0] n15678;
wire            n15679;
wire      [7:0] n1568;
wire      [7:0] n15680;
wire            n15681;
wire      [7:0] n15682;
wire            n15683;
wire      [7:0] n15684;
wire            n15685;
wire      [7:0] n15686;
wire            n15687;
wire      [7:0] n15688;
wire            n15689;
wire      [7:0] n1569;
wire      [7:0] n15690;
wire            n15691;
wire      [7:0] n15692;
wire            n15693;
wire      [7:0] n15694;
wire            n15695;
wire      [7:0] n15696;
wire            n15697;
wire      [7:0] n15698;
wire            n15699;
wire      [7:0] n1570;
wire      [7:0] n15700;
wire            n15701;
wire      [7:0] n15702;
wire            n15703;
wire      [7:0] n15704;
wire            n15705;
wire      [7:0] n15706;
wire            n15707;
wire      [7:0] n15708;
wire            n15709;
wire      [7:0] n1571;
wire      [7:0] n15710;
wire            n15711;
wire      [7:0] n15712;
wire            n15713;
wire      [7:0] n15714;
wire            n15715;
wire      [7:0] n15716;
wire            n15717;
wire      [7:0] n15718;
wire            n15719;
wire      [7:0] n1572;
wire      [7:0] n15720;
wire            n15721;
wire      [7:0] n15722;
wire            n15723;
wire      [7:0] n15724;
wire            n15725;
wire      [7:0] n15726;
wire            n15727;
wire      [7:0] n15728;
wire            n15729;
wire      [7:0] n1573;
wire      [7:0] n15730;
wire            n15731;
wire      [7:0] n15732;
wire            n15733;
wire      [7:0] n15734;
wire            n15735;
wire      [7:0] n15736;
wire            n15737;
wire      [7:0] n15738;
wire            n15739;
wire      [7:0] n1574;
wire      [7:0] n15740;
wire            n15741;
wire      [7:0] n15742;
wire            n15743;
wire      [7:0] n15744;
wire            n15745;
wire      [7:0] n15746;
wire            n15747;
wire      [7:0] n15748;
wire            n15749;
wire      [7:0] n1575;
wire      [7:0] n15750;
wire            n15751;
wire      [7:0] n15752;
wire            n15753;
wire      [7:0] n15754;
wire            n15755;
wire      [7:0] n15756;
wire            n15757;
wire      [7:0] n15758;
wire            n15759;
wire      [7:0] n1576;
wire      [7:0] n15760;
wire            n15761;
wire      [7:0] n15762;
wire            n15763;
wire      [7:0] n15764;
wire            n15765;
wire      [7:0] n15766;
wire            n15767;
wire      [7:0] n15768;
wire            n15769;
wire      [7:0] n1577;
wire      [7:0] n15770;
wire            n15771;
wire      [7:0] n15772;
wire            n15773;
wire      [7:0] n15774;
wire            n15775;
wire      [7:0] n15776;
wire            n15777;
wire      [7:0] n15778;
wire            n15779;
wire      [7:0] n1578;
wire      [7:0] n15780;
wire            n15781;
wire      [7:0] n15782;
wire            n15783;
wire      [7:0] n15784;
wire            n15785;
wire      [7:0] n15786;
wire            n15787;
wire      [7:0] n15788;
wire            n15789;
wire      [7:0] n1579;
wire      [7:0] n15790;
wire            n15791;
wire      [7:0] n15792;
wire            n15793;
wire      [7:0] n15794;
wire            n15795;
wire      [7:0] n15796;
wire            n15797;
wire      [7:0] n15798;
wire            n15799;
wire            n158;
wire      [7:0] n1580;
wire      [7:0] n15800;
wire            n15801;
wire      [7:0] n15802;
wire            n15803;
wire      [7:0] n15804;
wire            n15805;
wire      [7:0] n15806;
wire            n15807;
wire      [7:0] n15808;
wire            n15809;
wire      [7:0] n1581;
wire      [7:0] n15810;
wire            n15811;
wire      [7:0] n15812;
wire            n15813;
wire      [7:0] n15814;
wire            n15815;
wire      [7:0] n15816;
wire            n15817;
wire      [7:0] n15818;
wire            n15819;
wire      [7:0] n1582;
wire      [7:0] n15820;
wire            n15821;
wire      [7:0] n15822;
wire            n15823;
wire      [7:0] n15824;
wire            n15825;
wire      [7:0] n15826;
wire            n15827;
wire      [7:0] n15828;
wire            n15829;
wire      [7:0] n1583;
wire      [7:0] n15830;
wire            n15831;
wire      [7:0] n15832;
wire            n15833;
wire      [7:0] n15834;
wire            n15835;
wire      [7:0] n15836;
wire            n15837;
wire      [7:0] n15838;
wire            n15839;
wire      [7:0] n1584;
wire      [7:0] n15840;
wire            n15841;
wire      [7:0] n15842;
wire            n15843;
wire      [7:0] n15844;
wire            n15845;
wire      [7:0] n15846;
wire            n15847;
wire      [7:0] n15848;
wire            n15849;
wire      [7:0] n1585;
wire      [7:0] n15850;
wire            n15851;
wire      [7:0] n15852;
wire            n15853;
wire      [7:0] n15854;
wire            n15855;
wire      [7:0] n15856;
wire            n15857;
wire      [7:0] n15858;
wire            n15859;
wire      [7:0] n1586;
wire      [7:0] n15860;
wire            n15861;
wire      [7:0] n15862;
wire            n15863;
wire      [7:0] n15864;
wire            n15865;
wire      [7:0] n15866;
wire            n15867;
wire      [7:0] n15868;
wire            n15869;
wire      [7:0] n1587;
wire      [7:0] n15870;
wire            n15871;
wire      [7:0] n15872;
wire            n15873;
wire      [7:0] n15874;
wire            n15875;
wire      [7:0] n15876;
wire            n15877;
wire      [7:0] n15878;
wire            n15879;
wire      [7:0] n1588;
wire      [7:0] n15880;
wire            n15881;
wire      [7:0] n15882;
wire            n15883;
wire      [7:0] n15884;
wire            n15885;
wire      [7:0] n15886;
wire            n15887;
wire      [7:0] n15888;
wire            n15889;
wire      [7:0] n1589;
wire      [7:0] n15890;
wire            n15891;
wire      [7:0] n15892;
wire            n15893;
wire      [7:0] n15894;
wire            n15895;
wire      [7:0] n15896;
wire            n15897;
wire      [7:0] n15898;
wire            n15899;
wire      [7:0] n1590;
wire      [7:0] n15900;
wire            n15901;
wire      [7:0] n15902;
wire            n15903;
wire      [7:0] n15904;
wire            n15905;
wire      [7:0] n15906;
wire            n15907;
wire      [7:0] n15908;
wire            n15909;
wire      [7:0] n1591;
wire      [7:0] n15910;
wire            n15911;
wire      [7:0] n15912;
wire            n15913;
wire      [7:0] n15914;
wire            n15915;
wire      [7:0] n15916;
wire            n15917;
wire      [7:0] n15918;
wire            n15919;
wire      [7:0] n1592;
wire      [7:0] n15920;
wire            n15921;
wire      [7:0] n15922;
wire            n15923;
wire      [7:0] n15924;
wire            n15925;
wire      [7:0] n15926;
wire            n15927;
wire      [7:0] n15928;
wire            n15929;
wire      [7:0] n1593;
wire      [7:0] n15930;
wire            n15931;
wire      [7:0] n15932;
wire            n15933;
wire      [7:0] n15934;
wire            n15935;
wire      [7:0] n15936;
wire            n15937;
wire      [7:0] n15938;
wire            n15939;
wire      [7:0] n1594;
wire      [7:0] n15940;
wire            n15941;
wire      [7:0] n15942;
wire            n15943;
wire      [7:0] n15944;
wire            n15945;
wire      [7:0] n15946;
wire            n15947;
wire      [7:0] n15948;
wire            n15949;
wire      [7:0] n1595;
wire      [7:0] n15950;
wire            n15951;
wire      [7:0] n15952;
wire            n15953;
wire      [7:0] n15954;
wire            n15955;
wire      [7:0] n15956;
wire            n15957;
wire      [7:0] n15958;
wire            n15959;
wire      [7:0] n1596;
wire      [7:0] n15960;
wire            n15961;
wire      [7:0] n15962;
wire            n15963;
wire      [7:0] n15964;
wire            n15965;
wire      [7:0] n15966;
wire            n15967;
wire      [7:0] n15968;
wire            n15969;
wire      [7:0] n1597;
wire      [7:0] n15970;
wire            n15971;
wire      [7:0] n15972;
wire            n15973;
wire      [7:0] n15974;
wire            n15975;
wire      [7:0] n15976;
wire            n15977;
wire      [7:0] n15978;
wire            n15979;
wire      [7:0] n1598;
wire      [7:0] n15980;
wire            n15981;
wire      [7:0] n15982;
wire            n15983;
wire      [7:0] n15984;
wire            n15985;
wire      [7:0] n15986;
wire            n15987;
wire      [7:0] n15988;
wire            n15989;
wire      [7:0] n1599;
wire      [7:0] n15990;
wire            n15991;
wire      [7:0] n15992;
wire            n15993;
wire      [7:0] n15994;
wire            n15995;
wire      [7:0] n15996;
wire            n15997;
wire      [7:0] n15998;
wire            n15999;
wire            n16;
wire      [7:0] n160;
wire      [7:0] n1600;
wire      [7:0] n16000;
wire            n16001;
wire      [7:0] n16002;
wire            n16003;
wire      [7:0] n16004;
wire            n16005;
wire      [7:0] n16006;
wire            n16007;
wire      [7:0] n16008;
wire            n16009;
wire      [7:0] n1601;
wire      [7:0] n16010;
wire            n16011;
wire      [7:0] n16012;
wire            n16013;
wire      [7:0] n16014;
wire            n16015;
wire      [7:0] n16016;
wire            n16017;
wire      [7:0] n16018;
wire            n16019;
wire      [7:0] n1602;
wire      [7:0] n16020;
wire            n16021;
wire      [7:0] n16022;
wire            n16023;
wire      [7:0] n16024;
wire            n16025;
wire      [7:0] n16026;
wire            n16027;
wire      [7:0] n16028;
wire            n16029;
wire      [7:0] n1603;
wire      [7:0] n16030;
wire            n16031;
wire      [7:0] n16032;
wire            n16033;
wire      [7:0] n16034;
wire            n16035;
wire      [7:0] n16036;
wire            n16037;
wire      [7:0] n16038;
wire            n16039;
wire      [7:0] n1604;
wire      [7:0] n16040;
wire            n16041;
wire      [7:0] n16042;
wire            n16043;
wire      [7:0] n16044;
wire            n16045;
wire      [7:0] n16046;
wire            n16047;
wire      [7:0] n16048;
wire            n16049;
wire      [7:0] n1605;
wire      [7:0] n16050;
wire            n16051;
wire      [7:0] n16052;
wire            n16053;
wire      [7:0] n16054;
wire            n16055;
wire      [7:0] n16056;
wire            n16057;
wire      [7:0] n16058;
wire            n16059;
wire      [7:0] n1606;
wire      [7:0] n16060;
wire            n16061;
wire      [7:0] n16062;
wire            n16063;
wire      [7:0] n16064;
wire            n16065;
wire      [7:0] n16066;
wire            n16067;
wire      [7:0] n16068;
wire            n16069;
wire      [7:0] n1607;
wire      [7:0] n16070;
wire            n16071;
wire      [7:0] n16072;
wire            n16073;
wire      [7:0] n16074;
wire            n16075;
wire      [7:0] n16076;
wire            n16077;
wire      [7:0] n16078;
wire            n16079;
wire      [7:0] n1608;
wire      [7:0] n16080;
wire            n16081;
wire      [7:0] n16082;
wire            n16083;
wire      [7:0] n16084;
wire            n16085;
wire      [7:0] n16086;
wire            n16087;
wire      [7:0] n16088;
wire            n16089;
wire      [7:0] n1609;
wire      [7:0] n16090;
wire            n16091;
wire      [7:0] n16092;
wire            n16093;
wire      [7:0] n16094;
wire            n16095;
wire      [7:0] n16096;
wire            n16097;
wire      [7:0] n16098;
wire            n16099;
wire            n161;
wire      [7:0] n1610;
wire      [7:0] n16100;
wire            n16101;
wire      [7:0] n16102;
wire            n16103;
wire      [7:0] n16104;
wire            n16105;
wire      [7:0] n16106;
wire            n16107;
wire      [7:0] n16108;
wire            n16109;
wire      [7:0] n1611;
wire      [7:0] n16110;
wire            n16111;
wire      [7:0] n16112;
wire            n16113;
wire      [7:0] n16114;
wire            n16115;
wire      [7:0] n16116;
wire            n16117;
wire      [7:0] n16118;
wire            n16119;
wire      [7:0] n1612;
wire      [7:0] n16120;
wire            n16121;
wire      [7:0] n16122;
wire            n16123;
wire      [7:0] n16124;
wire            n16125;
wire      [7:0] n16126;
wire            n16127;
wire      [7:0] n16128;
wire            n16129;
wire      [7:0] n1613;
wire      [7:0] n16130;
wire            n16131;
wire      [7:0] n16132;
wire            n16133;
wire      [7:0] n16134;
wire            n16135;
wire      [7:0] n16136;
wire            n16137;
wire      [7:0] n16138;
wire            n16139;
wire      [7:0] n1614;
wire      [7:0] n16140;
wire            n16141;
wire      [7:0] n16142;
wire            n16143;
wire      [7:0] n16144;
wire            n16145;
wire      [7:0] n16146;
wire            n16147;
wire      [7:0] n16148;
wire            n16149;
wire      [7:0] n1615;
wire      [7:0] n16150;
wire            n16151;
wire      [7:0] n16152;
wire            n16153;
wire      [7:0] n16154;
wire            n16155;
wire      [7:0] n16156;
wire            n16157;
wire      [7:0] n16158;
wire            n16159;
wire      [7:0] n1616;
wire      [7:0] n16160;
wire            n16161;
wire      [7:0] n16162;
wire            n16163;
wire      [7:0] n16164;
wire            n16165;
wire      [7:0] n16166;
wire            n16167;
wire      [7:0] n16168;
wire            n16169;
wire      [7:0] n1617;
wire      [7:0] n16170;
wire            n16171;
wire      [7:0] n16172;
wire            n16173;
wire      [7:0] n16174;
wire            n16175;
wire      [7:0] n16176;
wire            n16177;
wire      [7:0] n16178;
wire            n16179;
wire      [7:0] n1618;
wire      [7:0] n16180;
wire            n16181;
wire      [7:0] n16182;
wire            n16183;
wire      [7:0] n16184;
wire            n16185;
wire      [7:0] n16186;
wire            n16187;
wire      [7:0] n16188;
wire      [7:0] n16189;
wire      [7:0] n1619;
wire      [7:0] n16190;
wire      [7:0] n16191;
wire      [7:0] n16192;
wire      [7:0] n16193;
wire      [7:0] n16194;
wire      [7:0] n16195;
wire      [7:0] n16196;
wire      [7:0] n16197;
wire      [7:0] n16198;
wire      [7:0] n16199;
wire      [7:0] n1620;
wire      [7:0] n16200;
wire      [7:0] n16201;
wire      [7:0] n16202;
wire      [7:0] n16203;
wire      [7:0] n16204;
wire      [7:0] n16205;
wire      [7:0] n16206;
wire      [7:0] n16207;
wire      [7:0] n16208;
wire      [7:0] n16209;
wire      [7:0] n1621;
wire      [7:0] n16210;
wire      [7:0] n16211;
wire      [7:0] n16212;
wire      [7:0] n16213;
wire      [7:0] n16214;
wire      [7:0] n16215;
wire      [7:0] n16216;
wire      [7:0] n16217;
wire      [7:0] n16218;
wire      [7:0] n16219;
wire      [7:0] n1622;
wire      [7:0] n16220;
wire      [7:0] n16221;
wire      [7:0] n16222;
wire      [7:0] n16223;
wire      [7:0] n16224;
wire      [7:0] n16225;
wire      [7:0] n16226;
wire      [7:0] n16227;
wire      [7:0] n16228;
wire      [7:0] n16229;
wire      [7:0] n1623;
wire      [7:0] n16230;
wire      [7:0] n16231;
wire      [7:0] n16232;
wire      [7:0] n16233;
wire      [7:0] n16234;
wire      [7:0] n16235;
wire      [7:0] n16236;
wire      [7:0] n16237;
wire      [7:0] n16238;
wire      [7:0] n16239;
wire      [7:0] n1624;
wire      [7:0] n16240;
wire      [7:0] n16241;
wire      [7:0] n16242;
wire      [7:0] n16243;
wire      [7:0] n16244;
wire      [7:0] n16245;
wire      [7:0] n16246;
wire      [7:0] n16247;
wire      [7:0] n16248;
wire      [7:0] n16249;
wire      [7:0] n1625;
wire      [7:0] n16250;
wire      [7:0] n16251;
wire      [7:0] n16252;
wire      [7:0] n16253;
wire      [7:0] n16254;
wire      [7:0] n16255;
wire      [7:0] n16256;
wire      [7:0] n16257;
wire      [7:0] n16258;
wire      [7:0] n16259;
wire      [7:0] n1626;
wire      [7:0] n16260;
wire      [7:0] n16261;
wire      [7:0] n16262;
wire      [7:0] n16263;
wire      [7:0] n16264;
wire      [7:0] n16265;
wire      [7:0] n16266;
wire      [7:0] n16267;
wire      [7:0] n16268;
wire      [7:0] n16269;
wire      [7:0] n1627;
wire      [7:0] n16270;
wire      [7:0] n16271;
wire      [7:0] n16272;
wire      [7:0] n16273;
wire      [7:0] n16274;
wire      [7:0] n16275;
wire      [7:0] n16276;
wire      [7:0] n16277;
wire      [7:0] n16278;
wire      [7:0] n16279;
wire      [7:0] n1628;
wire      [7:0] n16280;
wire      [7:0] n16281;
wire      [7:0] n16282;
wire      [7:0] n16283;
wire      [7:0] n16284;
wire      [7:0] n16285;
wire      [7:0] n16286;
wire      [7:0] n16287;
wire      [7:0] n16288;
wire      [7:0] n16289;
wire      [7:0] n1629;
wire      [7:0] n16290;
wire      [7:0] n16291;
wire      [7:0] n16292;
wire      [7:0] n16293;
wire      [7:0] n16294;
wire      [7:0] n16295;
wire      [7:0] n16296;
wire      [7:0] n16297;
wire      [7:0] n16298;
wire      [7:0] n16299;
wire      [7:0] n163;
wire      [7:0] n1630;
wire      [7:0] n16300;
wire      [7:0] n16301;
wire      [7:0] n16302;
wire      [7:0] n16303;
wire      [7:0] n16304;
wire      [7:0] n16305;
wire      [7:0] n16306;
wire      [7:0] n16307;
wire      [7:0] n16308;
wire      [7:0] n16309;
wire      [7:0] n1631;
wire      [7:0] n16310;
wire      [7:0] n16311;
wire      [7:0] n16312;
wire      [7:0] n16313;
wire      [7:0] n16314;
wire      [7:0] n16315;
wire      [7:0] n16316;
wire      [7:0] n16317;
wire      [7:0] n16318;
wire      [7:0] n16319;
wire      [7:0] n1632;
wire      [7:0] n16320;
wire      [7:0] n16321;
wire      [7:0] n16322;
wire      [7:0] n16323;
wire      [7:0] n16324;
wire      [7:0] n16325;
wire      [7:0] n16326;
wire      [7:0] n16327;
wire      [7:0] n16328;
wire      [7:0] n16329;
wire      [7:0] n1633;
wire      [7:0] n16330;
wire      [7:0] n16331;
wire      [7:0] n16332;
wire      [7:0] n16333;
wire      [7:0] n16334;
wire      [7:0] n16335;
wire      [7:0] n16336;
wire      [7:0] n16337;
wire      [7:0] n16338;
wire      [7:0] n16339;
wire      [7:0] n1634;
wire      [7:0] n16340;
wire      [7:0] n16341;
wire      [7:0] n16342;
wire      [7:0] n16343;
wire      [7:0] n16344;
wire      [7:0] n16345;
wire      [7:0] n16346;
wire      [7:0] n16347;
wire      [7:0] n16348;
wire      [7:0] n16349;
wire      [7:0] n1635;
wire      [7:0] n16350;
wire      [7:0] n16351;
wire      [7:0] n16352;
wire      [7:0] n16353;
wire      [7:0] n16354;
wire      [7:0] n16355;
wire      [7:0] n16356;
wire      [7:0] n16357;
wire      [7:0] n16358;
wire      [7:0] n16359;
wire      [7:0] n1636;
wire      [7:0] n16360;
wire      [7:0] n16361;
wire      [7:0] n16362;
wire      [7:0] n16363;
wire      [7:0] n16364;
wire      [7:0] n16365;
wire      [7:0] n16366;
wire      [7:0] n16367;
wire      [7:0] n16368;
wire      [7:0] n16369;
wire      [7:0] n1637;
wire      [7:0] n16370;
wire      [7:0] n16371;
wire      [7:0] n16372;
wire      [7:0] n16373;
wire      [7:0] n16374;
wire      [7:0] n16375;
wire      [7:0] n16376;
wire      [7:0] n16377;
wire      [7:0] n16378;
wire      [7:0] n16379;
wire      [7:0] n1638;
wire      [7:0] n16380;
wire      [7:0] n16381;
wire      [7:0] n16382;
wire      [7:0] n16383;
wire      [7:0] n16384;
wire      [7:0] n16385;
wire      [7:0] n16386;
wire      [7:0] n16387;
wire      [7:0] n16388;
wire      [7:0] n16389;
wire      [7:0] n1639;
wire      [7:0] n16390;
wire      [7:0] n16391;
wire      [7:0] n16392;
wire      [7:0] n16393;
wire      [7:0] n16394;
wire      [7:0] n16395;
wire      [7:0] n16396;
wire      [7:0] n16397;
wire      [7:0] n16398;
wire      [7:0] n16399;
wire      [7:0] n1640;
wire      [7:0] n16400;
wire      [7:0] n16401;
wire      [7:0] n16402;
wire      [7:0] n16403;
wire      [7:0] n16404;
wire      [7:0] n16405;
wire      [7:0] n16406;
wire      [7:0] n16407;
wire      [7:0] n16408;
wire      [7:0] n16409;
wire      [7:0] n1641;
wire      [7:0] n16410;
wire      [7:0] n16411;
wire      [7:0] n16412;
wire      [7:0] n16413;
wire      [7:0] n16414;
wire      [7:0] n16415;
wire      [7:0] n16416;
wire      [7:0] n16417;
wire      [7:0] n16418;
wire      [7:0] n16419;
wire      [7:0] n1642;
wire      [7:0] n16420;
wire      [7:0] n16421;
wire      [7:0] n16422;
wire      [7:0] n16423;
wire      [7:0] n16424;
wire      [7:0] n16425;
wire      [7:0] n16426;
wire      [7:0] n16427;
wire      [7:0] n16428;
wire      [7:0] n16429;
wire      [7:0] n1643;
wire      [7:0] n16430;
wire      [7:0] n16431;
wire      [7:0] n16432;
wire      [7:0] n16433;
wire      [7:0] n16434;
wire      [7:0] n16435;
wire      [7:0] n16436;
wire      [7:0] n16437;
wire      [7:0] n16438;
wire      [7:0] n16439;
wire      [7:0] n1644;
wire      [7:0] n16440;
wire      [7:0] n16441;
wire      [7:0] n16442;
wire      [7:0] n16443;
wire      [7:0] n16444;
wire      [7:0] n16445;
wire      [7:0] n16446;
wire     [71:0] n16447;
wire      [7:0] n16448;
wire            n16449;
wire      [7:0] n1645;
wire      [7:0] n16450;
wire            n16451;
wire      [7:0] n16452;
wire            n16453;
wire      [7:0] n16454;
wire            n16455;
wire      [7:0] n16456;
wire            n16457;
wire      [7:0] n16458;
wire            n16459;
wire      [7:0] n1646;
wire      [7:0] n16460;
wire            n16461;
wire      [7:0] n16462;
wire            n16463;
wire      [7:0] n16464;
wire            n16465;
wire      [7:0] n16466;
wire            n16467;
wire      [7:0] n16468;
wire            n16469;
wire      [7:0] n1647;
wire      [7:0] n16470;
wire            n16471;
wire      [7:0] n16472;
wire            n16473;
wire      [7:0] n16474;
wire            n16475;
wire      [7:0] n16476;
wire            n16477;
wire      [7:0] n16478;
wire            n16479;
wire      [7:0] n1648;
wire      [7:0] n16480;
wire            n16481;
wire      [7:0] n16482;
wire            n16483;
wire      [7:0] n16484;
wire            n16485;
wire      [7:0] n16486;
wire            n16487;
wire      [7:0] n16488;
wire            n16489;
wire      [7:0] n1649;
wire      [7:0] n16490;
wire            n16491;
wire      [7:0] n16492;
wire            n16493;
wire      [7:0] n16494;
wire            n16495;
wire      [7:0] n16496;
wire            n16497;
wire      [7:0] n16498;
wire            n16499;
wire            n165;
wire      [7:0] n1650;
wire      [7:0] n16500;
wire            n16501;
wire      [7:0] n16502;
wire            n16503;
wire      [7:0] n16504;
wire            n16505;
wire      [7:0] n16506;
wire            n16507;
wire      [7:0] n16508;
wire            n16509;
wire      [7:0] n1651;
wire      [7:0] n16510;
wire            n16511;
wire      [7:0] n16512;
wire            n16513;
wire      [7:0] n16514;
wire            n16515;
wire      [7:0] n16516;
wire            n16517;
wire      [7:0] n16518;
wire            n16519;
wire      [7:0] n1652;
wire      [7:0] n16520;
wire            n16521;
wire      [7:0] n16522;
wire            n16523;
wire      [7:0] n16524;
wire            n16525;
wire      [7:0] n16526;
wire            n16527;
wire      [7:0] n16528;
wire            n16529;
wire      [7:0] n1653;
wire      [7:0] n16530;
wire            n16531;
wire      [7:0] n16532;
wire            n16533;
wire      [7:0] n16534;
wire            n16535;
wire      [7:0] n16536;
wire            n16537;
wire      [7:0] n16538;
wire            n16539;
wire      [7:0] n1654;
wire      [7:0] n16540;
wire            n16541;
wire      [7:0] n16542;
wire            n16543;
wire      [7:0] n16544;
wire            n16545;
wire      [7:0] n16546;
wire            n16547;
wire      [7:0] n16548;
wire            n16549;
wire      [7:0] n1655;
wire      [7:0] n16550;
wire            n16551;
wire      [7:0] n16552;
wire            n16553;
wire      [7:0] n16554;
wire            n16555;
wire      [7:0] n16556;
wire            n16557;
wire      [7:0] n16558;
wire            n16559;
wire      [7:0] n1656;
wire      [7:0] n16560;
wire            n16561;
wire      [7:0] n16562;
wire            n16563;
wire      [7:0] n16564;
wire            n16565;
wire      [7:0] n16566;
wire            n16567;
wire      [7:0] n16568;
wire            n16569;
wire      [7:0] n1657;
wire      [7:0] n16570;
wire            n16571;
wire      [7:0] n16572;
wire            n16573;
wire      [7:0] n16574;
wire            n16575;
wire      [7:0] n16576;
wire            n16577;
wire      [7:0] n16578;
wire            n16579;
wire      [7:0] n1658;
wire      [7:0] n16580;
wire            n16581;
wire      [7:0] n16582;
wire            n16583;
wire      [7:0] n16584;
wire            n16585;
wire      [7:0] n16586;
wire            n16587;
wire      [7:0] n16588;
wire            n16589;
wire      [7:0] n1659;
wire      [7:0] n16590;
wire            n16591;
wire      [7:0] n16592;
wire            n16593;
wire      [7:0] n16594;
wire            n16595;
wire      [7:0] n16596;
wire            n16597;
wire      [7:0] n16598;
wire            n16599;
wire      [7:0] n166;
wire      [7:0] n1660;
wire      [7:0] n16600;
wire            n16601;
wire      [7:0] n16602;
wire            n16603;
wire      [7:0] n16604;
wire            n16605;
wire      [7:0] n16606;
wire            n16607;
wire      [7:0] n16608;
wire            n16609;
wire      [7:0] n1661;
wire      [7:0] n16610;
wire            n16611;
wire      [7:0] n16612;
wire            n16613;
wire      [7:0] n16614;
wire            n16615;
wire      [7:0] n16616;
wire            n16617;
wire      [7:0] n16618;
wire            n16619;
wire      [7:0] n1662;
wire      [7:0] n16620;
wire            n16621;
wire      [7:0] n16622;
wire            n16623;
wire      [7:0] n16624;
wire            n16625;
wire      [7:0] n16626;
wire            n16627;
wire      [7:0] n16628;
wire            n16629;
wire      [7:0] n1663;
wire      [7:0] n16630;
wire            n16631;
wire      [7:0] n16632;
wire            n16633;
wire      [7:0] n16634;
wire            n16635;
wire      [7:0] n16636;
wire            n16637;
wire      [7:0] n16638;
wire            n16639;
wire      [7:0] n1664;
wire      [7:0] n16640;
wire            n16641;
wire      [7:0] n16642;
wire            n16643;
wire      [7:0] n16644;
wire            n16645;
wire      [7:0] n16646;
wire            n16647;
wire      [7:0] n16648;
wire            n16649;
wire      [7:0] n1665;
wire      [7:0] n16650;
wire            n16651;
wire      [7:0] n16652;
wire            n16653;
wire      [7:0] n16654;
wire            n16655;
wire      [7:0] n16656;
wire            n16657;
wire      [7:0] n16658;
wire            n16659;
wire      [7:0] n1666;
wire      [7:0] n16660;
wire            n16661;
wire      [7:0] n16662;
wire            n16663;
wire      [7:0] n16664;
wire            n16665;
wire      [7:0] n16666;
wire            n16667;
wire      [7:0] n16668;
wire            n16669;
wire      [7:0] n1667;
wire      [7:0] n16670;
wire            n16671;
wire      [7:0] n16672;
wire            n16673;
wire      [7:0] n16674;
wire            n16675;
wire      [7:0] n16676;
wire            n16677;
wire      [7:0] n16678;
wire            n16679;
wire      [7:0] n1668;
wire      [7:0] n16680;
wire            n16681;
wire      [7:0] n16682;
wire            n16683;
wire      [7:0] n16684;
wire            n16685;
wire      [7:0] n16686;
wire            n16687;
wire      [7:0] n16688;
wire            n16689;
wire      [7:0] n1669;
wire      [7:0] n16690;
wire            n16691;
wire      [7:0] n16692;
wire            n16693;
wire      [7:0] n16694;
wire            n16695;
wire      [7:0] n16696;
wire            n16697;
wire      [7:0] n16698;
wire            n16699;
wire      [7:0] n1670;
wire      [7:0] n16700;
wire            n16701;
wire      [7:0] n16702;
wire            n16703;
wire      [7:0] n16704;
wire            n16705;
wire      [7:0] n16706;
wire            n16707;
wire      [7:0] n16708;
wire            n16709;
wire      [7:0] n1671;
wire      [7:0] n16710;
wire            n16711;
wire      [7:0] n16712;
wire            n16713;
wire      [7:0] n16714;
wire            n16715;
wire      [7:0] n16716;
wire            n16717;
wire      [7:0] n16718;
wire            n16719;
wire      [7:0] n1672;
wire      [7:0] n16720;
wire            n16721;
wire      [7:0] n16722;
wire            n16723;
wire      [7:0] n16724;
wire            n16725;
wire      [7:0] n16726;
wire            n16727;
wire      [7:0] n16728;
wire            n16729;
wire      [7:0] n1673;
wire      [7:0] n16730;
wire            n16731;
wire      [7:0] n16732;
wire            n16733;
wire      [7:0] n16734;
wire            n16735;
wire      [7:0] n16736;
wire            n16737;
wire      [7:0] n16738;
wire            n16739;
wire      [7:0] n1674;
wire      [7:0] n16740;
wire            n16741;
wire      [7:0] n16742;
wire            n16743;
wire      [7:0] n16744;
wire            n16745;
wire      [7:0] n16746;
wire            n16747;
wire      [7:0] n16748;
wire            n16749;
wire      [7:0] n1675;
wire      [7:0] n16750;
wire            n16751;
wire      [7:0] n16752;
wire            n16753;
wire      [7:0] n16754;
wire            n16755;
wire      [7:0] n16756;
wire            n16757;
wire      [7:0] n16758;
wire            n16759;
wire      [7:0] n1676;
wire      [7:0] n16760;
wire            n16761;
wire      [7:0] n16762;
wire            n16763;
wire      [7:0] n16764;
wire            n16765;
wire      [7:0] n16766;
wire            n16767;
wire      [7:0] n16768;
wire            n16769;
wire      [7:0] n1677;
wire      [7:0] n16770;
wire            n16771;
wire      [7:0] n16772;
wire            n16773;
wire      [7:0] n16774;
wire            n16775;
wire      [7:0] n16776;
wire            n16777;
wire      [7:0] n16778;
wire            n16779;
wire      [7:0] n1678;
wire      [7:0] n16780;
wire            n16781;
wire      [7:0] n16782;
wire            n16783;
wire      [7:0] n16784;
wire            n16785;
wire      [7:0] n16786;
wire            n16787;
wire      [7:0] n16788;
wire            n16789;
wire      [7:0] n1679;
wire      [7:0] n16790;
wire            n16791;
wire      [7:0] n16792;
wire            n16793;
wire      [7:0] n16794;
wire            n16795;
wire      [7:0] n16796;
wire            n16797;
wire      [7:0] n16798;
wire            n16799;
wire            n168;
wire      [7:0] n1680;
wire      [7:0] n16800;
wire            n16801;
wire      [7:0] n16802;
wire            n16803;
wire      [7:0] n16804;
wire            n16805;
wire      [7:0] n16806;
wire            n16807;
wire      [7:0] n16808;
wire            n16809;
wire      [7:0] n1681;
wire      [7:0] n16810;
wire            n16811;
wire      [7:0] n16812;
wire            n16813;
wire      [7:0] n16814;
wire            n16815;
wire      [7:0] n16816;
wire            n16817;
wire      [7:0] n16818;
wire            n16819;
wire      [7:0] n1682;
wire      [7:0] n16820;
wire            n16821;
wire      [7:0] n16822;
wire            n16823;
wire      [7:0] n16824;
wire            n16825;
wire      [7:0] n16826;
wire            n16827;
wire      [7:0] n16828;
wire            n16829;
wire      [7:0] n1683;
wire      [7:0] n16830;
wire            n16831;
wire      [7:0] n16832;
wire            n16833;
wire      [7:0] n16834;
wire            n16835;
wire      [7:0] n16836;
wire            n16837;
wire      [7:0] n16838;
wire            n16839;
wire      [7:0] n1684;
wire      [7:0] n16840;
wire            n16841;
wire      [7:0] n16842;
wire            n16843;
wire      [7:0] n16844;
wire            n16845;
wire      [7:0] n16846;
wire            n16847;
wire      [7:0] n16848;
wire            n16849;
wire      [7:0] n1685;
wire      [7:0] n16850;
wire            n16851;
wire      [7:0] n16852;
wire            n16853;
wire      [7:0] n16854;
wire            n16855;
wire      [7:0] n16856;
wire            n16857;
wire      [7:0] n16858;
wire            n16859;
wire      [7:0] n1686;
wire      [7:0] n16860;
wire            n16861;
wire      [7:0] n16862;
wire            n16863;
wire      [7:0] n16864;
wire            n16865;
wire      [7:0] n16866;
wire            n16867;
wire      [7:0] n16868;
wire            n16869;
wire      [7:0] n1687;
wire      [7:0] n16870;
wire            n16871;
wire      [7:0] n16872;
wire            n16873;
wire      [7:0] n16874;
wire            n16875;
wire      [7:0] n16876;
wire            n16877;
wire      [7:0] n16878;
wire            n16879;
wire      [7:0] n1688;
wire      [7:0] n16880;
wire            n16881;
wire      [7:0] n16882;
wire            n16883;
wire      [7:0] n16884;
wire            n16885;
wire      [7:0] n16886;
wire            n16887;
wire      [7:0] n16888;
wire            n16889;
wire      [7:0] n1689;
wire      [7:0] n16890;
wire            n16891;
wire      [7:0] n16892;
wire            n16893;
wire      [7:0] n16894;
wire            n16895;
wire      [7:0] n16896;
wire            n16897;
wire      [7:0] n16898;
wire            n16899;
wire      [7:0] n1690;
wire      [7:0] n16900;
wire            n16901;
wire      [7:0] n16902;
wire            n16903;
wire      [7:0] n16904;
wire            n16905;
wire      [7:0] n16906;
wire            n16907;
wire      [7:0] n16908;
wire            n16909;
wire      [7:0] n1691;
wire      [7:0] n16910;
wire            n16911;
wire      [7:0] n16912;
wire            n16913;
wire      [7:0] n16914;
wire            n16915;
wire      [7:0] n16916;
wire            n16917;
wire      [7:0] n16918;
wire            n16919;
wire      [7:0] n1692;
wire      [7:0] n16920;
wire            n16921;
wire      [7:0] n16922;
wire            n16923;
wire      [7:0] n16924;
wire            n16925;
wire      [7:0] n16926;
wire            n16927;
wire      [7:0] n16928;
wire            n16929;
wire      [7:0] n1693;
wire      [7:0] n16930;
wire            n16931;
wire      [7:0] n16932;
wire            n16933;
wire      [7:0] n16934;
wire            n16935;
wire      [7:0] n16936;
wire            n16937;
wire      [7:0] n16938;
wire            n16939;
wire      [7:0] n1694;
wire      [7:0] n16940;
wire            n16941;
wire      [7:0] n16942;
wire            n16943;
wire      [7:0] n16944;
wire            n16945;
wire      [7:0] n16946;
wire            n16947;
wire      [7:0] n16948;
wire            n16949;
wire      [7:0] n1695;
wire      [7:0] n16950;
wire            n16951;
wire      [7:0] n16952;
wire            n16953;
wire      [7:0] n16954;
wire            n16955;
wire      [7:0] n16956;
wire            n16957;
wire      [7:0] n16958;
wire            n16959;
wire      [7:0] n1696;
wire      [7:0] n16960;
wire      [7:0] n16961;
wire      [7:0] n16962;
wire      [7:0] n16963;
wire      [7:0] n16964;
wire      [7:0] n16965;
wire      [7:0] n16966;
wire      [7:0] n16967;
wire      [7:0] n16968;
wire      [7:0] n16969;
wire      [7:0] n1697;
wire      [7:0] n16970;
wire      [7:0] n16971;
wire      [7:0] n16972;
wire      [7:0] n16973;
wire      [7:0] n16974;
wire      [7:0] n16975;
wire      [7:0] n16976;
wire      [7:0] n16977;
wire      [7:0] n16978;
wire      [7:0] n16979;
wire      [7:0] n1698;
wire      [7:0] n16980;
wire      [7:0] n16981;
wire      [7:0] n16982;
wire      [7:0] n16983;
wire      [7:0] n16984;
wire      [7:0] n16985;
wire      [7:0] n16986;
wire      [7:0] n16987;
wire      [7:0] n16988;
wire      [7:0] n16989;
wire      [7:0] n1699;
wire      [7:0] n16990;
wire      [7:0] n16991;
wire      [7:0] n16992;
wire      [7:0] n16993;
wire      [7:0] n16994;
wire      [7:0] n16995;
wire      [7:0] n16996;
wire      [7:0] n16997;
wire      [7:0] n16998;
wire      [7:0] n16999;
wire      [7:0] n170;
wire      [7:0] n1700;
wire      [7:0] n17000;
wire      [7:0] n17001;
wire      [7:0] n17002;
wire      [7:0] n17003;
wire      [7:0] n17004;
wire      [7:0] n17005;
wire      [7:0] n17006;
wire      [7:0] n17007;
wire      [7:0] n17008;
wire      [7:0] n17009;
wire      [7:0] n1701;
wire      [7:0] n17010;
wire      [7:0] n17011;
wire      [7:0] n17012;
wire      [7:0] n17013;
wire      [7:0] n17014;
wire      [7:0] n17015;
wire      [7:0] n17016;
wire      [7:0] n17017;
wire      [7:0] n17018;
wire      [7:0] n17019;
wire      [7:0] n1702;
wire      [7:0] n17020;
wire      [7:0] n17021;
wire      [7:0] n17022;
wire      [7:0] n17023;
wire      [7:0] n17024;
wire      [7:0] n17025;
wire      [7:0] n17026;
wire      [7:0] n17027;
wire      [7:0] n17028;
wire      [7:0] n17029;
wire      [7:0] n1703;
wire      [7:0] n17030;
wire      [7:0] n17031;
wire      [7:0] n17032;
wire      [7:0] n17033;
wire      [7:0] n17034;
wire      [7:0] n17035;
wire      [7:0] n17036;
wire      [7:0] n17037;
wire      [7:0] n17038;
wire      [7:0] n17039;
wire      [7:0] n1704;
wire      [7:0] n17040;
wire      [7:0] n17041;
wire      [7:0] n17042;
wire      [7:0] n17043;
wire      [7:0] n17044;
wire      [7:0] n17045;
wire      [7:0] n17046;
wire      [7:0] n17047;
wire      [7:0] n17048;
wire      [7:0] n17049;
wire      [7:0] n1705;
wire      [7:0] n17050;
wire      [7:0] n17051;
wire      [7:0] n17052;
wire      [7:0] n17053;
wire      [7:0] n17054;
wire      [7:0] n17055;
wire      [7:0] n17056;
wire      [7:0] n17057;
wire      [7:0] n17058;
wire      [7:0] n17059;
wire      [7:0] n1706;
wire      [7:0] n17060;
wire      [7:0] n17061;
wire      [7:0] n17062;
wire      [7:0] n17063;
wire      [7:0] n17064;
wire      [7:0] n17065;
wire      [7:0] n17066;
wire      [7:0] n17067;
wire      [7:0] n17068;
wire      [7:0] n17069;
wire      [7:0] n1707;
wire      [7:0] n17070;
wire      [7:0] n17071;
wire      [7:0] n17072;
wire      [7:0] n17073;
wire      [7:0] n17074;
wire      [7:0] n17075;
wire      [7:0] n17076;
wire      [7:0] n17077;
wire      [7:0] n17078;
wire      [7:0] n17079;
wire      [7:0] n1708;
wire      [7:0] n17080;
wire      [7:0] n17081;
wire      [7:0] n17082;
wire      [7:0] n17083;
wire      [7:0] n17084;
wire      [7:0] n17085;
wire      [7:0] n17086;
wire      [7:0] n17087;
wire      [7:0] n17088;
wire      [7:0] n17089;
wire      [7:0] n1709;
wire      [7:0] n17090;
wire      [7:0] n17091;
wire      [7:0] n17092;
wire      [7:0] n17093;
wire      [7:0] n17094;
wire      [7:0] n17095;
wire      [7:0] n17096;
wire      [7:0] n17097;
wire      [7:0] n17098;
wire      [7:0] n17099;
wire      [7:0] n1710;
wire      [7:0] n17100;
wire      [7:0] n17101;
wire      [7:0] n17102;
wire      [7:0] n17103;
wire      [7:0] n17104;
wire      [7:0] n17105;
wire      [7:0] n17106;
wire      [7:0] n17107;
wire      [7:0] n17108;
wire      [7:0] n17109;
wire      [7:0] n1711;
wire      [7:0] n17110;
wire      [7:0] n17111;
wire      [7:0] n17112;
wire      [7:0] n17113;
wire      [7:0] n17114;
wire      [7:0] n17115;
wire      [7:0] n17116;
wire      [7:0] n17117;
wire      [7:0] n17118;
wire      [7:0] n17119;
wire      [7:0] n1712;
wire      [7:0] n17120;
wire      [7:0] n17121;
wire      [7:0] n17122;
wire      [7:0] n17123;
wire      [7:0] n17124;
wire      [7:0] n17125;
wire      [7:0] n17126;
wire      [7:0] n17127;
wire      [7:0] n17128;
wire      [7:0] n17129;
wire      [7:0] n1713;
wire      [7:0] n17130;
wire      [7:0] n17131;
wire      [7:0] n17132;
wire      [7:0] n17133;
wire      [7:0] n17134;
wire      [7:0] n17135;
wire      [7:0] n17136;
wire      [7:0] n17137;
wire      [7:0] n17138;
wire      [7:0] n17139;
wire      [7:0] n1714;
wire      [7:0] n17140;
wire      [7:0] n17141;
wire      [7:0] n17142;
wire      [7:0] n17143;
wire      [7:0] n17144;
wire      [7:0] n17145;
wire      [7:0] n17146;
wire      [7:0] n17147;
wire      [7:0] n17148;
wire      [7:0] n17149;
wire      [7:0] n1715;
wire      [7:0] n17150;
wire      [7:0] n17151;
wire      [7:0] n17152;
wire      [7:0] n17153;
wire      [7:0] n17154;
wire      [7:0] n17155;
wire      [7:0] n17156;
wire      [7:0] n17157;
wire      [7:0] n17158;
wire      [7:0] n17159;
wire      [7:0] n1716;
wire      [7:0] n17160;
wire      [7:0] n17161;
wire      [7:0] n17162;
wire      [7:0] n17163;
wire      [7:0] n17164;
wire      [7:0] n17165;
wire      [7:0] n17166;
wire      [7:0] n17167;
wire      [7:0] n17168;
wire      [7:0] n17169;
wire      [7:0] n1717;
wire      [7:0] n17170;
wire      [7:0] n17171;
wire      [7:0] n17172;
wire      [7:0] n17173;
wire      [7:0] n17174;
wire      [7:0] n17175;
wire      [7:0] n17176;
wire      [7:0] n17177;
wire      [7:0] n17178;
wire      [7:0] n17179;
wire      [7:0] n1718;
wire      [7:0] n17180;
wire      [7:0] n17181;
wire      [7:0] n17182;
wire      [7:0] n17183;
wire      [7:0] n17184;
wire      [7:0] n17185;
wire      [7:0] n17186;
wire      [7:0] n17187;
wire      [7:0] n17188;
wire      [7:0] n17189;
wire      [7:0] n1719;
wire      [7:0] n17190;
wire      [7:0] n17191;
wire      [7:0] n17192;
wire      [7:0] n17193;
wire      [7:0] n17194;
wire      [7:0] n17195;
wire      [7:0] n17196;
wire      [7:0] n17197;
wire      [7:0] n17198;
wire      [7:0] n17199;
wire            n172;
wire      [7:0] n1720;
wire      [7:0] n17200;
wire      [7:0] n17201;
wire      [7:0] n17202;
wire      [7:0] n17203;
wire      [7:0] n17204;
wire      [7:0] n17205;
wire      [7:0] n17206;
wire      [7:0] n17207;
wire      [7:0] n17208;
wire      [7:0] n17209;
wire      [7:0] n1721;
wire      [7:0] n17210;
wire      [7:0] n17211;
wire      [7:0] n17212;
wire      [7:0] n17213;
wire      [7:0] n17214;
wire      [7:0] n17215;
wire      [7:0] n17216;
wire      [7:0] n17217;
wire      [7:0] n17218;
wire            n17219;
wire      [7:0] n1722;
wire      [7:0] n17220;
wire            n17221;
wire      [7:0] n17222;
wire            n17223;
wire      [7:0] n17224;
wire            n17225;
wire      [7:0] n17226;
wire            n17227;
wire      [7:0] n17228;
wire            n17229;
wire      [7:0] n1723;
wire      [7:0] n17230;
wire            n17231;
wire      [7:0] n17232;
wire            n17233;
wire      [7:0] n17234;
wire            n17235;
wire      [7:0] n17236;
wire            n17237;
wire      [7:0] n17238;
wire            n17239;
wire      [7:0] n1724;
wire      [7:0] n17240;
wire            n17241;
wire      [7:0] n17242;
wire            n17243;
wire      [7:0] n17244;
wire            n17245;
wire      [7:0] n17246;
wire            n17247;
wire      [7:0] n17248;
wire            n17249;
wire      [7:0] n1725;
wire      [7:0] n17250;
wire            n17251;
wire      [7:0] n17252;
wire            n17253;
wire      [7:0] n17254;
wire            n17255;
wire      [7:0] n17256;
wire            n17257;
wire      [7:0] n17258;
wire            n17259;
wire      [7:0] n1726;
wire      [7:0] n17260;
wire            n17261;
wire      [7:0] n17262;
wire            n17263;
wire      [7:0] n17264;
wire            n17265;
wire      [7:0] n17266;
wire            n17267;
wire      [7:0] n17268;
wire            n17269;
wire      [7:0] n1727;
wire      [7:0] n17270;
wire            n17271;
wire      [7:0] n17272;
wire            n17273;
wire      [7:0] n17274;
wire            n17275;
wire      [7:0] n17276;
wire            n17277;
wire      [7:0] n17278;
wire            n17279;
wire      [7:0] n1728;
wire      [7:0] n17280;
wire            n17281;
wire      [7:0] n17282;
wire            n17283;
wire      [7:0] n17284;
wire            n17285;
wire      [7:0] n17286;
wire            n17287;
wire      [7:0] n17288;
wire            n17289;
wire      [7:0] n1729;
wire      [7:0] n17290;
wire            n17291;
wire      [7:0] n17292;
wire            n17293;
wire      [7:0] n17294;
wire            n17295;
wire      [7:0] n17296;
wire            n17297;
wire      [7:0] n17298;
wire            n17299;
wire      [7:0] n1730;
wire      [7:0] n17300;
wire            n17301;
wire      [7:0] n17302;
wire            n17303;
wire      [7:0] n17304;
wire            n17305;
wire      [7:0] n17306;
wire            n17307;
wire      [7:0] n17308;
wire            n17309;
wire      [7:0] n1731;
wire      [7:0] n17310;
wire            n17311;
wire      [7:0] n17312;
wire            n17313;
wire      [7:0] n17314;
wire            n17315;
wire      [7:0] n17316;
wire            n17317;
wire      [7:0] n17318;
wire            n17319;
wire      [7:0] n1732;
wire      [7:0] n17320;
wire            n17321;
wire      [7:0] n17322;
wire            n17323;
wire      [7:0] n17324;
wire            n17325;
wire      [7:0] n17326;
wire            n17327;
wire      [7:0] n17328;
wire            n17329;
wire      [7:0] n1733;
wire      [7:0] n17330;
wire            n17331;
wire      [7:0] n17332;
wire            n17333;
wire      [7:0] n17334;
wire            n17335;
wire      [7:0] n17336;
wire            n17337;
wire      [7:0] n17338;
wire            n17339;
wire      [7:0] n1734;
wire      [7:0] n17340;
wire            n17341;
wire      [7:0] n17342;
wire            n17343;
wire      [7:0] n17344;
wire            n17345;
wire      [7:0] n17346;
wire            n17347;
wire      [7:0] n17348;
wire            n17349;
wire      [7:0] n1735;
wire      [7:0] n17350;
wire            n17351;
wire      [7:0] n17352;
wire            n17353;
wire      [7:0] n17354;
wire            n17355;
wire      [7:0] n17356;
wire            n17357;
wire      [7:0] n17358;
wire            n17359;
wire      [7:0] n1736;
wire      [7:0] n17360;
wire            n17361;
wire      [7:0] n17362;
wire            n17363;
wire      [7:0] n17364;
wire            n17365;
wire      [7:0] n17366;
wire            n17367;
wire      [7:0] n17368;
wire            n17369;
wire      [7:0] n1737;
wire      [7:0] n17370;
wire            n17371;
wire      [7:0] n17372;
wire            n17373;
wire      [7:0] n17374;
wire            n17375;
wire      [7:0] n17376;
wire            n17377;
wire      [7:0] n17378;
wire            n17379;
wire      [7:0] n1738;
wire      [7:0] n17380;
wire            n17381;
wire      [7:0] n17382;
wire            n17383;
wire      [7:0] n17384;
wire            n17385;
wire      [7:0] n17386;
wire            n17387;
wire      [7:0] n17388;
wire            n17389;
wire      [7:0] n1739;
wire      [7:0] n17390;
wire            n17391;
wire      [7:0] n17392;
wire            n17393;
wire      [7:0] n17394;
wire            n17395;
wire      [7:0] n17396;
wire            n17397;
wire      [7:0] n17398;
wire            n17399;
wire      [7:0] n174;
wire      [7:0] n1740;
wire      [7:0] n17400;
wire            n17401;
wire      [7:0] n17402;
wire            n17403;
wire      [7:0] n17404;
wire            n17405;
wire      [7:0] n17406;
wire            n17407;
wire      [7:0] n17408;
wire            n17409;
wire      [7:0] n1741;
wire      [7:0] n17410;
wire            n17411;
wire      [7:0] n17412;
wire            n17413;
wire      [7:0] n17414;
wire            n17415;
wire      [7:0] n17416;
wire            n17417;
wire      [7:0] n17418;
wire            n17419;
wire      [7:0] n1742;
wire      [7:0] n17420;
wire            n17421;
wire      [7:0] n17422;
wire            n17423;
wire      [7:0] n17424;
wire            n17425;
wire      [7:0] n17426;
wire            n17427;
wire      [7:0] n17428;
wire            n17429;
wire      [7:0] n1743;
wire      [7:0] n17430;
wire            n17431;
wire      [7:0] n17432;
wire            n17433;
wire      [7:0] n17434;
wire            n17435;
wire      [7:0] n17436;
wire            n17437;
wire      [7:0] n17438;
wire            n17439;
wire      [7:0] n1744;
wire      [7:0] n17440;
wire            n17441;
wire      [7:0] n17442;
wire            n17443;
wire      [7:0] n17444;
wire            n17445;
wire      [7:0] n17446;
wire            n17447;
wire      [7:0] n17448;
wire            n17449;
wire      [7:0] n1745;
wire      [7:0] n17450;
wire            n17451;
wire      [7:0] n17452;
wire            n17453;
wire      [7:0] n17454;
wire            n17455;
wire      [7:0] n17456;
wire            n17457;
wire      [7:0] n17458;
wire            n17459;
wire      [7:0] n1746;
wire      [7:0] n17460;
wire            n17461;
wire      [7:0] n17462;
wire            n17463;
wire      [7:0] n17464;
wire            n17465;
wire      [7:0] n17466;
wire            n17467;
wire      [7:0] n17468;
wire            n17469;
wire      [7:0] n1747;
wire      [7:0] n17470;
wire            n17471;
wire      [7:0] n17472;
wire            n17473;
wire      [7:0] n17474;
wire            n17475;
wire      [7:0] n17476;
wire            n17477;
wire      [7:0] n17478;
wire            n17479;
wire      [7:0] n1748;
wire      [7:0] n17480;
wire            n17481;
wire      [7:0] n17482;
wire            n17483;
wire      [7:0] n17484;
wire            n17485;
wire      [7:0] n17486;
wire            n17487;
wire      [7:0] n17488;
wire            n17489;
wire      [7:0] n1749;
wire      [7:0] n17490;
wire            n17491;
wire      [7:0] n17492;
wire            n17493;
wire      [7:0] n17494;
wire            n17495;
wire      [7:0] n17496;
wire            n17497;
wire      [7:0] n17498;
wire            n17499;
wire      [7:0] n1750;
wire      [7:0] n17500;
wire            n17501;
wire      [7:0] n17502;
wire            n17503;
wire      [7:0] n17504;
wire            n17505;
wire      [7:0] n17506;
wire            n17507;
wire      [7:0] n17508;
wire            n17509;
wire      [7:0] n1751;
wire      [7:0] n17510;
wire            n17511;
wire      [7:0] n17512;
wire            n17513;
wire      [7:0] n17514;
wire            n17515;
wire      [7:0] n17516;
wire            n17517;
wire      [7:0] n17518;
wire            n17519;
wire      [7:0] n1752;
wire      [7:0] n17520;
wire            n17521;
wire      [7:0] n17522;
wire            n17523;
wire      [7:0] n17524;
wire            n17525;
wire      [7:0] n17526;
wire            n17527;
wire      [7:0] n17528;
wire            n17529;
wire      [7:0] n1753;
wire      [7:0] n17530;
wire            n17531;
wire      [7:0] n17532;
wire            n17533;
wire      [7:0] n17534;
wire            n17535;
wire      [7:0] n17536;
wire            n17537;
wire      [7:0] n17538;
wire            n17539;
wire      [7:0] n1754;
wire      [7:0] n17540;
wire            n17541;
wire      [7:0] n17542;
wire            n17543;
wire      [7:0] n17544;
wire            n17545;
wire      [7:0] n17546;
wire            n17547;
wire      [7:0] n17548;
wire            n17549;
wire      [7:0] n1755;
wire      [7:0] n17550;
wire            n17551;
wire      [7:0] n17552;
wire            n17553;
wire      [7:0] n17554;
wire            n17555;
wire      [7:0] n17556;
wire            n17557;
wire      [7:0] n17558;
wire            n17559;
wire      [7:0] n1756;
wire      [7:0] n17560;
wire            n17561;
wire      [7:0] n17562;
wire            n17563;
wire      [7:0] n17564;
wire            n17565;
wire      [7:0] n17566;
wire            n17567;
wire      [7:0] n17568;
wire            n17569;
wire      [7:0] n1757;
wire      [7:0] n17570;
wire            n17571;
wire      [7:0] n17572;
wire            n17573;
wire      [7:0] n17574;
wire            n17575;
wire      [7:0] n17576;
wire            n17577;
wire      [7:0] n17578;
wire            n17579;
wire      [7:0] n1758;
wire      [7:0] n17580;
wire            n17581;
wire      [7:0] n17582;
wire            n17583;
wire      [7:0] n17584;
wire            n17585;
wire      [7:0] n17586;
wire            n17587;
wire      [7:0] n17588;
wire            n17589;
wire      [7:0] n1759;
wire      [7:0] n17590;
wire            n17591;
wire      [7:0] n17592;
wire            n17593;
wire      [7:0] n17594;
wire            n17595;
wire      [7:0] n17596;
wire            n17597;
wire      [7:0] n17598;
wire            n17599;
wire            n176;
wire      [7:0] n1760;
wire      [7:0] n17600;
wire            n17601;
wire      [7:0] n17602;
wire            n17603;
wire      [7:0] n17604;
wire            n17605;
wire      [7:0] n17606;
wire            n17607;
wire      [7:0] n17608;
wire            n17609;
wire      [7:0] n1761;
wire      [7:0] n17610;
wire            n17611;
wire      [7:0] n17612;
wire            n17613;
wire      [7:0] n17614;
wire            n17615;
wire      [7:0] n17616;
wire            n17617;
wire      [7:0] n17618;
wire            n17619;
wire      [7:0] n1762;
wire      [7:0] n17620;
wire            n17621;
wire      [7:0] n17622;
wire            n17623;
wire      [7:0] n17624;
wire            n17625;
wire      [7:0] n17626;
wire            n17627;
wire      [7:0] n17628;
wire            n17629;
wire      [7:0] n1763;
wire      [7:0] n17630;
wire            n17631;
wire      [7:0] n17632;
wire            n17633;
wire      [7:0] n17634;
wire            n17635;
wire      [7:0] n17636;
wire            n17637;
wire      [7:0] n17638;
wire            n17639;
wire      [7:0] n1764;
wire      [7:0] n17640;
wire            n17641;
wire      [7:0] n17642;
wire            n17643;
wire      [7:0] n17644;
wire            n17645;
wire      [7:0] n17646;
wire            n17647;
wire      [7:0] n17648;
wire            n17649;
wire      [7:0] n1765;
wire      [7:0] n17650;
wire            n17651;
wire      [7:0] n17652;
wire            n17653;
wire      [7:0] n17654;
wire            n17655;
wire      [7:0] n17656;
wire            n17657;
wire      [7:0] n17658;
wire            n17659;
wire      [7:0] n1766;
wire      [7:0] n17660;
wire            n17661;
wire      [7:0] n17662;
wire            n17663;
wire      [7:0] n17664;
wire            n17665;
wire      [7:0] n17666;
wire            n17667;
wire      [7:0] n17668;
wire            n17669;
wire      [7:0] n1767;
wire      [7:0] n17670;
wire            n17671;
wire      [7:0] n17672;
wire            n17673;
wire      [7:0] n17674;
wire            n17675;
wire      [7:0] n17676;
wire            n17677;
wire      [7:0] n17678;
wire            n17679;
wire      [7:0] n1768;
wire      [7:0] n17680;
wire            n17681;
wire      [7:0] n17682;
wire            n17683;
wire      [7:0] n17684;
wire            n17685;
wire      [7:0] n17686;
wire            n17687;
wire      [7:0] n17688;
wire            n17689;
wire      [7:0] n1769;
wire      [7:0] n17690;
wire            n17691;
wire      [7:0] n17692;
wire            n17693;
wire      [7:0] n17694;
wire            n17695;
wire      [7:0] n17696;
wire            n17697;
wire      [7:0] n17698;
wire            n17699;
wire      [7:0] n1770;
wire      [7:0] n17700;
wire            n17701;
wire      [7:0] n17702;
wire            n17703;
wire      [7:0] n17704;
wire            n17705;
wire      [7:0] n17706;
wire            n17707;
wire      [7:0] n17708;
wire            n17709;
wire      [7:0] n1771;
wire      [7:0] n17710;
wire            n17711;
wire      [7:0] n17712;
wire            n17713;
wire      [7:0] n17714;
wire            n17715;
wire      [7:0] n17716;
wire            n17717;
wire      [7:0] n17718;
wire            n17719;
wire      [7:0] n1772;
wire      [7:0] n17720;
wire            n17721;
wire      [7:0] n17722;
wire            n17723;
wire      [7:0] n17724;
wire            n17725;
wire      [7:0] n17726;
wire            n17727;
wire      [7:0] n17728;
wire            n17729;
wire      [7:0] n1773;
wire      [7:0] n17730;
wire      [7:0] n17731;
wire      [7:0] n17732;
wire      [7:0] n17733;
wire      [7:0] n17734;
wire      [7:0] n17735;
wire      [7:0] n17736;
wire      [7:0] n17737;
wire      [7:0] n17738;
wire      [7:0] n17739;
wire      [7:0] n1774;
wire      [7:0] n17740;
wire      [7:0] n17741;
wire      [7:0] n17742;
wire      [7:0] n17743;
wire      [7:0] n17744;
wire      [7:0] n17745;
wire      [7:0] n17746;
wire      [7:0] n17747;
wire      [7:0] n17748;
wire      [7:0] n17749;
wire      [7:0] n1775;
wire      [7:0] n17750;
wire      [7:0] n17751;
wire      [7:0] n17752;
wire      [7:0] n17753;
wire      [7:0] n17754;
wire      [7:0] n17755;
wire      [7:0] n17756;
wire      [7:0] n17757;
wire      [7:0] n17758;
wire      [7:0] n17759;
wire      [7:0] n1776;
wire      [7:0] n17760;
wire      [7:0] n17761;
wire      [7:0] n17762;
wire      [7:0] n17763;
wire      [7:0] n17764;
wire      [7:0] n17765;
wire      [7:0] n17766;
wire      [7:0] n17767;
wire      [7:0] n17768;
wire      [7:0] n17769;
wire      [7:0] n1777;
wire      [7:0] n17770;
wire      [7:0] n17771;
wire      [7:0] n17772;
wire      [7:0] n17773;
wire      [7:0] n17774;
wire      [7:0] n17775;
wire      [7:0] n17776;
wire      [7:0] n17777;
wire      [7:0] n17778;
wire      [7:0] n17779;
wire      [7:0] n1778;
wire      [7:0] n17780;
wire      [7:0] n17781;
wire      [7:0] n17782;
wire      [7:0] n17783;
wire      [7:0] n17784;
wire      [7:0] n17785;
wire      [7:0] n17786;
wire      [7:0] n17787;
wire      [7:0] n17788;
wire      [7:0] n17789;
wire      [7:0] n1779;
wire      [7:0] n17790;
wire      [7:0] n17791;
wire      [7:0] n17792;
wire      [7:0] n17793;
wire      [7:0] n17794;
wire      [7:0] n17795;
wire      [7:0] n17796;
wire      [7:0] n17797;
wire      [7:0] n17798;
wire      [7:0] n17799;
wire      [7:0] n178;
wire      [7:0] n1780;
wire      [7:0] n17800;
wire      [7:0] n17801;
wire      [7:0] n17802;
wire      [7:0] n17803;
wire      [7:0] n17804;
wire      [7:0] n17805;
wire      [7:0] n17806;
wire      [7:0] n17807;
wire      [7:0] n17808;
wire      [7:0] n17809;
wire      [7:0] n1781;
wire      [7:0] n17810;
wire      [7:0] n17811;
wire      [7:0] n17812;
wire      [7:0] n17813;
wire      [7:0] n17814;
wire      [7:0] n17815;
wire      [7:0] n17816;
wire      [7:0] n17817;
wire      [7:0] n17818;
wire      [7:0] n17819;
wire      [7:0] n1782;
wire      [7:0] n17820;
wire      [7:0] n17821;
wire      [7:0] n17822;
wire      [7:0] n17823;
wire      [7:0] n17824;
wire      [7:0] n17825;
wire      [7:0] n17826;
wire      [7:0] n17827;
wire      [7:0] n17828;
wire      [7:0] n17829;
wire      [7:0] n1783;
wire      [7:0] n17830;
wire      [7:0] n17831;
wire      [7:0] n17832;
wire      [7:0] n17833;
wire      [7:0] n17834;
wire      [7:0] n17835;
wire      [7:0] n17836;
wire      [7:0] n17837;
wire      [7:0] n17838;
wire      [7:0] n17839;
wire      [7:0] n1784;
wire      [7:0] n17840;
wire      [7:0] n17841;
wire      [7:0] n17842;
wire      [7:0] n17843;
wire      [7:0] n17844;
wire      [7:0] n17845;
wire      [7:0] n17846;
wire      [7:0] n17847;
wire      [7:0] n17848;
wire      [7:0] n17849;
wire      [7:0] n1785;
wire      [7:0] n17850;
wire      [7:0] n17851;
wire      [7:0] n17852;
wire      [7:0] n17853;
wire      [7:0] n17854;
wire      [7:0] n17855;
wire      [7:0] n17856;
wire      [7:0] n17857;
wire      [7:0] n17858;
wire      [7:0] n17859;
wire      [7:0] n1786;
wire      [7:0] n17860;
wire      [7:0] n17861;
wire      [7:0] n17862;
wire      [7:0] n17863;
wire      [7:0] n17864;
wire      [7:0] n17865;
wire      [7:0] n17866;
wire      [7:0] n17867;
wire      [7:0] n17868;
wire      [7:0] n17869;
wire      [7:0] n1787;
wire      [7:0] n17870;
wire      [7:0] n17871;
wire      [7:0] n17872;
wire      [7:0] n17873;
wire      [7:0] n17874;
wire      [7:0] n17875;
wire      [7:0] n17876;
wire      [7:0] n17877;
wire      [7:0] n17878;
wire      [7:0] n17879;
wire      [7:0] n1788;
wire      [7:0] n17880;
wire      [7:0] n17881;
wire      [7:0] n17882;
wire      [7:0] n17883;
wire      [7:0] n17884;
wire      [7:0] n17885;
wire      [7:0] n17886;
wire      [7:0] n17887;
wire      [7:0] n17888;
wire      [7:0] n17889;
wire      [7:0] n1789;
wire      [7:0] n17890;
wire      [7:0] n17891;
wire      [7:0] n17892;
wire      [7:0] n17893;
wire      [7:0] n17894;
wire      [7:0] n17895;
wire      [7:0] n17896;
wire      [7:0] n17897;
wire      [7:0] n17898;
wire      [7:0] n17899;
wire            n179;
wire      [7:0] n1790;
wire      [7:0] n17900;
wire      [7:0] n17901;
wire      [7:0] n17902;
wire      [7:0] n17903;
wire      [7:0] n17904;
wire      [7:0] n17905;
wire      [7:0] n17906;
wire      [7:0] n17907;
wire      [7:0] n17908;
wire      [7:0] n17909;
wire      [7:0] n1791;
wire      [7:0] n17910;
wire      [7:0] n17911;
wire      [7:0] n17912;
wire      [7:0] n17913;
wire      [7:0] n17914;
wire      [7:0] n17915;
wire      [7:0] n17916;
wire      [7:0] n17917;
wire      [7:0] n17918;
wire      [7:0] n17919;
wire      [7:0] n1792;
wire      [7:0] n17920;
wire      [7:0] n17921;
wire      [7:0] n17922;
wire      [7:0] n17923;
wire      [7:0] n17924;
wire      [7:0] n17925;
wire      [7:0] n17926;
wire      [7:0] n17927;
wire      [7:0] n17928;
wire      [7:0] n17929;
wire      [7:0] n1793;
wire      [7:0] n17930;
wire      [7:0] n17931;
wire      [7:0] n17932;
wire      [7:0] n17933;
wire      [7:0] n17934;
wire      [7:0] n17935;
wire      [7:0] n17936;
wire      [7:0] n17937;
wire      [7:0] n17938;
wire      [7:0] n17939;
wire      [7:0] n1794;
wire      [7:0] n17940;
wire      [7:0] n17941;
wire      [7:0] n17942;
wire      [7:0] n17943;
wire      [7:0] n17944;
wire      [7:0] n17945;
wire      [7:0] n17946;
wire      [7:0] n17947;
wire      [7:0] n17948;
wire      [7:0] n17949;
wire      [7:0] n1795;
wire      [7:0] n17950;
wire      [7:0] n17951;
wire      [7:0] n17952;
wire      [7:0] n17953;
wire      [7:0] n17954;
wire      [7:0] n17955;
wire      [7:0] n17956;
wire      [7:0] n17957;
wire      [7:0] n17958;
wire      [7:0] n17959;
wire            n1796;
wire      [7:0] n17960;
wire      [7:0] n17961;
wire      [7:0] n17962;
wire      [7:0] n17963;
wire      [7:0] n17964;
wire      [7:0] n17965;
wire      [7:0] n17966;
wire      [7:0] n17967;
wire      [7:0] n17968;
wire      [7:0] n17969;
wire      [7:0] n1797;
wire      [7:0] n17970;
wire      [7:0] n17971;
wire      [7:0] n17972;
wire      [7:0] n17973;
wire      [7:0] n17974;
wire      [7:0] n17975;
wire      [7:0] n17976;
wire      [7:0] n17977;
wire      [7:0] n17978;
wire      [7:0] n17979;
wire            n1798;
wire      [7:0] n17980;
wire      [7:0] n17981;
wire      [7:0] n17982;
wire      [7:0] n17983;
wire      [7:0] n17984;
wire      [7:0] n17985;
wire      [7:0] n17986;
wire      [7:0] n17987;
wire      [7:0] n17988;
wire      [7:0] n17989;
wire      [7:0] n1799;
wire     [79:0] n17990;
wire      [7:0] n17991;
wire      [7:0] n17992;
wire            n17993;
wire      [7:0] n17994;
wire            n17995;
wire      [7:0] n17996;
wire            n17997;
wire      [7:0] n17998;
wire            n17999;
wire      [7:0] n18;
wire            n1800;
wire      [7:0] n18000;
wire            n18001;
wire      [7:0] n18002;
wire            n18003;
wire      [7:0] n18004;
wire            n18005;
wire      [7:0] n18006;
wire            n18007;
wire      [7:0] n18008;
wire            n18009;
wire      [7:0] n1801;
wire      [7:0] n18010;
wire            n18011;
wire      [7:0] n18012;
wire            n18013;
wire      [7:0] n18014;
wire            n18015;
wire      [7:0] n18016;
wire            n18017;
wire      [7:0] n18018;
wire            n18019;
wire            n1802;
wire      [7:0] n18020;
wire            n18021;
wire      [7:0] n18022;
wire            n18023;
wire      [7:0] n18024;
wire            n18025;
wire      [7:0] n18026;
wire            n18027;
wire      [7:0] n18028;
wire            n18029;
wire      [7:0] n1803;
wire      [7:0] n18030;
wire            n18031;
wire      [7:0] n18032;
wire            n18033;
wire      [7:0] n18034;
wire            n18035;
wire      [7:0] n18036;
wire            n18037;
wire      [7:0] n18038;
wire            n18039;
wire            n1804;
wire      [7:0] n18040;
wire            n18041;
wire      [7:0] n18042;
wire            n18043;
wire      [7:0] n18044;
wire            n18045;
wire      [7:0] n18046;
wire            n18047;
wire      [7:0] n18048;
wire            n18049;
wire      [7:0] n1805;
wire      [7:0] n18050;
wire            n18051;
wire      [7:0] n18052;
wire            n18053;
wire      [7:0] n18054;
wire            n18055;
wire      [7:0] n18056;
wire            n18057;
wire      [7:0] n18058;
wire            n18059;
wire            n1806;
wire      [7:0] n18060;
wire            n18061;
wire      [7:0] n18062;
wire            n18063;
wire      [7:0] n18064;
wire            n18065;
wire      [7:0] n18066;
wire            n18067;
wire      [7:0] n18068;
wire            n18069;
wire      [7:0] n1807;
wire      [7:0] n18070;
wire            n18071;
wire      [7:0] n18072;
wire            n18073;
wire      [7:0] n18074;
wire            n18075;
wire      [7:0] n18076;
wire            n18077;
wire      [7:0] n18078;
wire            n18079;
wire            n1808;
wire      [7:0] n18080;
wire            n18081;
wire      [7:0] n18082;
wire            n18083;
wire      [7:0] n18084;
wire            n18085;
wire      [7:0] n18086;
wire            n18087;
wire      [7:0] n18088;
wire            n18089;
wire      [7:0] n1809;
wire      [7:0] n18090;
wire            n18091;
wire      [7:0] n18092;
wire            n18093;
wire      [7:0] n18094;
wire            n18095;
wire      [7:0] n18096;
wire            n18097;
wire      [7:0] n18098;
wire            n18099;
wire      [7:0] n181;
wire            n1810;
wire      [7:0] n18100;
wire            n18101;
wire      [7:0] n18102;
wire            n18103;
wire      [7:0] n18104;
wire            n18105;
wire      [7:0] n18106;
wire            n18107;
wire      [7:0] n18108;
wire            n18109;
wire      [7:0] n1811;
wire      [7:0] n18110;
wire            n18111;
wire      [7:0] n18112;
wire            n18113;
wire      [7:0] n18114;
wire            n18115;
wire      [7:0] n18116;
wire            n18117;
wire      [7:0] n18118;
wire            n18119;
wire            n1812;
wire      [7:0] n18120;
wire            n18121;
wire      [7:0] n18122;
wire            n18123;
wire      [7:0] n18124;
wire            n18125;
wire      [7:0] n18126;
wire            n18127;
wire      [7:0] n18128;
wire            n18129;
wire      [7:0] n1813;
wire      [7:0] n18130;
wire            n18131;
wire      [7:0] n18132;
wire            n18133;
wire      [7:0] n18134;
wire            n18135;
wire      [7:0] n18136;
wire            n18137;
wire      [7:0] n18138;
wire            n18139;
wire            n1814;
wire      [7:0] n18140;
wire            n18141;
wire      [7:0] n18142;
wire            n18143;
wire      [7:0] n18144;
wire            n18145;
wire      [7:0] n18146;
wire            n18147;
wire      [7:0] n18148;
wire            n18149;
wire      [7:0] n1815;
wire      [7:0] n18150;
wire            n18151;
wire      [7:0] n18152;
wire            n18153;
wire      [7:0] n18154;
wire            n18155;
wire      [7:0] n18156;
wire            n18157;
wire      [7:0] n18158;
wire            n18159;
wire            n1816;
wire      [7:0] n18160;
wire            n18161;
wire      [7:0] n18162;
wire            n18163;
wire      [7:0] n18164;
wire            n18165;
wire      [7:0] n18166;
wire            n18167;
wire      [7:0] n18168;
wire            n18169;
wire      [7:0] n1817;
wire      [7:0] n18170;
wire            n18171;
wire      [7:0] n18172;
wire            n18173;
wire      [7:0] n18174;
wire            n18175;
wire      [7:0] n18176;
wire            n18177;
wire      [7:0] n18178;
wire            n18179;
wire            n1818;
wire      [7:0] n18180;
wire            n18181;
wire      [7:0] n18182;
wire            n18183;
wire      [7:0] n18184;
wire            n18185;
wire      [7:0] n18186;
wire            n18187;
wire      [7:0] n18188;
wire            n18189;
wire      [7:0] n1819;
wire      [7:0] n18190;
wire            n18191;
wire      [7:0] n18192;
wire            n18193;
wire      [7:0] n18194;
wire            n18195;
wire      [7:0] n18196;
wire            n18197;
wire      [7:0] n18198;
wire            n18199;
wire            n1820;
wire      [7:0] n18200;
wire            n18201;
wire      [7:0] n18202;
wire            n18203;
wire      [7:0] n18204;
wire            n18205;
wire      [7:0] n18206;
wire            n18207;
wire      [7:0] n18208;
wire            n18209;
wire      [7:0] n1821;
wire      [7:0] n18210;
wire            n18211;
wire      [7:0] n18212;
wire            n18213;
wire      [7:0] n18214;
wire            n18215;
wire      [7:0] n18216;
wire            n18217;
wire      [7:0] n18218;
wire            n18219;
wire            n1822;
wire      [7:0] n18220;
wire            n18221;
wire      [7:0] n18222;
wire            n18223;
wire      [7:0] n18224;
wire            n18225;
wire      [7:0] n18226;
wire            n18227;
wire      [7:0] n18228;
wire            n18229;
wire      [7:0] n1823;
wire      [7:0] n18230;
wire            n18231;
wire      [7:0] n18232;
wire            n18233;
wire      [7:0] n18234;
wire            n18235;
wire      [7:0] n18236;
wire            n18237;
wire      [7:0] n18238;
wire            n18239;
wire            n1824;
wire      [7:0] n18240;
wire            n18241;
wire      [7:0] n18242;
wire            n18243;
wire      [7:0] n18244;
wire            n18245;
wire      [7:0] n18246;
wire            n18247;
wire      [7:0] n18248;
wire            n18249;
wire      [7:0] n1825;
wire      [7:0] n18250;
wire            n18251;
wire      [7:0] n18252;
wire            n18253;
wire      [7:0] n18254;
wire            n18255;
wire      [7:0] n18256;
wire            n18257;
wire      [7:0] n18258;
wire            n18259;
wire            n1826;
wire      [7:0] n18260;
wire            n18261;
wire      [7:0] n18262;
wire            n18263;
wire      [7:0] n18264;
wire            n18265;
wire      [7:0] n18266;
wire            n18267;
wire      [7:0] n18268;
wire            n18269;
wire      [7:0] n1827;
wire      [7:0] n18270;
wire            n18271;
wire      [7:0] n18272;
wire            n18273;
wire      [7:0] n18274;
wire            n18275;
wire      [7:0] n18276;
wire            n18277;
wire      [7:0] n18278;
wire            n18279;
wire            n1828;
wire      [7:0] n18280;
wire            n18281;
wire      [7:0] n18282;
wire            n18283;
wire      [7:0] n18284;
wire            n18285;
wire      [7:0] n18286;
wire            n18287;
wire      [7:0] n18288;
wire            n18289;
wire      [7:0] n1829;
wire      [7:0] n18290;
wire            n18291;
wire      [7:0] n18292;
wire            n18293;
wire      [7:0] n18294;
wire            n18295;
wire      [7:0] n18296;
wire            n18297;
wire      [7:0] n18298;
wire            n18299;
wire            n183;
wire            n1830;
wire      [7:0] n18300;
wire            n18301;
wire      [7:0] n18302;
wire            n18303;
wire      [7:0] n18304;
wire            n18305;
wire      [7:0] n18306;
wire            n18307;
wire      [7:0] n18308;
wire            n18309;
wire      [7:0] n1831;
wire      [7:0] n18310;
wire            n18311;
wire      [7:0] n18312;
wire            n18313;
wire      [7:0] n18314;
wire            n18315;
wire      [7:0] n18316;
wire            n18317;
wire      [7:0] n18318;
wire            n18319;
wire            n1832;
wire      [7:0] n18320;
wire            n18321;
wire      [7:0] n18322;
wire            n18323;
wire      [7:0] n18324;
wire            n18325;
wire      [7:0] n18326;
wire            n18327;
wire      [7:0] n18328;
wire            n18329;
wire      [7:0] n1833;
wire      [7:0] n18330;
wire            n18331;
wire      [7:0] n18332;
wire            n18333;
wire      [7:0] n18334;
wire            n18335;
wire      [7:0] n18336;
wire            n18337;
wire      [7:0] n18338;
wire            n18339;
wire            n1834;
wire      [7:0] n18340;
wire            n18341;
wire      [7:0] n18342;
wire            n18343;
wire      [7:0] n18344;
wire            n18345;
wire      [7:0] n18346;
wire            n18347;
wire      [7:0] n18348;
wire            n18349;
wire      [7:0] n1835;
wire      [7:0] n18350;
wire            n18351;
wire      [7:0] n18352;
wire            n18353;
wire      [7:0] n18354;
wire            n18355;
wire      [7:0] n18356;
wire            n18357;
wire      [7:0] n18358;
wire            n18359;
wire            n1836;
wire      [7:0] n18360;
wire            n18361;
wire      [7:0] n18362;
wire            n18363;
wire      [7:0] n18364;
wire            n18365;
wire      [7:0] n18366;
wire            n18367;
wire      [7:0] n18368;
wire            n18369;
wire      [7:0] n1837;
wire      [7:0] n18370;
wire            n18371;
wire      [7:0] n18372;
wire            n18373;
wire      [7:0] n18374;
wire            n18375;
wire      [7:0] n18376;
wire            n18377;
wire      [7:0] n18378;
wire            n18379;
wire            n1838;
wire      [7:0] n18380;
wire            n18381;
wire      [7:0] n18382;
wire            n18383;
wire      [7:0] n18384;
wire            n18385;
wire      [7:0] n18386;
wire            n18387;
wire      [7:0] n18388;
wire            n18389;
wire      [7:0] n1839;
wire      [7:0] n18390;
wire            n18391;
wire      [7:0] n18392;
wire            n18393;
wire      [7:0] n18394;
wire            n18395;
wire      [7:0] n18396;
wire            n18397;
wire      [7:0] n18398;
wire            n18399;
wire            n1840;
wire      [7:0] n18400;
wire            n18401;
wire      [7:0] n18402;
wire            n18403;
wire      [7:0] n18404;
wire            n18405;
wire      [7:0] n18406;
wire            n18407;
wire      [7:0] n18408;
wire            n18409;
wire      [7:0] n1841;
wire      [7:0] n18410;
wire            n18411;
wire      [7:0] n18412;
wire            n18413;
wire      [7:0] n18414;
wire            n18415;
wire      [7:0] n18416;
wire            n18417;
wire      [7:0] n18418;
wire            n18419;
wire            n1842;
wire      [7:0] n18420;
wire            n18421;
wire      [7:0] n18422;
wire            n18423;
wire      [7:0] n18424;
wire            n18425;
wire      [7:0] n18426;
wire            n18427;
wire      [7:0] n18428;
wire            n18429;
wire      [7:0] n1843;
wire      [7:0] n18430;
wire            n18431;
wire      [7:0] n18432;
wire            n18433;
wire      [7:0] n18434;
wire            n18435;
wire      [7:0] n18436;
wire            n18437;
wire      [7:0] n18438;
wire            n18439;
wire            n1844;
wire      [7:0] n18440;
wire            n18441;
wire      [7:0] n18442;
wire            n18443;
wire      [7:0] n18444;
wire            n18445;
wire      [7:0] n18446;
wire            n18447;
wire      [7:0] n18448;
wire            n18449;
wire      [7:0] n1845;
wire      [7:0] n18450;
wire            n18451;
wire      [7:0] n18452;
wire            n18453;
wire      [7:0] n18454;
wire            n18455;
wire      [7:0] n18456;
wire            n18457;
wire      [7:0] n18458;
wire            n18459;
wire            n1846;
wire      [7:0] n18460;
wire            n18461;
wire      [7:0] n18462;
wire            n18463;
wire      [7:0] n18464;
wire            n18465;
wire      [7:0] n18466;
wire            n18467;
wire      [7:0] n18468;
wire            n18469;
wire      [7:0] n1847;
wire      [7:0] n18470;
wire            n18471;
wire      [7:0] n18472;
wire            n18473;
wire      [7:0] n18474;
wire            n18475;
wire      [7:0] n18476;
wire            n18477;
wire      [7:0] n18478;
wire            n18479;
wire            n1848;
wire      [7:0] n18480;
wire            n18481;
wire      [7:0] n18482;
wire            n18483;
wire      [7:0] n18484;
wire            n18485;
wire      [7:0] n18486;
wire            n18487;
wire      [7:0] n18488;
wire            n18489;
wire      [7:0] n1849;
wire      [7:0] n18490;
wire            n18491;
wire      [7:0] n18492;
wire            n18493;
wire      [7:0] n18494;
wire            n18495;
wire      [7:0] n18496;
wire            n18497;
wire      [7:0] n18498;
wire            n18499;
wire      [7:0] n185;
wire            n1850;
wire      [7:0] n18500;
wire            n18501;
wire      [7:0] n18502;
wire            n18503;
wire      [7:0] n18504;
wire      [7:0] n18505;
wire      [7:0] n18506;
wire      [7:0] n18507;
wire      [7:0] n18508;
wire      [7:0] n18509;
wire      [7:0] n1851;
wire      [7:0] n18510;
wire      [7:0] n18511;
wire      [7:0] n18512;
wire      [7:0] n18513;
wire      [7:0] n18514;
wire      [7:0] n18515;
wire      [7:0] n18516;
wire      [7:0] n18517;
wire      [7:0] n18518;
wire      [7:0] n18519;
wire            n1852;
wire      [7:0] n18520;
wire      [7:0] n18521;
wire      [7:0] n18522;
wire      [7:0] n18523;
wire      [7:0] n18524;
wire      [7:0] n18525;
wire      [7:0] n18526;
wire      [7:0] n18527;
wire      [7:0] n18528;
wire      [7:0] n18529;
wire      [7:0] n1853;
wire      [7:0] n18530;
wire      [7:0] n18531;
wire      [7:0] n18532;
wire      [7:0] n18533;
wire      [7:0] n18534;
wire      [7:0] n18535;
wire      [7:0] n18536;
wire      [7:0] n18537;
wire      [7:0] n18538;
wire      [7:0] n18539;
wire            n1854;
wire      [7:0] n18540;
wire      [7:0] n18541;
wire      [7:0] n18542;
wire      [7:0] n18543;
wire      [7:0] n18544;
wire      [7:0] n18545;
wire      [7:0] n18546;
wire      [7:0] n18547;
wire      [7:0] n18548;
wire      [7:0] n18549;
wire      [7:0] n1855;
wire      [7:0] n18550;
wire      [7:0] n18551;
wire      [7:0] n18552;
wire      [7:0] n18553;
wire      [7:0] n18554;
wire      [7:0] n18555;
wire      [7:0] n18556;
wire      [7:0] n18557;
wire      [7:0] n18558;
wire      [7:0] n18559;
wire            n1856;
wire      [7:0] n18560;
wire      [7:0] n18561;
wire      [7:0] n18562;
wire      [7:0] n18563;
wire      [7:0] n18564;
wire      [7:0] n18565;
wire      [7:0] n18566;
wire      [7:0] n18567;
wire      [7:0] n18568;
wire      [7:0] n18569;
wire      [7:0] n1857;
wire      [7:0] n18570;
wire      [7:0] n18571;
wire      [7:0] n18572;
wire      [7:0] n18573;
wire      [7:0] n18574;
wire      [7:0] n18575;
wire      [7:0] n18576;
wire      [7:0] n18577;
wire      [7:0] n18578;
wire      [7:0] n18579;
wire            n1858;
wire      [7:0] n18580;
wire      [7:0] n18581;
wire      [7:0] n18582;
wire      [7:0] n18583;
wire      [7:0] n18584;
wire      [7:0] n18585;
wire      [7:0] n18586;
wire      [7:0] n18587;
wire      [7:0] n18588;
wire      [7:0] n18589;
wire      [7:0] n1859;
wire      [7:0] n18590;
wire      [7:0] n18591;
wire      [7:0] n18592;
wire      [7:0] n18593;
wire      [7:0] n18594;
wire      [7:0] n18595;
wire      [7:0] n18596;
wire      [7:0] n18597;
wire      [7:0] n18598;
wire      [7:0] n18599;
wire            n186;
wire            n1860;
wire      [7:0] n18600;
wire      [7:0] n18601;
wire      [7:0] n18602;
wire      [7:0] n18603;
wire      [7:0] n18604;
wire      [7:0] n18605;
wire      [7:0] n18606;
wire      [7:0] n18607;
wire      [7:0] n18608;
wire      [7:0] n18609;
wire      [7:0] n1861;
wire      [7:0] n18610;
wire      [7:0] n18611;
wire      [7:0] n18612;
wire      [7:0] n18613;
wire      [7:0] n18614;
wire      [7:0] n18615;
wire      [7:0] n18616;
wire      [7:0] n18617;
wire      [7:0] n18618;
wire      [7:0] n18619;
wire            n1862;
wire      [7:0] n18620;
wire      [7:0] n18621;
wire      [7:0] n18622;
wire      [7:0] n18623;
wire      [7:0] n18624;
wire      [7:0] n18625;
wire      [7:0] n18626;
wire      [7:0] n18627;
wire      [7:0] n18628;
wire      [7:0] n18629;
wire      [7:0] n1863;
wire      [7:0] n18630;
wire      [7:0] n18631;
wire      [7:0] n18632;
wire      [7:0] n18633;
wire      [7:0] n18634;
wire      [7:0] n18635;
wire      [7:0] n18636;
wire      [7:0] n18637;
wire      [7:0] n18638;
wire      [7:0] n18639;
wire            n1864;
wire      [7:0] n18640;
wire      [7:0] n18641;
wire      [7:0] n18642;
wire      [7:0] n18643;
wire      [7:0] n18644;
wire      [7:0] n18645;
wire      [7:0] n18646;
wire      [7:0] n18647;
wire      [7:0] n18648;
wire      [7:0] n18649;
wire      [7:0] n1865;
wire      [7:0] n18650;
wire      [7:0] n18651;
wire      [7:0] n18652;
wire      [7:0] n18653;
wire      [7:0] n18654;
wire      [7:0] n18655;
wire      [7:0] n18656;
wire      [7:0] n18657;
wire      [7:0] n18658;
wire      [7:0] n18659;
wire            n1866;
wire      [7:0] n18660;
wire      [7:0] n18661;
wire      [7:0] n18662;
wire      [7:0] n18663;
wire      [7:0] n18664;
wire      [7:0] n18665;
wire      [7:0] n18666;
wire      [7:0] n18667;
wire      [7:0] n18668;
wire      [7:0] n18669;
wire      [7:0] n1867;
wire      [7:0] n18670;
wire      [7:0] n18671;
wire      [7:0] n18672;
wire      [7:0] n18673;
wire      [7:0] n18674;
wire      [7:0] n18675;
wire      [7:0] n18676;
wire      [7:0] n18677;
wire      [7:0] n18678;
wire      [7:0] n18679;
wire            n1868;
wire      [7:0] n18680;
wire      [7:0] n18681;
wire      [7:0] n18682;
wire      [7:0] n18683;
wire      [7:0] n18684;
wire      [7:0] n18685;
wire      [7:0] n18686;
wire      [7:0] n18687;
wire      [7:0] n18688;
wire      [7:0] n18689;
wire      [7:0] n1869;
wire      [7:0] n18690;
wire      [7:0] n18691;
wire      [7:0] n18692;
wire      [7:0] n18693;
wire      [7:0] n18694;
wire      [7:0] n18695;
wire      [7:0] n18696;
wire      [7:0] n18697;
wire      [7:0] n18698;
wire      [7:0] n18699;
wire      [7:0] n187;
wire            n1870;
wire      [7:0] n18700;
wire      [7:0] n18701;
wire      [7:0] n18702;
wire      [7:0] n18703;
wire      [7:0] n18704;
wire      [7:0] n18705;
wire      [7:0] n18706;
wire      [7:0] n18707;
wire      [7:0] n18708;
wire      [7:0] n18709;
wire      [7:0] n1871;
wire      [7:0] n18710;
wire      [7:0] n18711;
wire      [7:0] n18712;
wire      [7:0] n18713;
wire      [7:0] n18714;
wire      [7:0] n18715;
wire      [7:0] n18716;
wire      [7:0] n18717;
wire      [7:0] n18718;
wire      [7:0] n18719;
wire            n1872;
wire      [7:0] n18720;
wire      [7:0] n18721;
wire      [7:0] n18722;
wire      [7:0] n18723;
wire      [7:0] n18724;
wire      [7:0] n18725;
wire      [7:0] n18726;
wire      [7:0] n18727;
wire      [7:0] n18728;
wire      [7:0] n18729;
wire      [7:0] n1873;
wire      [7:0] n18730;
wire      [7:0] n18731;
wire      [7:0] n18732;
wire      [7:0] n18733;
wire      [7:0] n18734;
wire      [7:0] n18735;
wire      [7:0] n18736;
wire      [7:0] n18737;
wire      [7:0] n18738;
wire      [7:0] n18739;
wire            n1874;
wire      [7:0] n18740;
wire      [7:0] n18741;
wire      [7:0] n18742;
wire      [7:0] n18743;
wire      [7:0] n18744;
wire      [7:0] n18745;
wire      [7:0] n18746;
wire      [7:0] n18747;
wire      [7:0] n18748;
wire      [7:0] n18749;
wire      [7:0] n1875;
wire      [7:0] n18750;
wire      [7:0] n18751;
wire      [7:0] n18752;
wire      [7:0] n18753;
wire      [7:0] n18754;
wire      [7:0] n18755;
wire      [7:0] n18756;
wire      [7:0] n18757;
wire      [7:0] n18758;
wire      [7:0] n18759;
wire            n1876;
wire      [7:0] n18760;
wire      [7:0] n18761;
wire      [7:0] n18762;
wire      [7:0] n18763;
wire      [7:0] n18764;
wire     [87:0] n18765;
wire      [7:0] n18766;
wire      [7:0] n18767;
wire      [7:0] n18768;
wire      [7:0] n18769;
wire      [7:0] n1877;
wire      [7:0] n18770;
wire      [7:0] n18771;
wire     [95:0] n18772;
wire      [7:0] n18773;
wire            n18774;
wire      [7:0] n18775;
wire            n18776;
wire      [7:0] n18777;
wire            n18778;
wire      [7:0] n18779;
wire            n1878;
wire            n18780;
wire      [7:0] n18781;
wire            n18782;
wire      [7:0] n18783;
wire            n18784;
wire      [7:0] n18785;
wire            n18786;
wire      [7:0] n18787;
wire            n18788;
wire      [7:0] n18789;
wire      [7:0] n1879;
wire            n18790;
wire      [7:0] n18791;
wire            n18792;
wire      [7:0] n18793;
wire            n18794;
wire      [7:0] n18795;
wire            n18796;
wire      [7:0] n18797;
wire            n18798;
wire      [7:0] n18799;
wire            n1880;
wire            n18800;
wire      [7:0] n18801;
wire            n18802;
wire      [7:0] n18803;
wire            n18804;
wire      [7:0] n18805;
wire            n18806;
wire      [7:0] n18807;
wire            n18808;
wire      [7:0] n18809;
wire      [7:0] n1881;
wire            n18810;
wire      [7:0] n18811;
wire            n18812;
wire      [7:0] n18813;
wire            n18814;
wire      [7:0] n18815;
wire            n18816;
wire      [7:0] n18817;
wire            n18818;
wire      [7:0] n18819;
wire            n1882;
wire            n18820;
wire      [7:0] n18821;
wire            n18822;
wire      [7:0] n18823;
wire            n18824;
wire      [7:0] n18825;
wire            n18826;
wire      [7:0] n18827;
wire            n18828;
wire      [7:0] n18829;
wire      [7:0] n1883;
wire            n18830;
wire      [7:0] n18831;
wire            n18832;
wire      [7:0] n18833;
wire            n18834;
wire      [7:0] n18835;
wire            n18836;
wire      [7:0] n18837;
wire            n18838;
wire      [7:0] n18839;
wire            n1884;
wire            n18840;
wire      [7:0] n18841;
wire            n18842;
wire      [7:0] n18843;
wire            n18844;
wire      [7:0] n18845;
wire            n18846;
wire      [7:0] n18847;
wire            n18848;
wire      [7:0] n18849;
wire      [7:0] n1885;
wire            n18850;
wire      [7:0] n18851;
wire            n18852;
wire      [7:0] n18853;
wire            n18854;
wire      [7:0] n18855;
wire            n18856;
wire      [7:0] n18857;
wire            n18858;
wire      [7:0] n18859;
wire            n1886;
wire            n18860;
wire      [7:0] n18861;
wire            n18862;
wire      [7:0] n18863;
wire            n18864;
wire      [7:0] n18865;
wire            n18866;
wire      [7:0] n18867;
wire            n18868;
wire      [7:0] n18869;
wire      [7:0] n1887;
wire            n18870;
wire      [7:0] n18871;
wire            n18872;
wire      [7:0] n18873;
wire            n18874;
wire      [7:0] n18875;
wire            n18876;
wire      [7:0] n18877;
wire            n18878;
wire      [7:0] n18879;
wire            n1888;
wire            n18880;
wire      [7:0] n18881;
wire            n18882;
wire      [7:0] n18883;
wire            n18884;
wire      [7:0] n18885;
wire            n18886;
wire      [7:0] n18887;
wire            n18888;
wire      [7:0] n18889;
wire      [7:0] n1889;
wire            n18890;
wire      [7:0] n18891;
wire            n18892;
wire      [7:0] n18893;
wire            n18894;
wire      [7:0] n18895;
wire            n18896;
wire      [7:0] n18897;
wire            n18898;
wire      [7:0] n18899;
wire            n189;
wire            n1890;
wire            n18900;
wire      [7:0] n18901;
wire            n18902;
wire      [7:0] n18903;
wire            n18904;
wire      [7:0] n18905;
wire            n18906;
wire      [7:0] n18907;
wire            n18908;
wire      [7:0] n18909;
wire      [7:0] n1891;
wire            n18910;
wire      [7:0] n18911;
wire            n18912;
wire      [7:0] n18913;
wire            n18914;
wire      [7:0] n18915;
wire            n18916;
wire      [7:0] n18917;
wire            n18918;
wire      [7:0] n18919;
wire            n1892;
wire            n18920;
wire      [7:0] n18921;
wire            n18922;
wire      [7:0] n18923;
wire            n18924;
wire      [7:0] n18925;
wire            n18926;
wire      [7:0] n18927;
wire            n18928;
wire      [7:0] n18929;
wire      [7:0] n1893;
wire            n18930;
wire      [7:0] n18931;
wire            n18932;
wire      [7:0] n18933;
wire            n18934;
wire      [7:0] n18935;
wire            n18936;
wire      [7:0] n18937;
wire            n18938;
wire      [7:0] n18939;
wire            n1894;
wire            n18940;
wire      [7:0] n18941;
wire            n18942;
wire      [7:0] n18943;
wire            n18944;
wire      [7:0] n18945;
wire            n18946;
wire      [7:0] n18947;
wire            n18948;
wire      [7:0] n18949;
wire      [7:0] n1895;
wire            n18950;
wire      [7:0] n18951;
wire            n18952;
wire      [7:0] n18953;
wire            n18954;
wire      [7:0] n18955;
wire            n18956;
wire      [7:0] n18957;
wire            n18958;
wire      [7:0] n18959;
wire            n1896;
wire            n18960;
wire      [7:0] n18961;
wire            n18962;
wire      [7:0] n18963;
wire            n18964;
wire      [7:0] n18965;
wire            n18966;
wire      [7:0] n18967;
wire            n18968;
wire      [7:0] n18969;
wire      [7:0] n1897;
wire            n18970;
wire      [7:0] n18971;
wire            n18972;
wire      [7:0] n18973;
wire            n18974;
wire      [7:0] n18975;
wire            n18976;
wire      [7:0] n18977;
wire            n18978;
wire      [7:0] n18979;
wire            n1898;
wire            n18980;
wire      [7:0] n18981;
wire            n18982;
wire      [7:0] n18983;
wire            n18984;
wire      [7:0] n18985;
wire            n18986;
wire      [7:0] n18987;
wire            n18988;
wire      [7:0] n18989;
wire      [7:0] n1899;
wire            n18990;
wire      [7:0] n18991;
wire            n18992;
wire      [7:0] n18993;
wire            n18994;
wire      [7:0] n18995;
wire            n18996;
wire      [7:0] n18997;
wire            n18998;
wire      [7:0] n18999;
wire            n1900;
wire            n19000;
wire      [7:0] n19001;
wire            n19002;
wire      [7:0] n19003;
wire            n19004;
wire      [7:0] n19005;
wire            n19006;
wire      [7:0] n19007;
wire            n19008;
wire      [7:0] n19009;
wire      [7:0] n1901;
wire            n19010;
wire      [7:0] n19011;
wire            n19012;
wire      [7:0] n19013;
wire            n19014;
wire      [7:0] n19015;
wire            n19016;
wire      [7:0] n19017;
wire            n19018;
wire      [7:0] n19019;
wire            n1902;
wire            n19020;
wire      [7:0] n19021;
wire            n19022;
wire      [7:0] n19023;
wire            n19024;
wire      [7:0] n19025;
wire            n19026;
wire      [7:0] n19027;
wire            n19028;
wire      [7:0] n19029;
wire      [7:0] n1903;
wire            n19030;
wire      [7:0] n19031;
wire            n19032;
wire      [7:0] n19033;
wire            n19034;
wire      [7:0] n19035;
wire            n19036;
wire      [7:0] n19037;
wire            n19038;
wire      [7:0] n19039;
wire            n1904;
wire            n19040;
wire      [7:0] n19041;
wire            n19042;
wire      [7:0] n19043;
wire            n19044;
wire      [7:0] n19045;
wire            n19046;
wire      [7:0] n19047;
wire            n19048;
wire      [7:0] n19049;
wire      [7:0] n1905;
wire            n19050;
wire      [7:0] n19051;
wire            n19052;
wire      [7:0] n19053;
wire            n19054;
wire      [7:0] n19055;
wire            n19056;
wire      [7:0] n19057;
wire            n19058;
wire      [7:0] n19059;
wire            n1906;
wire            n19060;
wire      [7:0] n19061;
wire            n19062;
wire      [7:0] n19063;
wire            n19064;
wire      [7:0] n19065;
wire            n19066;
wire      [7:0] n19067;
wire            n19068;
wire      [7:0] n19069;
wire      [7:0] n1907;
wire            n19070;
wire      [7:0] n19071;
wire            n19072;
wire      [7:0] n19073;
wire            n19074;
wire      [7:0] n19075;
wire            n19076;
wire      [7:0] n19077;
wire            n19078;
wire      [7:0] n19079;
wire            n1908;
wire            n19080;
wire      [7:0] n19081;
wire            n19082;
wire      [7:0] n19083;
wire            n19084;
wire      [7:0] n19085;
wire            n19086;
wire      [7:0] n19087;
wire            n19088;
wire      [7:0] n19089;
wire      [7:0] n1909;
wire            n19090;
wire      [7:0] n19091;
wire            n19092;
wire      [7:0] n19093;
wire            n19094;
wire      [7:0] n19095;
wire            n19096;
wire      [7:0] n19097;
wire            n19098;
wire      [7:0] n19099;
wire      [7:0] n191;
wire            n1910;
wire            n19100;
wire      [7:0] n19101;
wire            n19102;
wire      [7:0] n19103;
wire            n19104;
wire      [7:0] n19105;
wire            n19106;
wire      [7:0] n19107;
wire            n19108;
wire      [7:0] n19109;
wire      [7:0] n1911;
wire            n19110;
wire      [7:0] n19111;
wire            n19112;
wire      [7:0] n19113;
wire            n19114;
wire      [7:0] n19115;
wire            n19116;
wire      [7:0] n19117;
wire            n19118;
wire      [7:0] n19119;
wire            n1912;
wire            n19120;
wire      [7:0] n19121;
wire            n19122;
wire      [7:0] n19123;
wire            n19124;
wire      [7:0] n19125;
wire            n19126;
wire      [7:0] n19127;
wire            n19128;
wire      [7:0] n19129;
wire      [7:0] n1913;
wire            n19130;
wire      [7:0] n19131;
wire            n19132;
wire      [7:0] n19133;
wire            n19134;
wire      [7:0] n19135;
wire            n19136;
wire      [7:0] n19137;
wire            n19138;
wire      [7:0] n19139;
wire            n1914;
wire            n19140;
wire      [7:0] n19141;
wire            n19142;
wire      [7:0] n19143;
wire            n19144;
wire      [7:0] n19145;
wire            n19146;
wire      [7:0] n19147;
wire            n19148;
wire      [7:0] n19149;
wire      [7:0] n1915;
wire            n19150;
wire      [7:0] n19151;
wire            n19152;
wire      [7:0] n19153;
wire            n19154;
wire      [7:0] n19155;
wire            n19156;
wire      [7:0] n19157;
wire            n19158;
wire      [7:0] n19159;
wire            n1916;
wire            n19160;
wire      [7:0] n19161;
wire            n19162;
wire      [7:0] n19163;
wire            n19164;
wire      [7:0] n19165;
wire            n19166;
wire      [7:0] n19167;
wire            n19168;
wire      [7:0] n19169;
wire      [7:0] n1917;
wire            n19170;
wire      [7:0] n19171;
wire            n19172;
wire      [7:0] n19173;
wire            n19174;
wire      [7:0] n19175;
wire            n19176;
wire      [7:0] n19177;
wire            n19178;
wire      [7:0] n19179;
wire            n1918;
wire            n19180;
wire      [7:0] n19181;
wire            n19182;
wire      [7:0] n19183;
wire            n19184;
wire      [7:0] n19185;
wire            n19186;
wire      [7:0] n19187;
wire            n19188;
wire      [7:0] n19189;
wire      [7:0] n1919;
wire            n19190;
wire      [7:0] n19191;
wire            n19192;
wire      [7:0] n19193;
wire            n19194;
wire      [7:0] n19195;
wire            n19196;
wire      [7:0] n19197;
wire            n19198;
wire      [7:0] n19199;
wire            n1920;
wire            n19200;
wire      [7:0] n19201;
wire            n19202;
wire      [7:0] n19203;
wire            n19204;
wire      [7:0] n19205;
wire            n19206;
wire      [7:0] n19207;
wire            n19208;
wire      [7:0] n19209;
wire      [7:0] n1921;
wire            n19210;
wire      [7:0] n19211;
wire            n19212;
wire      [7:0] n19213;
wire            n19214;
wire      [7:0] n19215;
wire            n19216;
wire      [7:0] n19217;
wire            n19218;
wire      [7:0] n19219;
wire            n1922;
wire            n19220;
wire      [7:0] n19221;
wire            n19222;
wire      [7:0] n19223;
wire            n19224;
wire      [7:0] n19225;
wire            n19226;
wire      [7:0] n19227;
wire            n19228;
wire      [7:0] n19229;
wire      [7:0] n1923;
wire            n19230;
wire      [7:0] n19231;
wire            n19232;
wire      [7:0] n19233;
wire            n19234;
wire      [7:0] n19235;
wire            n19236;
wire      [7:0] n19237;
wire            n19238;
wire      [7:0] n19239;
wire            n1924;
wire            n19240;
wire      [7:0] n19241;
wire            n19242;
wire      [7:0] n19243;
wire            n19244;
wire      [7:0] n19245;
wire            n19246;
wire      [7:0] n19247;
wire            n19248;
wire      [7:0] n19249;
wire      [7:0] n1925;
wire            n19250;
wire      [7:0] n19251;
wire            n19252;
wire      [7:0] n19253;
wire            n19254;
wire      [7:0] n19255;
wire            n19256;
wire      [7:0] n19257;
wire            n19258;
wire      [7:0] n19259;
wire            n1926;
wire            n19260;
wire      [7:0] n19261;
wire            n19262;
wire      [7:0] n19263;
wire            n19264;
wire      [7:0] n19265;
wire            n19266;
wire      [7:0] n19267;
wire            n19268;
wire      [7:0] n19269;
wire      [7:0] n1927;
wire            n19270;
wire      [7:0] n19271;
wire            n19272;
wire      [7:0] n19273;
wire            n19274;
wire      [7:0] n19275;
wire            n19276;
wire      [7:0] n19277;
wire            n19278;
wire      [7:0] n19279;
wire            n1928;
wire            n19280;
wire      [7:0] n19281;
wire            n19282;
wire      [7:0] n19283;
wire            n19284;
wire      [7:0] n19285;
wire      [7:0] n19286;
wire      [7:0] n19287;
wire      [7:0] n19288;
wire      [7:0] n19289;
wire      [7:0] n1929;
wire      [7:0] n19290;
wire      [7:0] n19291;
wire      [7:0] n19292;
wire      [7:0] n19293;
wire      [7:0] n19294;
wire      [7:0] n19295;
wire      [7:0] n19296;
wire      [7:0] n19297;
wire      [7:0] n19298;
wire      [7:0] n19299;
wire            n193;
wire            n1930;
wire      [7:0] n19300;
wire      [7:0] n19301;
wire      [7:0] n19302;
wire      [7:0] n19303;
wire      [7:0] n19304;
wire      [7:0] n19305;
wire      [7:0] n19306;
wire      [7:0] n19307;
wire      [7:0] n19308;
wire      [7:0] n19309;
wire      [7:0] n1931;
wire      [7:0] n19310;
wire      [7:0] n19311;
wire      [7:0] n19312;
wire      [7:0] n19313;
wire      [7:0] n19314;
wire      [7:0] n19315;
wire      [7:0] n19316;
wire      [7:0] n19317;
wire      [7:0] n19318;
wire      [7:0] n19319;
wire            n1932;
wire      [7:0] n19320;
wire      [7:0] n19321;
wire      [7:0] n19322;
wire      [7:0] n19323;
wire      [7:0] n19324;
wire      [7:0] n19325;
wire      [7:0] n19326;
wire      [7:0] n19327;
wire      [7:0] n19328;
wire      [7:0] n19329;
wire      [7:0] n1933;
wire      [7:0] n19330;
wire      [7:0] n19331;
wire      [7:0] n19332;
wire      [7:0] n19333;
wire      [7:0] n19334;
wire      [7:0] n19335;
wire      [7:0] n19336;
wire      [7:0] n19337;
wire      [7:0] n19338;
wire      [7:0] n19339;
wire            n1934;
wire      [7:0] n19340;
wire      [7:0] n19341;
wire      [7:0] n19342;
wire      [7:0] n19343;
wire      [7:0] n19344;
wire      [7:0] n19345;
wire      [7:0] n19346;
wire      [7:0] n19347;
wire      [7:0] n19348;
wire      [7:0] n19349;
wire      [7:0] n1935;
wire      [7:0] n19350;
wire      [7:0] n19351;
wire      [7:0] n19352;
wire      [7:0] n19353;
wire      [7:0] n19354;
wire      [7:0] n19355;
wire      [7:0] n19356;
wire      [7:0] n19357;
wire      [7:0] n19358;
wire      [7:0] n19359;
wire            n1936;
wire      [7:0] n19360;
wire      [7:0] n19361;
wire      [7:0] n19362;
wire      [7:0] n19363;
wire      [7:0] n19364;
wire      [7:0] n19365;
wire      [7:0] n19366;
wire      [7:0] n19367;
wire      [7:0] n19368;
wire      [7:0] n19369;
wire      [7:0] n1937;
wire      [7:0] n19370;
wire      [7:0] n19371;
wire      [7:0] n19372;
wire      [7:0] n19373;
wire      [7:0] n19374;
wire      [7:0] n19375;
wire      [7:0] n19376;
wire      [7:0] n19377;
wire      [7:0] n19378;
wire      [7:0] n19379;
wire            n1938;
wire      [7:0] n19380;
wire      [7:0] n19381;
wire      [7:0] n19382;
wire      [7:0] n19383;
wire      [7:0] n19384;
wire      [7:0] n19385;
wire      [7:0] n19386;
wire      [7:0] n19387;
wire      [7:0] n19388;
wire      [7:0] n19389;
wire      [7:0] n1939;
wire      [7:0] n19390;
wire      [7:0] n19391;
wire      [7:0] n19392;
wire      [7:0] n19393;
wire      [7:0] n19394;
wire      [7:0] n19395;
wire      [7:0] n19396;
wire      [7:0] n19397;
wire      [7:0] n19398;
wire      [7:0] n19399;
wire            n1940;
wire      [7:0] n19400;
wire      [7:0] n19401;
wire      [7:0] n19402;
wire      [7:0] n19403;
wire      [7:0] n19404;
wire      [7:0] n19405;
wire      [7:0] n19406;
wire      [7:0] n19407;
wire      [7:0] n19408;
wire      [7:0] n19409;
wire      [7:0] n1941;
wire      [7:0] n19410;
wire      [7:0] n19411;
wire      [7:0] n19412;
wire      [7:0] n19413;
wire      [7:0] n19414;
wire      [7:0] n19415;
wire      [7:0] n19416;
wire      [7:0] n19417;
wire      [7:0] n19418;
wire      [7:0] n19419;
wire            n1942;
wire      [7:0] n19420;
wire      [7:0] n19421;
wire      [7:0] n19422;
wire      [7:0] n19423;
wire      [7:0] n19424;
wire      [7:0] n19425;
wire      [7:0] n19426;
wire      [7:0] n19427;
wire      [7:0] n19428;
wire      [7:0] n19429;
wire      [7:0] n1943;
wire      [7:0] n19430;
wire      [7:0] n19431;
wire      [7:0] n19432;
wire      [7:0] n19433;
wire      [7:0] n19434;
wire      [7:0] n19435;
wire      [7:0] n19436;
wire      [7:0] n19437;
wire      [7:0] n19438;
wire      [7:0] n19439;
wire            n1944;
wire      [7:0] n19440;
wire      [7:0] n19441;
wire      [7:0] n19442;
wire      [7:0] n19443;
wire      [7:0] n19444;
wire      [7:0] n19445;
wire      [7:0] n19446;
wire      [7:0] n19447;
wire      [7:0] n19448;
wire      [7:0] n19449;
wire      [7:0] n1945;
wire      [7:0] n19450;
wire      [7:0] n19451;
wire      [7:0] n19452;
wire      [7:0] n19453;
wire      [7:0] n19454;
wire      [7:0] n19455;
wire      [7:0] n19456;
wire      [7:0] n19457;
wire      [7:0] n19458;
wire      [7:0] n19459;
wire            n1946;
wire      [7:0] n19460;
wire      [7:0] n19461;
wire      [7:0] n19462;
wire      [7:0] n19463;
wire      [7:0] n19464;
wire      [7:0] n19465;
wire      [7:0] n19466;
wire      [7:0] n19467;
wire      [7:0] n19468;
wire      [7:0] n19469;
wire      [7:0] n1947;
wire      [7:0] n19470;
wire      [7:0] n19471;
wire      [7:0] n19472;
wire      [7:0] n19473;
wire      [7:0] n19474;
wire      [7:0] n19475;
wire      [7:0] n19476;
wire      [7:0] n19477;
wire      [7:0] n19478;
wire      [7:0] n19479;
wire            n1948;
wire      [7:0] n19480;
wire      [7:0] n19481;
wire      [7:0] n19482;
wire      [7:0] n19483;
wire      [7:0] n19484;
wire      [7:0] n19485;
wire      [7:0] n19486;
wire      [7:0] n19487;
wire      [7:0] n19488;
wire      [7:0] n19489;
wire      [7:0] n1949;
wire      [7:0] n19490;
wire      [7:0] n19491;
wire      [7:0] n19492;
wire      [7:0] n19493;
wire      [7:0] n19494;
wire      [7:0] n19495;
wire      [7:0] n19496;
wire      [7:0] n19497;
wire      [7:0] n19498;
wire      [7:0] n19499;
wire      [7:0] n195;
wire            n1950;
wire      [7:0] n19500;
wire      [7:0] n19501;
wire      [7:0] n19502;
wire      [7:0] n19503;
wire      [7:0] n19504;
wire      [7:0] n19505;
wire      [7:0] n19506;
wire      [7:0] n19507;
wire      [7:0] n19508;
wire      [7:0] n19509;
wire      [7:0] n1951;
wire      [7:0] n19510;
wire      [7:0] n19511;
wire      [7:0] n19512;
wire      [7:0] n19513;
wire      [7:0] n19514;
wire      [7:0] n19515;
wire      [7:0] n19516;
wire      [7:0] n19517;
wire      [7:0] n19518;
wire      [7:0] n19519;
wire            n1952;
wire      [7:0] n19520;
wire      [7:0] n19521;
wire      [7:0] n19522;
wire      [7:0] n19523;
wire      [7:0] n19524;
wire      [7:0] n19525;
wire      [7:0] n19526;
wire      [7:0] n19527;
wire      [7:0] n19528;
wire      [7:0] n19529;
wire      [7:0] n1953;
wire      [7:0] n19530;
wire      [7:0] n19531;
wire      [7:0] n19532;
wire      [7:0] n19533;
wire      [7:0] n19534;
wire      [7:0] n19535;
wire      [7:0] n19536;
wire      [7:0] n19537;
wire      [7:0] n19538;
wire      [7:0] n19539;
wire            n1954;
wire      [7:0] n19540;
wire      [7:0] n19541;
wire            n19542;
wire      [7:0] n19543;
wire            n19544;
wire      [7:0] n19545;
wire            n19546;
wire      [7:0] n19547;
wire            n19548;
wire      [7:0] n19549;
wire      [7:0] n1955;
wire            n19550;
wire      [7:0] n19551;
wire            n19552;
wire      [7:0] n19553;
wire            n19554;
wire      [7:0] n19555;
wire            n19556;
wire      [7:0] n19557;
wire            n19558;
wire      [7:0] n19559;
wire            n1956;
wire            n19560;
wire      [7:0] n19561;
wire            n19562;
wire      [7:0] n19563;
wire            n19564;
wire      [7:0] n19565;
wire            n19566;
wire      [7:0] n19567;
wire            n19568;
wire      [7:0] n19569;
wire      [7:0] n1957;
wire            n19570;
wire      [7:0] n19571;
wire            n19572;
wire      [7:0] n19573;
wire            n19574;
wire      [7:0] n19575;
wire            n19576;
wire      [7:0] n19577;
wire            n19578;
wire      [7:0] n19579;
wire            n1958;
wire            n19580;
wire      [7:0] n19581;
wire            n19582;
wire      [7:0] n19583;
wire            n19584;
wire      [7:0] n19585;
wire            n19586;
wire      [7:0] n19587;
wire            n19588;
wire      [7:0] n19589;
wire      [7:0] n1959;
wire            n19590;
wire      [7:0] n19591;
wire            n19592;
wire      [7:0] n19593;
wire            n19594;
wire      [7:0] n19595;
wire            n19596;
wire      [7:0] n19597;
wire            n19598;
wire      [7:0] n19599;
wire            n1960;
wire            n19600;
wire      [7:0] n19601;
wire            n19602;
wire      [7:0] n19603;
wire            n19604;
wire      [7:0] n19605;
wire            n19606;
wire      [7:0] n19607;
wire            n19608;
wire      [7:0] n19609;
wire      [7:0] n1961;
wire            n19610;
wire      [7:0] n19611;
wire            n19612;
wire      [7:0] n19613;
wire            n19614;
wire      [7:0] n19615;
wire            n19616;
wire      [7:0] n19617;
wire            n19618;
wire      [7:0] n19619;
wire            n1962;
wire            n19620;
wire      [7:0] n19621;
wire            n19622;
wire      [7:0] n19623;
wire            n19624;
wire      [7:0] n19625;
wire            n19626;
wire      [7:0] n19627;
wire            n19628;
wire      [7:0] n19629;
wire      [7:0] n1963;
wire            n19630;
wire      [7:0] n19631;
wire            n19632;
wire      [7:0] n19633;
wire            n19634;
wire      [7:0] n19635;
wire            n19636;
wire      [7:0] n19637;
wire            n19638;
wire      [7:0] n19639;
wire            n1964;
wire            n19640;
wire      [7:0] n19641;
wire            n19642;
wire      [7:0] n19643;
wire            n19644;
wire      [7:0] n19645;
wire            n19646;
wire      [7:0] n19647;
wire            n19648;
wire      [7:0] n19649;
wire      [7:0] n1965;
wire            n19650;
wire      [7:0] n19651;
wire            n19652;
wire      [7:0] n19653;
wire            n19654;
wire      [7:0] n19655;
wire            n19656;
wire      [7:0] n19657;
wire            n19658;
wire      [7:0] n19659;
wire            n1966;
wire            n19660;
wire      [7:0] n19661;
wire            n19662;
wire      [7:0] n19663;
wire            n19664;
wire      [7:0] n19665;
wire            n19666;
wire      [7:0] n19667;
wire            n19668;
wire      [7:0] n19669;
wire      [7:0] n1967;
wire            n19670;
wire      [7:0] n19671;
wire            n19672;
wire      [7:0] n19673;
wire            n19674;
wire      [7:0] n19675;
wire            n19676;
wire      [7:0] n19677;
wire            n19678;
wire      [7:0] n19679;
wire            n1968;
wire            n19680;
wire      [7:0] n19681;
wire            n19682;
wire      [7:0] n19683;
wire            n19684;
wire      [7:0] n19685;
wire            n19686;
wire      [7:0] n19687;
wire            n19688;
wire      [7:0] n19689;
wire      [7:0] n1969;
wire            n19690;
wire      [7:0] n19691;
wire            n19692;
wire      [7:0] n19693;
wire            n19694;
wire      [7:0] n19695;
wire            n19696;
wire      [7:0] n19697;
wire            n19698;
wire      [7:0] n19699;
wire            n197;
wire            n1970;
wire            n19700;
wire      [7:0] n19701;
wire            n19702;
wire      [7:0] n19703;
wire            n19704;
wire      [7:0] n19705;
wire            n19706;
wire      [7:0] n19707;
wire            n19708;
wire      [7:0] n19709;
wire      [7:0] n1971;
wire            n19710;
wire      [7:0] n19711;
wire            n19712;
wire      [7:0] n19713;
wire            n19714;
wire      [7:0] n19715;
wire            n19716;
wire      [7:0] n19717;
wire            n19718;
wire      [7:0] n19719;
wire            n1972;
wire            n19720;
wire      [7:0] n19721;
wire            n19722;
wire      [7:0] n19723;
wire            n19724;
wire      [7:0] n19725;
wire            n19726;
wire      [7:0] n19727;
wire            n19728;
wire      [7:0] n19729;
wire      [7:0] n1973;
wire            n19730;
wire      [7:0] n19731;
wire            n19732;
wire      [7:0] n19733;
wire            n19734;
wire      [7:0] n19735;
wire            n19736;
wire      [7:0] n19737;
wire            n19738;
wire      [7:0] n19739;
wire            n1974;
wire            n19740;
wire      [7:0] n19741;
wire            n19742;
wire      [7:0] n19743;
wire            n19744;
wire      [7:0] n19745;
wire            n19746;
wire      [7:0] n19747;
wire            n19748;
wire      [7:0] n19749;
wire      [7:0] n1975;
wire            n19750;
wire      [7:0] n19751;
wire            n19752;
wire      [7:0] n19753;
wire            n19754;
wire      [7:0] n19755;
wire            n19756;
wire      [7:0] n19757;
wire            n19758;
wire      [7:0] n19759;
wire            n1976;
wire            n19760;
wire      [7:0] n19761;
wire            n19762;
wire      [7:0] n19763;
wire            n19764;
wire      [7:0] n19765;
wire            n19766;
wire      [7:0] n19767;
wire            n19768;
wire      [7:0] n19769;
wire      [7:0] n1977;
wire            n19770;
wire      [7:0] n19771;
wire            n19772;
wire      [7:0] n19773;
wire            n19774;
wire      [7:0] n19775;
wire            n19776;
wire      [7:0] n19777;
wire            n19778;
wire      [7:0] n19779;
wire            n1978;
wire            n19780;
wire      [7:0] n19781;
wire            n19782;
wire      [7:0] n19783;
wire            n19784;
wire      [7:0] n19785;
wire            n19786;
wire      [7:0] n19787;
wire            n19788;
wire      [7:0] n19789;
wire      [7:0] n1979;
wire            n19790;
wire      [7:0] n19791;
wire            n19792;
wire      [7:0] n19793;
wire            n19794;
wire      [7:0] n19795;
wire            n19796;
wire      [7:0] n19797;
wire            n19798;
wire      [7:0] n19799;
wire            n1980;
wire            n19800;
wire      [7:0] n19801;
wire            n19802;
wire      [7:0] n19803;
wire            n19804;
wire      [7:0] n19805;
wire            n19806;
wire      [7:0] n19807;
wire            n19808;
wire      [7:0] n19809;
wire      [7:0] n1981;
wire            n19810;
wire      [7:0] n19811;
wire            n19812;
wire      [7:0] n19813;
wire            n19814;
wire      [7:0] n19815;
wire            n19816;
wire      [7:0] n19817;
wire            n19818;
wire      [7:0] n19819;
wire            n1982;
wire            n19820;
wire      [7:0] n19821;
wire            n19822;
wire      [7:0] n19823;
wire            n19824;
wire      [7:0] n19825;
wire            n19826;
wire      [7:0] n19827;
wire            n19828;
wire      [7:0] n19829;
wire      [7:0] n1983;
wire            n19830;
wire      [7:0] n19831;
wire            n19832;
wire      [7:0] n19833;
wire            n19834;
wire      [7:0] n19835;
wire            n19836;
wire      [7:0] n19837;
wire            n19838;
wire      [7:0] n19839;
wire            n1984;
wire            n19840;
wire      [7:0] n19841;
wire            n19842;
wire      [7:0] n19843;
wire            n19844;
wire      [7:0] n19845;
wire            n19846;
wire      [7:0] n19847;
wire            n19848;
wire      [7:0] n19849;
wire      [7:0] n1985;
wire            n19850;
wire      [7:0] n19851;
wire            n19852;
wire      [7:0] n19853;
wire            n19854;
wire      [7:0] n19855;
wire            n19856;
wire      [7:0] n19857;
wire            n19858;
wire      [7:0] n19859;
wire            n1986;
wire            n19860;
wire      [7:0] n19861;
wire            n19862;
wire      [7:0] n19863;
wire            n19864;
wire      [7:0] n19865;
wire            n19866;
wire      [7:0] n19867;
wire            n19868;
wire      [7:0] n19869;
wire      [7:0] n1987;
wire            n19870;
wire      [7:0] n19871;
wire            n19872;
wire      [7:0] n19873;
wire            n19874;
wire      [7:0] n19875;
wire            n19876;
wire      [7:0] n19877;
wire            n19878;
wire      [7:0] n19879;
wire            n1988;
wire            n19880;
wire      [7:0] n19881;
wire            n19882;
wire      [7:0] n19883;
wire            n19884;
wire      [7:0] n19885;
wire            n19886;
wire      [7:0] n19887;
wire            n19888;
wire      [7:0] n19889;
wire      [7:0] n1989;
wire            n19890;
wire      [7:0] n19891;
wire            n19892;
wire      [7:0] n19893;
wire            n19894;
wire      [7:0] n19895;
wire            n19896;
wire      [7:0] n19897;
wire            n19898;
wire      [7:0] n19899;
wire      [7:0] n199;
wire            n1990;
wire            n19900;
wire      [7:0] n19901;
wire            n19902;
wire      [7:0] n19903;
wire            n19904;
wire      [7:0] n19905;
wire            n19906;
wire      [7:0] n19907;
wire            n19908;
wire      [7:0] n19909;
wire      [7:0] n1991;
wire            n19910;
wire      [7:0] n19911;
wire            n19912;
wire      [7:0] n19913;
wire            n19914;
wire      [7:0] n19915;
wire            n19916;
wire      [7:0] n19917;
wire            n19918;
wire      [7:0] n19919;
wire            n1992;
wire            n19920;
wire      [7:0] n19921;
wire            n19922;
wire      [7:0] n19923;
wire            n19924;
wire      [7:0] n19925;
wire            n19926;
wire      [7:0] n19927;
wire            n19928;
wire      [7:0] n19929;
wire      [7:0] n1993;
wire            n19930;
wire      [7:0] n19931;
wire            n19932;
wire      [7:0] n19933;
wire            n19934;
wire      [7:0] n19935;
wire            n19936;
wire      [7:0] n19937;
wire            n19938;
wire      [7:0] n19939;
wire            n1994;
wire            n19940;
wire      [7:0] n19941;
wire            n19942;
wire      [7:0] n19943;
wire            n19944;
wire      [7:0] n19945;
wire            n19946;
wire      [7:0] n19947;
wire            n19948;
wire      [7:0] n19949;
wire      [7:0] n1995;
wire            n19950;
wire      [7:0] n19951;
wire            n19952;
wire      [7:0] n19953;
wire            n19954;
wire      [7:0] n19955;
wire            n19956;
wire      [7:0] n19957;
wire            n19958;
wire      [7:0] n19959;
wire            n1996;
wire            n19960;
wire      [7:0] n19961;
wire            n19962;
wire      [7:0] n19963;
wire            n19964;
wire      [7:0] n19965;
wire            n19966;
wire      [7:0] n19967;
wire            n19968;
wire      [7:0] n19969;
wire      [7:0] n1997;
wire            n19970;
wire      [7:0] n19971;
wire            n19972;
wire      [7:0] n19973;
wire            n19974;
wire      [7:0] n19975;
wire            n19976;
wire      [7:0] n19977;
wire            n19978;
wire      [7:0] n19979;
wire            n1998;
wire            n19980;
wire      [7:0] n19981;
wire            n19982;
wire      [7:0] n19983;
wire            n19984;
wire      [7:0] n19985;
wire            n19986;
wire      [7:0] n19987;
wire            n19988;
wire      [7:0] n19989;
wire      [7:0] n1999;
wire            n19990;
wire      [7:0] n19991;
wire            n19992;
wire      [7:0] n19993;
wire            n19994;
wire      [7:0] n19995;
wire            n19996;
wire      [7:0] n19997;
wire            n19998;
wire      [7:0] n19999;
wire      [7:0] n2;
wire            n20;
wire            n200;
wire            n2000;
wire            n20000;
wire      [7:0] n20001;
wire            n20002;
wire      [7:0] n20003;
wire            n20004;
wire      [7:0] n20005;
wire            n20006;
wire      [7:0] n20007;
wire            n20008;
wire      [7:0] n20009;
wire      [7:0] n2001;
wire            n20010;
wire      [7:0] n20011;
wire            n20012;
wire      [7:0] n20013;
wire            n20014;
wire      [7:0] n20015;
wire            n20016;
wire      [7:0] n20017;
wire            n20018;
wire      [7:0] n20019;
wire            n2002;
wire            n20020;
wire      [7:0] n20021;
wire            n20022;
wire      [7:0] n20023;
wire            n20024;
wire      [7:0] n20025;
wire            n20026;
wire      [7:0] n20027;
wire            n20028;
wire      [7:0] n20029;
wire      [7:0] n2003;
wire            n20030;
wire      [7:0] n20031;
wire            n20032;
wire      [7:0] n20033;
wire            n20034;
wire      [7:0] n20035;
wire            n20036;
wire      [7:0] n20037;
wire            n20038;
wire      [7:0] n20039;
wire            n2004;
wire            n20040;
wire      [7:0] n20041;
wire            n20042;
wire      [7:0] n20043;
wire            n20044;
wire      [7:0] n20045;
wire            n20046;
wire      [7:0] n20047;
wire            n20048;
wire      [7:0] n20049;
wire      [7:0] n2005;
wire            n20050;
wire      [7:0] n20051;
wire            n20052;
wire      [7:0] n20053;
wire      [7:0] n20054;
wire      [7:0] n20055;
wire      [7:0] n20056;
wire      [7:0] n20057;
wire      [7:0] n20058;
wire      [7:0] n20059;
wire            n2006;
wire      [7:0] n20060;
wire      [7:0] n20061;
wire      [7:0] n20062;
wire      [7:0] n20063;
wire      [7:0] n20064;
wire      [7:0] n20065;
wire      [7:0] n20066;
wire      [7:0] n20067;
wire      [7:0] n20068;
wire      [7:0] n20069;
wire      [7:0] n2007;
wire      [7:0] n20070;
wire      [7:0] n20071;
wire      [7:0] n20072;
wire      [7:0] n20073;
wire      [7:0] n20074;
wire      [7:0] n20075;
wire      [7:0] n20076;
wire      [7:0] n20077;
wire      [7:0] n20078;
wire      [7:0] n20079;
wire            n2008;
wire      [7:0] n20080;
wire      [7:0] n20081;
wire      [7:0] n20082;
wire      [7:0] n20083;
wire      [7:0] n20084;
wire      [7:0] n20085;
wire      [7:0] n20086;
wire      [7:0] n20087;
wire      [7:0] n20088;
wire      [7:0] n20089;
wire      [7:0] n2009;
wire      [7:0] n20090;
wire      [7:0] n20091;
wire      [7:0] n20092;
wire      [7:0] n20093;
wire      [7:0] n20094;
wire      [7:0] n20095;
wire      [7:0] n20096;
wire      [7:0] n20097;
wire      [7:0] n20098;
wire      [7:0] n20099;
wire            n2010;
wire      [7:0] n20100;
wire      [7:0] n20101;
wire      [7:0] n20102;
wire      [7:0] n20103;
wire      [7:0] n20104;
wire      [7:0] n20105;
wire      [7:0] n20106;
wire      [7:0] n20107;
wire      [7:0] n20108;
wire      [7:0] n20109;
wire      [7:0] n2011;
wire      [7:0] n20110;
wire      [7:0] n20111;
wire      [7:0] n20112;
wire      [7:0] n20113;
wire      [7:0] n20114;
wire      [7:0] n20115;
wire      [7:0] n20116;
wire      [7:0] n20117;
wire      [7:0] n20118;
wire      [7:0] n20119;
wire            n2012;
wire      [7:0] n20120;
wire      [7:0] n20121;
wire      [7:0] n20122;
wire      [7:0] n20123;
wire      [7:0] n20124;
wire      [7:0] n20125;
wire      [7:0] n20126;
wire      [7:0] n20127;
wire      [7:0] n20128;
wire      [7:0] n20129;
wire      [7:0] n2013;
wire      [7:0] n20130;
wire      [7:0] n20131;
wire      [7:0] n20132;
wire      [7:0] n20133;
wire      [7:0] n20134;
wire      [7:0] n20135;
wire      [7:0] n20136;
wire      [7:0] n20137;
wire      [7:0] n20138;
wire      [7:0] n20139;
wire            n2014;
wire      [7:0] n20140;
wire      [7:0] n20141;
wire      [7:0] n20142;
wire      [7:0] n20143;
wire      [7:0] n20144;
wire      [7:0] n20145;
wire      [7:0] n20146;
wire      [7:0] n20147;
wire      [7:0] n20148;
wire      [7:0] n20149;
wire      [7:0] n2015;
wire      [7:0] n20150;
wire      [7:0] n20151;
wire      [7:0] n20152;
wire      [7:0] n20153;
wire      [7:0] n20154;
wire      [7:0] n20155;
wire      [7:0] n20156;
wire      [7:0] n20157;
wire      [7:0] n20158;
wire      [7:0] n20159;
wire            n2016;
wire      [7:0] n20160;
wire      [7:0] n20161;
wire      [7:0] n20162;
wire      [7:0] n20163;
wire      [7:0] n20164;
wire      [7:0] n20165;
wire      [7:0] n20166;
wire      [7:0] n20167;
wire      [7:0] n20168;
wire      [7:0] n20169;
wire      [7:0] n2017;
wire      [7:0] n20170;
wire      [7:0] n20171;
wire      [7:0] n20172;
wire      [7:0] n20173;
wire      [7:0] n20174;
wire      [7:0] n20175;
wire      [7:0] n20176;
wire      [7:0] n20177;
wire      [7:0] n20178;
wire      [7:0] n20179;
wire            n2018;
wire      [7:0] n20180;
wire      [7:0] n20181;
wire      [7:0] n20182;
wire      [7:0] n20183;
wire      [7:0] n20184;
wire      [7:0] n20185;
wire      [7:0] n20186;
wire      [7:0] n20187;
wire      [7:0] n20188;
wire      [7:0] n20189;
wire      [7:0] n2019;
wire      [7:0] n20190;
wire      [7:0] n20191;
wire      [7:0] n20192;
wire      [7:0] n20193;
wire      [7:0] n20194;
wire      [7:0] n20195;
wire      [7:0] n20196;
wire      [7:0] n20197;
wire      [7:0] n20198;
wire      [7:0] n20199;
wire      [7:0] n202;
wire            n2020;
wire      [7:0] n20200;
wire      [7:0] n20201;
wire      [7:0] n20202;
wire      [7:0] n20203;
wire      [7:0] n20204;
wire      [7:0] n20205;
wire      [7:0] n20206;
wire      [7:0] n20207;
wire      [7:0] n20208;
wire      [7:0] n20209;
wire      [7:0] n2021;
wire      [7:0] n20210;
wire      [7:0] n20211;
wire      [7:0] n20212;
wire      [7:0] n20213;
wire      [7:0] n20214;
wire      [7:0] n20215;
wire      [7:0] n20216;
wire      [7:0] n20217;
wire      [7:0] n20218;
wire      [7:0] n20219;
wire            n2022;
wire      [7:0] n20220;
wire      [7:0] n20221;
wire      [7:0] n20222;
wire      [7:0] n20223;
wire      [7:0] n20224;
wire      [7:0] n20225;
wire      [7:0] n20226;
wire      [7:0] n20227;
wire      [7:0] n20228;
wire      [7:0] n20229;
wire      [7:0] n2023;
wire      [7:0] n20230;
wire      [7:0] n20231;
wire      [7:0] n20232;
wire      [7:0] n20233;
wire      [7:0] n20234;
wire      [7:0] n20235;
wire      [7:0] n20236;
wire      [7:0] n20237;
wire      [7:0] n20238;
wire      [7:0] n20239;
wire            n2024;
wire      [7:0] n20240;
wire      [7:0] n20241;
wire      [7:0] n20242;
wire      [7:0] n20243;
wire      [7:0] n20244;
wire      [7:0] n20245;
wire      [7:0] n20246;
wire      [7:0] n20247;
wire      [7:0] n20248;
wire      [7:0] n20249;
wire      [7:0] n2025;
wire      [7:0] n20250;
wire      [7:0] n20251;
wire      [7:0] n20252;
wire      [7:0] n20253;
wire      [7:0] n20254;
wire      [7:0] n20255;
wire      [7:0] n20256;
wire      [7:0] n20257;
wire      [7:0] n20258;
wire      [7:0] n20259;
wire            n2026;
wire      [7:0] n20260;
wire      [7:0] n20261;
wire      [7:0] n20262;
wire      [7:0] n20263;
wire      [7:0] n20264;
wire      [7:0] n20265;
wire      [7:0] n20266;
wire      [7:0] n20267;
wire      [7:0] n20268;
wire      [7:0] n20269;
wire      [7:0] n2027;
wire      [7:0] n20270;
wire      [7:0] n20271;
wire      [7:0] n20272;
wire      [7:0] n20273;
wire      [7:0] n20274;
wire      [7:0] n20275;
wire      [7:0] n20276;
wire      [7:0] n20277;
wire      [7:0] n20278;
wire      [7:0] n20279;
wire            n2028;
wire      [7:0] n20280;
wire      [7:0] n20281;
wire      [7:0] n20282;
wire      [7:0] n20283;
wire      [7:0] n20284;
wire      [7:0] n20285;
wire      [7:0] n20286;
wire      [7:0] n20287;
wire      [7:0] n20288;
wire      [7:0] n20289;
wire      [7:0] n2029;
wire      [7:0] n20290;
wire      [7:0] n20291;
wire      [7:0] n20292;
wire      [7:0] n20293;
wire      [7:0] n20294;
wire      [7:0] n20295;
wire      [7:0] n20296;
wire      [7:0] n20297;
wire      [7:0] n20298;
wire      [7:0] n20299;
wire            n2030;
wire      [7:0] n20300;
wire      [7:0] n20301;
wire      [7:0] n20302;
wire      [7:0] n20303;
wire      [7:0] n20304;
wire      [7:0] n20305;
wire      [7:0] n20306;
wire      [7:0] n20307;
wire      [7:0] n20308;
wire      [7:0] n20309;
wire      [7:0] n2031;
wire      [7:0] n20310;
wire            n20311;
wire      [7:0] n20312;
wire            n20313;
wire      [7:0] n20314;
wire            n20315;
wire      [7:0] n20316;
wire            n20317;
wire      [7:0] n20318;
wire            n20319;
wire            n2032;
wire      [7:0] n20320;
wire            n20321;
wire      [7:0] n20322;
wire            n20323;
wire      [7:0] n20324;
wire            n20325;
wire      [7:0] n20326;
wire            n20327;
wire      [7:0] n20328;
wire            n20329;
wire      [7:0] n2033;
wire      [7:0] n20330;
wire            n20331;
wire      [7:0] n20332;
wire            n20333;
wire      [7:0] n20334;
wire            n20335;
wire      [7:0] n20336;
wire            n20337;
wire      [7:0] n20338;
wire            n20339;
wire            n2034;
wire      [7:0] n20340;
wire            n20341;
wire      [7:0] n20342;
wire            n20343;
wire      [7:0] n20344;
wire            n20345;
wire      [7:0] n20346;
wire            n20347;
wire      [7:0] n20348;
wire            n20349;
wire      [7:0] n2035;
wire      [7:0] n20350;
wire            n20351;
wire      [7:0] n20352;
wire            n20353;
wire      [7:0] n20354;
wire            n20355;
wire      [7:0] n20356;
wire            n20357;
wire      [7:0] n20358;
wire            n20359;
wire            n2036;
wire      [7:0] n20360;
wire            n20361;
wire      [7:0] n20362;
wire            n20363;
wire      [7:0] n20364;
wire            n20365;
wire      [7:0] n20366;
wire            n20367;
wire      [7:0] n20368;
wire            n20369;
wire      [7:0] n2037;
wire      [7:0] n20370;
wire            n20371;
wire      [7:0] n20372;
wire            n20373;
wire      [7:0] n20374;
wire            n20375;
wire      [7:0] n20376;
wire            n20377;
wire      [7:0] n20378;
wire            n20379;
wire            n2038;
wire      [7:0] n20380;
wire            n20381;
wire      [7:0] n20382;
wire            n20383;
wire      [7:0] n20384;
wire            n20385;
wire      [7:0] n20386;
wire            n20387;
wire      [7:0] n20388;
wire            n20389;
wire      [7:0] n2039;
wire      [7:0] n20390;
wire            n20391;
wire      [7:0] n20392;
wire            n20393;
wire      [7:0] n20394;
wire            n20395;
wire      [7:0] n20396;
wire            n20397;
wire      [7:0] n20398;
wire            n20399;
wire            n204;
wire            n2040;
wire      [7:0] n20400;
wire            n20401;
wire      [7:0] n20402;
wire            n20403;
wire      [7:0] n20404;
wire            n20405;
wire      [7:0] n20406;
wire            n20407;
wire      [7:0] n20408;
wire            n20409;
wire      [7:0] n2041;
wire      [7:0] n20410;
wire            n20411;
wire      [7:0] n20412;
wire            n20413;
wire      [7:0] n20414;
wire            n20415;
wire      [7:0] n20416;
wire            n20417;
wire      [7:0] n20418;
wire            n20419;
wire            n2042;
wire      [7:0] n20420;
wire            n20421;
wire      [7:0] n20422;
wire            n20423;
wire      [7:0] n20424;
wire            n20425;
wire      [7:0] n20426;
wire            n20427;
wire      [7:0] n20428;
wire            n20429;
wire      [7:0] n2043;
wire      [7:0] n20430;
wire            n20431;
wire      [7:0] n20432;
wire            n20433;
wire      [7:0] n20434;
wire            n20435;
wire      [7:0] n20436;
wire            n20437;
wire      [7:0] n20438;
wire            n20439;
wire            n2044;
wire      [7:0] n20440;
wire            n20441;
wire      [7:0] n20442;
wire            n20443;
wire      [7:0] n20444;
wire            n20445;
wire      [7:0] n20446;
wire            n20447;
wire      [7:0] n20448;
wire            n20449;
wire      [7:0] n2045;
wire      [7:0] n20450;
wire            n20451;
wire      [7:0] n20452;
wire            n20453;
wire      [7:0] n20454;
wire            n20455;
wire      [7:0] n20456;
wire            n20457;
wire      [7:0] n20458;
wire            n20459;
wire            n2046;
wire      [7:0] n20460;
wire            n20461;
wire      [7:0] n20462;
wire            n20463;
wire      [7:0] n20464;
wire            n20465;
wire      [7:0] n20466;
wire            n20467;
wire      [7:0] n20468;
wire            n20469;
wire      [7:0] n2047;
wire      [7:0] n20470;
wire            n20471;
wire      [7:0] n20472;
wire            n20473;
wire      [7:0] n20474;
wire            n20475;
wire      [7:0] n20476;
wire            n20477;
wire      [7:0] n20478;
wire            n20479;
wire            n2048;
wire      [7:0] n20480;
wire            n20481;
wire      [7:0] n20482;
wire            n20483;
wire      [7:0] n20484;
wire            n20485;
wire      [7:0] n20486;
wire            n20487;
wire      [7:0] n20488;
wire            n20489;
wire      [7:0] n2049;
wire      [7:0] n20490;
wire            n20491;
wire      [7:0] n20492;
wire            n20493;
wire      [7:0] n20494;
wire            n20495;
wire      [7:0] n20496;
wire            n20497;
wire      [7:0] n20498;
wire            n20499;
wire            n2050;
wire      [7:0] n20500;
wire            n20501;
wire      [7:0] n20502;
wire            n20503;
wire      [7:0] n20504;
wire            n20505;
wire      [7:0] n20506;
wire            n20507;
wire      [7:0] n20508;
wire            n20509;
wire      [7:0] n2051;
wire      [7:0] n20510;
wire            n20511;
wire      [7:0] n20512;
wire            n20513;
wire      [7:0] n20514;
wire            n20515;
wire      [7:0] n20516;
wire            n20517;
wire      [7:0] n20518;
wire            n20519;
wire            n2052;
wire      [7:0] n20520;
wire            n20521;
wire      [7:0] n20522;
wire            n20523;
wire      [7:0] n20524;
wire            n20525;
wire      [7:0] n20526;
wire            n20527;
wire      [7:0] n20528;
wire            n20529;
wire      [7:0] n2053;
wire      [7:0] n20530;
wire            n20531;
wire      [7:0] n20532;
wire            n20533;
wire      [7:0] n20534;
wire            n20535;
wire      [7:0] n20536;
wire            n20537;
wire      [7:0] n20538;
wire            n20539;
wire            n2054;
wire      [7:0] n20540;
wire            n20541;
wire      [7:0] n20542;
wire            n20543;
wire      [7:0] n20544;
wire            n20545;
wire      [7:0] n20546;
wire            n20547;
wire      [7:0] n20548;
wire            n20549;
wire      [7:0] n2055;
wire      [7:0] n20550;
wire            n20551;
wire      [7:0] n20552;
wire            n20553;
wire      [7:0] n20554;
wire            n20555;
wire      [7:0] n20556;
wire            n20557;
wire      [7:0] n20558;
wire            n20559;
wire            n2056;
wire      [7:0] n20560;
wire            n20561;
wire      [7:0] n20562;
wire            n20563;
wire      [7:0] n20564;
wire            n20565;
wire      [7:0] n20566;
wire            n20567;
wire      [7:0] n20568;
wire            n20569;
wire      [7:0] n2057;
wire      [7:0] n20570;
wire            n20571;
wire      [7:0] n20572;
wire            n20573;
wire      [7:0] n20574;
wire            n20575;
wire      [7:0] n20576;
wire            n20577;
wire      [7:0] n20578;
wire            n20579;
wire            n2058;
wire      [7:0] n20580;
wire            n20581;
wire      [7:0] n20582;
wire            n20583;
wire      [7:0] n20584;
wire            n20585;
wire      [7:0] n20586;
wire            n20587;
wire      [7:0] n20588;
wire            n20589;
wire      [7:0] n2059;
wire      [7:0] n20590;
wire            n20591;
wire      [7:0] n20592;
wire            n20593;
wire      [7:0] n20594;
wire            n20595;
wire      [7:0] n20596;
wire            n20597;
wire      [7:0] n20598;
wire            n20599;
wire      [7:0] n206;
wire            n2060;
wire      [7:0] n20600;
wire            n20601;
wire      [7:0] n20602;
wire            n20603;
wire      [7:0] n20604;
wire            n20605;
wire      [7:0] n20606;
wire            n20607;
wire      [7:0] n20608;
wire            n20609;
wire      [7:0] n2061;
wire      [7:0] n20610;
wire            n20611;
wire      [7:0] n20612;
wire            n20613;
wire      [7:0] n20614;
wire            n20615;
wire      [7:0] n20616;
wire            n20617;
wire      [7:0] n20618;
wire            n20619;
wire            n2062;
wire      [7:0] n20620;
wire            n20621;
wire      [7:0] n20622;
wire            n20623;
wire      [7:0] n20624;
wire            n20625;
wire      [7:0] n20626;
wire            n20627;
wire      [7:0] n20628;
wire            n20629;
wire      [7:0] n2063;
wire      [7:0] n20630;
wire            n20631;
wire      [7:0] n20632;
wire            n20633;
wire      [7:0] n20634;
wire            n20635;
wire      [7:0] n20636;
wire            n20637;
wire      [7:0] n20638;
wire            n20639;
wire            n2064;
wire      [7:0] n20640;
wire            n20641;
wire      [7:0] n20642;
wire            n20643;
wire      [7:0] n20644;
wire            n20645;
wire      [7:0] n20646;
wire            n20647;
wire      [7:0] n20648;
wire            n20649;
wire      [7:0] n2065;
wire      [7:0] n20650;
wire            n20651;
wire      [7:0] n20652;
wire            n20653;
wire      [7:0] n20654;
wire            n20655;
wire      [7:0] n20656;
wire            n20657;
wire      [7:0] n20658;
wire            n20659;
wire            n2066;
wire      [7:0] n20660;
wire            n20661;
wire      [7:0] n20662;
wire            n20663;
wire      [7:0] n20664;
wire            n20665;
wire      [7:0] n20666;
wire            n20667;
wire      [7:0] n20668;
wire            n20669;
wire      [7:0] n2067;
wire      [7:0] n20670;
wire            n20671;
wire      [7:0] n20672;
wire            n20673;
wire      [7:0] n20674;
wire            n20675;
wire      [7:0] n20676;
wire            n20677;
wire      [7:0] n20678;
wire            n20679;
wire            n2068;
wire      [7:0] n20680;
wire            n20681;
wire      [7:0] n20682;
wire            n20683;
wire      [7:0] n20684;
wire            n20685;
wire      [7:0] n20686;
wire            n20687;
wire      [7:0] n20688;
wire            n20689;
wire      [7:0] n2069;
wire      [7:0] n20690;
wire            n20691;
wire      [7:0] n20692;
wire            n20693;
wire      [7:0] n20694;
wire            n20695;
wire      [7:0] n20696;
wire            n20697;
wire      [7:0] n20698;
wire            n20699;
wire            n2070;
wire      [7:0] n20700;
wire            n20701;
wire      [7:0] n20702;
wire            n20703;
wire      [7:0] n20704;
wire            n20705;
wire      [7:0] n20706;
wire            n20707;
wire      [7:0] n20708;
wire            n20709;
wire      [7:0] n2071;
wire      [7:0] n20710;
wire            n20711;
wire      [7:0] n20712;
wire            n20713;
wire      [7:0] n20714;
wire            n20715;
wire      [7:0] n20716;
wire            n20717;
wire      [7:0] n20718;
wire            n20719;
wire            n2072;
wire      [7:0] n20720;
wire            n20721;
wire      [7:0] n20722;
wire            n20723;
wire      [7:0] n20724;
wire            n20725;
wire      [7:0] n20726;
wire            n20727;
wire      [7:0] n20728;
wire            n20729;
wire      [7:0] n2073;
wire      [7:0] n20730;
wire            n20731;
wire      [7:0] n20732;
wire            n20733;
wire      [7:0] n20734;
wire            n20735;
wire      [7:0] n20736;
wire            n20737;
wire      [7:0] n20738;
wire            n20739;
wire            n2074;
wire      [7:0] n20740;
wire            n20741;
wire      [7:0] n20742;
wire            n20743;
wire      [7:0] n20744;
wire            n20745;
wire      [7:0] n20746;
wire            n20747;
wire      [7:0] n20748;
wire            n20749;
wire      [7:0] n2075;
wire      [7:0] n20750;
wire            n20751;
wire      [7:0] n20752;
wire            n20753;
wire      [7:0] n20754;
wire            n20755;
wire      [7:0] n20756;
wire            n20757;
wire      [7:0] n20758;
wire            n20759;
wire            n2076;
wire      [7:0] n20760;
wire            n20761;
wire      [7:0] n20762;
wire            n20763;
wire      [7:0] n20764;
wire            n20765;
wire      [7:0] n20766;
wire            n20767;
wire      [7:0] n20768;
wire            n20769;
wire      [7:0] n2077;
wire      [7:0] n20770;
wire            n20771;
wire      [7:0] n20772;
wire            n20773;
wire      [7:0] n20774;
wire            n20775;
wire      [7:0] n20776;
wire            n20777;
wire      [7:0] n20778;
wire            n20779;
wire            n2078;
wire      [7:0] n20780;
wire            n20781;
wire      [7:0] n20782;
wire            n20783;
wire      [7:0] n20784;
wire            n20785;
wire      [7:0] n20786;
wire            n20787;
wire      [7:0] n20788;
wire            n20789;
wire      [7:0] n2079;
wire      [7:0] n20790;
wire            n20791;
wire      [7:0] n20792;
wire            n20793;
wire      [7:0] n20794;
wire            n20795;
wire      [7:0] n20796;
wire            n20797;
wire      [7:0] n20798;
wire            n20799;
wire            n208;
wire            n2080;
wire      [7:0] n20800;
wire            n20801;
wire      [7:0] n20802;
wire            n20803;
wire      [7:0] n20804;
wire            n20805;
wire      [7:0] n20806;
wire            n20807;
wire      [7:0] n20808;
wire            n20809;
wire      [7:0] n2081;
wire      [7:0] n20810;
wire            n20811;
wire      [7:0] n20812;
wire            n20813;
wire      [7:0] n20814;
wire            n20815;
wire      [7:0] n20816;
wire            n20817;
wire      [7:0] n20818;
wire            n20819;
wire            n2082;
wire      [7:0] n20820;
wire            n20821;
wire      [7:0] n20822;
wire      [7:0] n20823;
wire      [7:0] n20824;
wire      [7:0] n20825;
wire      [7:0] n20826;
wire      [7:0] n20827;
wire      [7:0] n20828;
wire      [7:0] n20829;
wire      [7:0] n2083;
wire      [7:0] n20830;
wire      [7:0] n20831;
wire      [7:0] n20832;
wire      [7:0] n20833;
wire      [7:0] n20834;
wire      [7:0] n20835;
wire      [7:0] n20836;
wire      [7:0] n20837;
wire      [7:0] n20838;
wire      [7:0] n20839;
wire            n2084;
wire      [7:0] n20840;
wire      [7:0] n20841;
wire      [7:0] n20842;
wire      [7:0] n20843;
wire      [7:0] n20844;
wire      [7:0] n20845;
wire      [7:0] n20846;
wire      [7:0] n20847;
wire      [7:0] n20848;
wire      [7:0] n20849;
wire      [7:0] n2085;
wire      [7:0] n20850;
wire      [7:0] n20851;
wire      [7:0] n20852;
wire      [7:0] n20853;
wire      [7:0] n20854;
wire      [7:0] n20855;
wire      [7:0] n20856;
wire      [7:0] n20857;
wire      [7:0] n20858;
wire      [7:0] n20859;
wire            n2086;
wire      [7:0] n20860;
wire      [7:0] n20861;
wire      [7:0] n20862;
wire      [7:0] n20863;
wire      [7:0] n20864;
wire      [7:0] n20865;
wire      [7:0] n20866;
wire      [7:0] n20867;
wire      [7:0] n20868;
wire      [7:0] n20869;
wire      [7:0] n2087;
wire      [7:0] n20870;
wire      [7:0] n20871;
wire      [7:0] n20872;
wire      [7:0] n20873;
wire      [7:0] n20874;
wire      [7:0] n20875;
wire      [7:0] n20876;
wire      [7:0] n20877;
wire      [7:0] n20878;
wire      [7:0] n20879;
wire            n2088;
wire      [7:0] n20880;
wire      [7:0] n20881;
wire      [7:0] n20882;
wire      [7:0] n20883;
wire      [7:0] n20884;
wire      [7:0] n20885;
wire      [7:0] n20886;
wire      [7:0] n20887;
wire      [7:0] n20888;
wire      [7:0] n20889;
wire      [7:0] n2089;
wire      [7:0] n20890;
wire      [7:0] n20891;
wire      [7:0] n20892;
wire      [7:0] n20893;
wire      [7:0] n20894;
wire      [7:0] n20895;
wire      [7:0] n20896;
wire      [7:0] n20897;
wire      [7:0] n20898;
wire      [7:0] n20899;
wire      [7:0] n209;
wire            n2090;
wire      [7:0] n20900;
wire      [7:0] n20901;
wire      [7:0] n20902;
wire      [7:0] n20903;
wire      [7:0] n20904;
wire      [7:0] n20905;
wire      [7:0] n20906;
wire      [7:0] n20907;
wire      [7:0] n20908;
wire      [7:0] n20909;
wire      [7:0] n2091;
wire      [7:0] n20910;
wire      [7:0] n20911;
wire      [7:0] n20912;
wire      [7:0] n20913;
wire      [7:0] n20914;
wire      [7:0] n20915;
wire      [7:0] n20916;
wire      [7:0] n20917;
wire      [7:0] n20918;
wire      [7:0] n20919;
wire            n2092;
wire      [7:0] n20920;
wire      [7:0] n20921;
wire      [7:0] n20922;
wire      [7:0] n20923;
wire      [7:0] n20924;
wire      [7:0] n20925;
wire      [7:0] n20926;
wire      [7:0] n20927;
wire      [7:0] n20928;
wire      [7:0] n20929;
wire      [7:0] n2093;
wire      [7:0] n20930;
wire      [7:0] n20931;
wire      [7:0] n20932;
wire      [7:0] n20933;
wire      [7:0] n20934;
wire      [7:0] n20935;
wire      [7:0] n20936;
wire      [7:0] n20937;
wire      [7:0] n20938;
wire      [7:0] n20939;
wire            n2094;
wire      [7:0] n20940;
wire      [7:0] n20941;
wire      [7:0] n20942;
wire      [7:0] n20943;
wire      [7:0] n20944;
wire      [7:0] n20945;
wire      [7:0] n20946;
wire      [7:0] n20947;
wire      [7:0] n20948;
wire      [7:0] n20949;
wire      [7:0] n2095;
wire      [7:0] n20950;
wire      [7:0] n20951;
wire      [7:0] n20952;
wire      [7:0] n20953;
wire      [7:0] n20954;
wire      [7:0] n20955;
wire      [7:0] n20956;
wire      [7:0] n20957;
wire      [7:0] n20958;
wire      [7:0] n20959;
wire            n2096;
wire      [7:0] n20960;
wire      [7:0] n20961;
wire      [7:0] n20962;
wire      [7:0] n20963;
wire      [7:0] n20964;
wire      [7:0] n20965;
wire      [7:0] n20966;
wire      [7:0] n20967;
wire      [7:0] n20968;
wire      [7:0] n20969;
wire      [7:0] n2097;
wire      [7:0] n20970;
wire      [7:0] n20971;
wire      [7:0] n20972;
wire      [7:0] n20973;
wire      [7:0] n20974;
wire      [7:0] n20975;
wire      [7:0] n20976;
wire      [7:0] n20977;
wire      [7:0] n20978;
wire      [7:0] n20979;
wire            n2098;
wire      [7:0] n20980;
wire      [7:0] n20981;
wire      [7:0] n20982;
wire      [7:0] n20983;
wire      [7:0] n20984;
wire      [7:0] n20985;
wire      [7:0] n20986;
wire      [7:0] n20987;
wire      [7:0] n20988;
wire      [7:0] n20989;
wire      [7:0] n2099;
wire      [7:0] n20990;
wire      [7:0] n20991;
wire      [7:0] n20992;
wire      [7:0] n20993;
wire      [7:0] n20994;
wire      [7:0] n20995;
wire      [7:0] n20996;
wire      [7:0] n20997;
wire      [7:0] n20998;
wire      [7:0] n20999;
wire            n210;
wire            n2100;
wire      [7:0] n21000;
wire      [7:0] n21001;
wire      [7:0] n21002;
wire      [7:0] n21003;
wire      [7:0] n21004;
wire      [7:0] n21005;
wire      [7:0] n21006;
wire      [7:0] n21007;
wire      [7:0] n21008;
wire      [7:0] n21009;
wire      [7:0] n2101;
wire      [7:0] n21010;
wire      [7:0] n21011;
wire      [7:0] n21012;
wire      [7:0] n21013;
wire      [7:0] n21014;
wire      [7:0] n21015;
wire      [7:0] n21016;
wire      [7:0] n21017;
wire      [7:0] n21018;
wire      [7:0] n21019;
wire            n2102;
wire      [7:0] n21020;
wire      [7:0] n21021;
wire      [7:0] n21022;
wire      [7:0] n21023;
wire      [7:0] n21024;
wire      [7:0] n21025;
wire      [7:0] n21026;
wire      [7:0] n21027;
wire      [7:0] n21028;
wire      [7:0] n21029;
wire      [7:0] n2103;
wire      [7:0] n21030;
wire      [7:0] n21031;
wire      [7:0] n21032;
wire      [7:0] n21033;
wire      [7:0] n21034;
wire      [7:0] n21035;
wire      [7:0] n21036;
wire      [7:0] n21037;
wire      [7:0] n21038;
wire      [7:0] n21039;
wire            n2104;
wire      [7:0] n21040;
wire      [7:0] n21041;
wire      [7:0] n21042;
wire      [7:0] n21043;
wire      [7:0] n21044;
wire      [7:0] n21045;
wire      [7:0] n21046;
wire      [7:0] n21047;
wire      [7:0] n21048;
wire      [7:0] n21049;
wire      [7:0] n2105;
wire      [7:0] n21050;
wire      [7:0] n21051;
wire      [7:0] n21052;
wire      [7:0] n21053;
wire      [7:0] n21054;
wire      [7:0] n21055;
wire      [7:0] n21056;
wire      [7:0] n21057;
wire      [7:0] n21058;
wire      [7:0] n21059;
wire            n2106;
wire      [7:0] n21060;
wire      [7:0] n21061;
wire      [7:0] n21062;
wire      [7:0] n21063;
wire      [7:0] n21064;
wire      [7:0] n21065;
wire      [7:0] n21066;
wire      [7:0] n21067;
wire      [7:0] n21068;
wire      [7:0] n21069;
wire      [7:0] n2107;
wire      [7:0] n21070;
wire      [7:0] n21071;
wire      [7:0] n21072;
wire      [7:0] n21073;
wire      [7:0] n21074;
wire      [7:0] n21075;
wire      [7:0] n21076;
wire      [7:0] n21077;
wire      [7:0] n21078;
wire      [7:0] n21079;
wire            n2108;
wire            n21080;
wire      [7:0] n21081;
wire            n21082;
wire      [7:0] n21083;
wire            n21084;
wire      [7:0] n21085;
wire            n21086;
wire      [7:0] n21087;
wire            n21088;
wire      [7:0] n21089;
wire      [7:0] n2109;
wire            n21090;
wire      [7:0] n21091;
wire            n21092;
wire      [7:0] n21093;
wire            n21094;
wire      [7:0] n21095;
wire            n21096;
wire      [7:0] n21097;
wire            n21098;
wire      [7:0] n21099;
wire            n2110;
wire            n21100;
wire      [7:0] n21101;
wire            n21102;
wire      [7:0] n21103;
wire            n21104;
wire      [7:0] n21105;
wire            n21106;
wire      [7:0] n21107;
wire            n21108;
wire      [7:0] n21109;
wire      [7:0] n2111;
wire            n21110;
wire      [7:0] n21111;
wire            n21112;
wire      [7:0] n21113;
wire            n21114;
wire      [7:0] n21115;
wire            n21116;
wire      [7:0] n21117;
wire            n21118;
wire      [7:0] n21119;
wire            n2112;
wire            n21120;
wire      [7:0] n21121;
wire            n21122;
wire      [7:0] n21123;
wire            n21124;
wire      [7:0] n21125;
wire            n21126;
wire      [7:0] n21127;
wire            n21128;
wire      [7:0] n21129;
wire      [7:0] n2113;
wire            n21130;
wire      [7:0] n21131;
wire            n21132;
wire      [7:0] n21133;
wire            n21134;
wire      [7:0] n21135;
wire            n21136;
wire      [7:0] n21137;
wire            n21138;
wire      [7:0] n21139;
wire            n2114;
wire            n21140;
wire      [7:0] n21141;
wire            n21142;
wire      [7:0] n21143;
wire            n21144;
wire      [7:0] n21145;
wire            n21146;
wire      [7:0] n21147;
wire            n21148;
wire      [7:0] n21149;
wire      [7:0] n2115;
wire            n21150;
wire      [7:0] n21151;
wire            n21152;
wire      [7:0] n21153;
wire            n21154;
wire      [7:0] n21155;
wire            n21156;
wire      [7:0] n21157;
wire            n21158;
wire      [7:0] n21159;
wire            n2116;
wire            n21160;
wire      [7:0] n21161;
wire            n21162;
wire      [7:0] n21163;
wire            n21164;
wire      [7:0] n21165;
wire            n21166;
wire      [7:0] n21167;
wire            n21168;
wire      [7:0] n21169;
wire      [7:0] n2117;
wire            n21170;
wire      [7:0] n21171;
wire            n21172;
wire      [7:0] n21173;
wire            n21174;
wire      [7:0] n21175;
wire            n21176;
wire      [7:0] n21177;
wire            n21178;
wire      [7:0] n21179;
wire            n2118;
wire            n21180;
wire      [7:0] n21181;
wire            n21182;
wire      [7:0] n21183;
wire            n21184;
wire      [7:0] n21185;
wire            n21186;
wire      [7:0] n21187;
wire            n21188;
wire      [7:0] n21189;
wire      [7:0] n2119;
wire            n21190;
wire      [7:0] n21191;
wire            n21192;
wire      [7:0] n21193;
wire            n21194;
wire      [7:0] n21195;
wire            n21196;
wire      [7:0] n21197;
wire            n21198;
wire      [7:0] n21199;
wire      [7:0] n212;
wire            n2120;
wire            n21200;
wire      [7:0] n21201;
wire            n21202;
wire      [7:0] n21203;
wire            n21204;
wire      [7:0] n21205;
wire            n21206;
wire      [7:0] n21207;
wire            n21208;
wire      [7:0] n21209;
wire      [7:0] n2121;
wire            n21210;
wire      [7:0] n21211;
wire            n21212;
wire      [7:0] n21213;
wire            n21214;
wire      [7:0] n21215;
wire            n21216;
wire      [7:0] n21217;
wire            n21218;
wire      [7:0] n21219;
wire            n2122;
wire            n21220;
wire      [7:0] n21221;
wire            n21222;
wire      [7:0] n21223;
wire            n21224;
wire      [7:0] n21225;
wire            n21226;
wire      [7:0] n21227;
wire            n21228;
wire      [7:0] n21229;
wire      [7:0] n2123;
wire            n21230;
wire      [7:0] n21231;
wire            n21232;
wire      [7:0] n21233;
wire            n21234;
wire      [7:0] n21235;
wire            n21236;
wire      [7:0] n21237;
wire            n21238;
wire      [7:0] n21239;
wire            n2124;
wire            n21240;
wire      [7:0] n21241;
wire            n21242;
wire      [7:0] n21243;
wire            n21244;
wire      [7:0] n21245;
wire            n21246;
wire      [7:0] n21247;
wire            n21248;
wire      [7:0] n21249;
wire      [7:0] n2125;
wire            n21250;
wire      [7:0] n21251;
wire            n21252;
wire      [7:0] n21253;
wire            n21254;
wire      [7:0] n21255;
wire            n21256;
wire      [7:0] n21257;
wire            n21258;
wire      [7:0] n21259;
wire            n2126;
wire            n21260;
wire      [7:0] n21261;
wire            n21262;
wire      [7:0] n21263;
wire            n21264;
wire      [7:0] n21265;
wire            n21266;
wire      [7:0] n21267;
wire            n21268;
wire      [7:0] n21269;
wire      [7:0] n2127;
wire            n21270;
wire      [7:0] n21271;
wire            n21272;
wire      [7:0] n21273;
wire            n21274;
wire      [7:0] n21275;
wire            n21276;
wire      [7:0] n21277;
wire            n21278;
wire      [7:0] n21279;
wire            n2128;
wire            n21280;
wire      [7:0] n21281;
wire            n21282;
wire      [7:0] n21283;
wire            n21284;
wire      [7:0] n21285;
wire            n21286;
wire      [7:0] n21287;
wire            n21288;
wire      [7:0] n21289;
wire      [7:0] n2129;
wire            n21290;
wire      [7:0] n21291;
wire            n21292;
wire      [7:0] n21293;
wire            n21294;
wire      [7:0] n21295;
wire            n21296;
wire      [7:0] n21297;
wire            n21298;
wire      [7:0] n21299;
wire            n2130;
wire            n21300;
wire      [7:0] n21301;
wire            n21302;
wire      [7:0] n21303;
wire            n21304;
wire      [7:0] n21305;
wire            n21306;
wire      [7:0] n21307;
wire            n21308;
wire      [7:0] n21309;
wire      [7:0] n2131;
wire            n21310;
wire      [7:0] n21311;
wire            n21312;
wire      [7:0] n21313;
wire            n21314;
wire      [7:0] n21315;
wire            n21316;
wire      [7:0] n21317;
wire            n21318;
wire      [7:0] n21319;
wire            n2132;
wire            n21320;
wire      [7:0] n21321;
wire            n21322;
wire      [7:0] n21323;
wire            n21324;
wire      [7:0] n21325;
wire            n21326;
wire      [7:0] n21327;
wire            n21328;
wire      [7:0] n21329;
wire      [7:0] n2133;
wire            n21330;
wire      [7:0] n21331;
wire            n21332;
wire      [7:0] n21333;
wire            n21334;
wire      [7:0] n21335;
wire            n21336;
wire      [7:0] n21337;
wire            n21338;
wire      [7:0] n21339;
wire            n2134;
wire            n21340;
wire      [7:0] n21341;
wire            n21342;
wire      [7:0] n21343;
wire            n21344;
wire      [7:0] n21345;
wire            n21346;
wire      [7:0] n21347;
wire            n21348;
wire      [7:0] n21349;
wire      [7:0] n2135;
wire            n21350;
wire      [7:0] n21351;
wire            n21352;
wire      [7:0] n21353;
wire            n21354;
wire      [7:0] n21355;
wire            n21356;
wire      [7:0] n21357;
wire            n21358;
wire      [7:0] n21359;
wire            n2136;
wire            n21360;
wire      [7:0] n21361;
wire            n21362;
wire      [7:0] n21363;
wire            n21364;
wire      [7:0] n21365;
wire            n21366;
wire      [7:0] n21367;
wire            n21368;
wire      [7:0] n21369;
wire      [7:0] n2137;
wire            n21370;
wire      [7:0] n21371;
wire            n21372;
wire      [7:0] n21373;
wire            n21374;
wire      [7:0] n21375;
wire            n21376;
wire      [7:0] n21377;
wire            n21378;
wire      [7:0] n21379;
wire            n2138;
wire            n21380;
wire      [7:0] n21381;
wire            n21382;
wire      [7:0] n21383;
wire            n21384;
wire      [7:0] n21385;
wire            n21386;
wire      [7:0] n21387;
wire            n21388;
wire      [7:0] n21389;
wire      [7:0] n2139;
wire            n21390;
wire      [7:0] n21391;
wire            n21392;
wire      [7:0] n21393;
wire            n21394;
wire      [7:0] n21395;
wire            n21396;
wire      [7:0] n21397;
wire            n21398;
wire      [7:0] n21399;
wire            n214;
wire            n2140;
wire            n21400;
wire      [7:0] n21401;
wire            n21402;
wire      [7:0] n21403;
wire            n21404;
wire      [7:0] n21405;
wire            n21406;
wire      [7:0] n21407;
wire            n21408;
wire      [7:0] n21409;
wire      [7:0] n2141;
wire            n21410;
wire      [7:0] n21411;
wire            n21412;
wire      [7:0] n21413;
wire            n21414;
wire      [7:0] n21415;
wire            n21416;
wire      [7:0] n21417;
wire            n21418;
wire      [7:0] n21419;
wire            n2142;
wire            n21420;
wire      [7:0] n21421;
wire            n21422;
wire      [7:0] n21423;
wire            n21424;
wire      [7:0] n21425;
wire            n21426;
wire      [7:0] n21427;
wire            n21428;
wire      [7:0] n21429;
wire      [7:0] n2143;
wire            n21430;
wire      [7:0] n21431;
wire            n21432;
wire      [7:0] n21433;
wire            n21434;
wire      [7:0] n21435;
wire            n21436;
wire      [7:0] n21437;
wire            n21438;
wire      [7:0] n21439;
wire            n2144;
wire            n21440;
wire      [7:0] n21441;
wire            n21442;
wire      [7:0] n21443;
wire            n21444;
wire      [7:0] n21445;
wire            n21446;
wire      [7:0] n21447;
wire            n21448;
wire      [7:0] n21449;
wire      [7:0] n2145;
wire            n21450;
wire      [7:0] n21451;
wire            n21452;
wire      [7:0] n21453;
wire            n21454;
wire      [7:0] n21455;
wire            n21456;
wire      [7:0] n21457;
wire            n21458;
wire      [7:0] n21459;
wire            n2146;
wire            n21460;
wire      [7:0] n21461;
wire            n21462;
wire      [7:0] n21463;
wire            n21464;
wire      [7:0] n21465;
wire            n21466;
wire      [7:0] n21467;
wire            n21468;
wire      [7:0] n21469;
wire      [7:0] n2147;
wire            n21470;
wire      [7:0] n21471;
wire            n21472;
wire      [7:0] n21473;
wire            n21474;
wire      [7:0] n21475;
wire            n21476;
wire      [7:0] n21477;
wire            n21478;
wire      [7:0] n21479;
wire            n2148;
wire            n21480;
wire      [7:0] n21481;
wire            n21482;
wire      [7:0] n21483;
wire            n21484;
wire      [7:0] n21485;
wire            n21486;
wire      [7:0] n21487;
wire            n21488;
wire      [7:0] n21489;
wire      [7:0] n2149;
wire            n21490;
wire      [7:0] n21491;
wire            n21492;
wire      [7:0] n21493;
wire            n21494;
wire      [7:0] n21495;
wire            n21496;
wire      [7:0] n21497;
wire            n21498;
wire      [7:0] n21499;
wire      [7:0] n215;
wire            n2150;
wire            n21500;
wire      [7:0] n21501;
wire            n21502;
wire      [7:0] n21503;
wire            n21504;
wire      [7:0] n21505;
wire            n21506;
wire      [7:0] n21507;
wire            n21508;
wire      [7:0] n21509;
wire      [7:0] n2151;
wire            n21510;
wire      [7:0] n21511;
wire            n21512;
wire      [7:0] n21513;
wire            n21514;
wire      [7:0] n21515;
wire            n21516;
wire      [7:0] n21517;
wire            n21518;
wire      [7:0] n21519;
wire            n2152;
wire            n21520;
wire      [7:0] n21521;
wire            n21522;
wire      [7:0] n21523;
wire            n21524;
wire      [7:0] n21525;
wire            n21526;
wire      [7:0] n21527;
wire            n21528;
wire      [7:0] n21529;
wire      [7:0] n2153;
wire            n21530;
wire      [7:0] n21531;
wire            n21532;
wire      [7:0] n21533;
wire            n21534;
wire      [7:0] n21535;
wire            n21536;
wire      [7:0] n21537;
wire            n21538;
wire      [7:0] n21539;
wire            n2154;
wire            n21540;
wire      [7:0] n21541;
wire            n21542;
wire      [7:0] n21543;
wire            n21544;
wire      [7:0] n21545;
wire            n21546;
wire      [7:0] n21547;
wire            n21548;
wire      [7:0] n21549;
wire      [7:0] n2155;
wire            n21550;
wire      [7:0] n21551;
wire            n21552;
wire      [7:0] n21553;
wire            n21554;
wire      [7:0] n21555;
wire            n21556;
wire      [7:0] n21557;
wire            n21558;
wire      [7:0] n21559;
wire            n2156;
wire            n21560;
wire      [7:0] n21561;
wire            n21562;
wire      [7:0] n21563;
wire            n21564;
wire      [7:0] n21565;
wire            n21566;
wire      [7:0] n21567;
wire            n21568;
wire      [7:0] n21569;
wire      [7:0] n2157;
wire            n21570;
wire      [7:0] n21571;
wire            n21572;
wire      [7:0] n21573;
wire            n21574;
wire      [7:0] n21575;
wire            n21576;
wire      [7:0] n21577;
wire            n21578;
wire      [7:0] n21579;
wire            n2158;
wire            n21580;
wire      [7:0] n21581;
wire            n21582;
wire      [7:0] n21583;
wire            n21584;
wire      [7:0] n21585;
wire            n21586;
wire      [7:0] n21587;
wire            n21588;
wire      [7:0] n21589;
wire      [7:0] n2159;
wire            n21590;
wire      [7:0] n21591;
wire      [7:0] n21592;
wire      [7:0] n21593;
wire      [7:0] n21594;
wire      [7:0] n21595;
wire      [7:0] n21596;
wire      [7:0] n21597;
wire      [7:0] n21598;
wire      [7:0] n21599;
wire            n2160;
wire      [7:0] n21600;
wire      [7:0] n21601;
wire      [7:0] n21602;
wire      [7:0] n21603;
wire      [7:0] n21604;
wire      [7:0] n21605;
wire      [7:0] n21606;
wire      [7:0] n21607;
wire      [7:0] n21608;
wire      [7:0] n21609;
wire      [7:0] n2161;
wire      [7:0] n21610;
wire      [7:0] n21611;
wire      [7:0] n21612;
wire      [7:0] n21613;
wire      [7:0] n21614;
wire      [7:0] n21615;
wire      [7:0] n21616;
wire      [7:0] n21617;
wire      [7:0] n21618;
wire      [7:0] n21619;
wire            n2162;
wire      [7:0] n21620;
wire      [7:0] n21621;
wire      [7:0] n21622;
wire      [7:0] n21623;
wire      [7:0] n21624;
wire      [7:0] n21625;
wire      [7:0] n21626;
wire      [7:0] n21627;
wire      [7:0] n21628;
wire      [7:0] n21629;
wire      [7:0] n2163;
wire      [7:0] n21630;
wire      [7:0] n21631;
wire      [7:0] n21632;
wire      [7:0] n21633;
wire      [7:0] n21634;
wire      [7:0] n21635;
wire      [7:0] n21636;
wire      [7:0] n21637;
wire      [7:0] n21638;
wire      [7:0] n21639;
wire            n2164;
wire      [7:0] n21640;
wire      [7:0] n21641;
wire      [7:0] n21642;
wire      [7:0] n21643;
wire      [7:0] n21644;
wire      [7:0] n21645;
wire      [7:0] n21646;
wire      [7:0] n21647;
wire      [7:0] n21648;
wire      [7:0] n21649;
wire      [7:0] n2165;
wire      [7:0] n21650;
wire      [7:0] n21651;
wire      [7:0] n21652;
wire      [7:0] n21653;
wire      [7:0] n21654;
wire      [7:0] n21655;
wire      [7:0] n21656;
wire      [7:0] n21657;
wire      [7:0] n21658;
wire      [7:0] n21659;
wire            n2166;
wire      [7:0] n21660;
wire      [7:0] n21661;
wire      [7:0] n21662;
wire      [7:0] n21663;
wire      [7:0] n21664;
wire      [7:0] n21665;
wire      [7:0] n21666;
wire      [7:0] n21667;
wire      [7:0] n21668;
wire      [7:0] n21669;
wire      [7:0] n2167;
wire      [7:0] n21670;
wire      [7:0] n21671;
wire      [7:0] n21672;
wire      [7:0] n21673;
wire      [7:0] n21674;
wire      [7:0] n21675;
wire      [7:0] n21676;
wire      [7:0] n21677;
wire      [7:0] n21678;
wire      [7:0] n21679;
wire            n2168;
wire      [7:0] n21680;
wire      [7:0] n21681;
wire      [7:0] n21682;
wire      [7:0] n21683;
wire      [7:0] n21684;
wire      [7:0] n21685;
wire      [7:0] n21686;
wire      [7:0] n21687;
wire      [7:0] n21688;
wire      [7:0] n21689;
wire      [7:0] n2169;
wire      [7:0] n21690;
wire      [7:0] n21691;
wire      [7:0] n21692;
wire      [7:0] n21693;
wire      [7:0] n21694;
wire      [7:0] n21695;
wire      [7:0] n21696;
wire      [7:0] n21697;
wire      [7:0] n21698;
wire      [7:0] n21699;
wire            n217;
wire            n2170;
wire      [7:0] n21700;
wire      [7:0] n21701;
wire      [7:0] n21702;
wire      [7:0] n21703;
wire      [7:0] n21704;
wire      [7:0] n21705;
wire      [7:0] n21706;
wire      [7:0] n21707;
wire      [7:0] n21708;
wire      [7:0] n21709;
wire      [7:0] n2171;
wire      [7:0] n21710;
wire      [7:0] n21711;
wire      [7:0] n21712;
wire      [7:0] n21713;
wire      [7:0] n21714;
wire      [7:0] n21715;
wire      [7:0] n21716;
wire      [7:0] n21717;
wire      [7:0] n21718;
wire      [7:0] n21719;
wire            n2172;
wire      [7:0] n21720;
wire      [7:0] n21721;
wire      [7:0] n21722;
wire      [7:0] n21723;
wire      [7:0] n21724;
wire      [7:0] n21725;
wire      [7:0] n21726;
wire      [7:0] n21727;
wire      [7:0] n21728;
wire      [7:0] n21729;
wire      [7:0] n2173;
wire      [7:0] n21730;
wire      [7:0] n21731;
wire      [7:0] n21732;
wire      [7:0] n21733;
wire      [7:0] n21734;
wire      [7:0] n21735;
wire      [7:0] n21736;
wire      [7:0] n21737;
wire      [7:0] n21738;
wire      [7:0] n21739;
wire            n2174;
wire      [7:0] n21740;
wire      [7:0] n21741;
wire      [7:0] n21742;
wire      [7:0] n21743;
wire      [7:0] n21744;
wire      [7:0] n21745;
wire      [7:0] n21746;
wire      [7:0] n21747;
wire      [7:0] n21748;
wire      [7:0] n21749;
wire      [7:0] n2175;
wire      [7:0] n21750;
wire      [7:0] n21751;
wire      [7:0] n21752;
wire      [7:0] n21753;
wire      [7:0] n21754;
wire      [7:0] n21755;
wire      [7:0] n21756;
wire      [7:0] n21757;
wire      [7:0] n21758;
wire      [7:0] n21759;
wire            n2176;
wire      [7:0] n21760;
wire      [7:0] n21761;
wire      [7:0] n21762;
wire      [7:0] n21763;
wire      [7:0] n21764;
wire      [7:0] n21765;
wire      [7:0] n21766;
wire      [7:0] n21767;
wire      [7:0] n21768;
wire      [7:0] n21769;
wire      [7:0] n2177;
wire      [7:0] n21770;
wire      [7:0] n21771;
wire      [7:0] n21772;
wire      [7:0] n21773;
wire      [7:0] n21774;
wire      [7:0] n21775;
wire      [7:0] n21776;
wire      [7:0] n21777;
wire      [7:0] n21778;
wire      [7:0] n21779;
wire            n2178;
wire      [7:0] n21780;
wire      [7:0] n21781;
wire      [7:0] n21782;
wire      [7:0] n21783;
wire      [7:0] n21784;
wire      [7:0] n21785;
wire      [7:0] n21786;
wire      [7:0] n21787;
wire      [7:0] n21788;
wire      [7:0] n21789;
wire      [7:0] n2179;
wire      [7:0] n21790;
wire      [7:0] n21791;
wire      [7:0] n21792;
wire      [7:0] n21793;
wire      [7:0] n21794;
wire      [7:0] n21795;
wire      [7:0] n21796;
wire      [7:0] n21797;
wire      [7:0] n21798;
wire      [7:0] n21799;
wire            n2180;
wire      [7:0] n21800;
wire      [7:0] n21801;
wire      [7:0] n21802;
wire      [7:0] n21803;
wire      [7:0] n21804;
wire      [7:0] n21805;
wire      [7:0] n21806;
wire      [7:0] n21807;
wire      [7:0] n21808;
wire      [7:0] n21809;
wire      [7:0] n2181;
wire      [7:0] n21810;
wire      [7:0] n21811;
wire      [7:0] n21812;
wire      [7:0] n21813;
wire      [7:0] n21814;
wire      [7:0] n21815;
wire      [7:0] n21816;
wire      [7:0] n21817;
wire      [7:0] n21818;
wire      [7:0] n21819;
wire            n2182;
wire      [7:0] n21820;
wire      [7:0] n21821;
wire      [7:0] n21822;
wire      [7:0] n21823;
wire      [7:0] n21824;
wire      [7:0] n21825;
wire      [7:0] n21826;
wire      [7:0] n21827;
wire      [7:0] n21828;
wire      [7:0] n21829;
wire      [7:0] n2183;
wire      [7:0] n21830;
wire      [7:0] n21831;
wire      [7:0] n21832;
wire      [7:0] n21833;
wire      [7:0] n21834;
wire      [7:0] n21835;
wire      [7:0] n21836;
wire      [7:0] n21837;
wire      [7:0] n21838;
wire      [7:0] n21839;
wire            n2184;
wire      [7:0] n21840;
wire      [7:0] n21841;
wire      [7:0] n21842;
wire      [7:0] n21843;
wire      [7:0] n21844;
wire      [7:0] n21845;
wire      [7:0] n21846;
wire      [7:0] n21847;
wire      [7:0] n21848;
wire            n21849;
wire      [7:0] n2185;
wire      [7:0] n21850;
wire            n21851;
wire      [7:0] n21852;
wire            n21853;
wire      [7:0] n21854;
wire            n21855;
wire      [7:0] n21856;
wire            n21857;
wire      [7:0] n21858;
wire            n21859;
wire            n2186;
wire      [7:0] n21860;
wire            n21861;
wire      [7:0] n21862;
wire            n21863;
wire      [7:0] n21864;
wire            n21865;
wire      [7:0] n21866;
wire            n21867;
wire      [7:0] n21868;
wire            n21869;
wire      [7:0] n2187;
wire      [7:0] n21870;
wire            n21871;
wire      [7:0] n21872;
wire            n21873;
wire      [7:0] n21874;
wire            n21875;
wire      [7:0] n21876;
wire            n21877;
wire      [7:0] n21878;
wire            n21879;
wire            n2188;
wire      [7:0] n21880;
wire            n21881;
wire      [7:0] n21882;
wire            n21883;
wire      [7:0] n21884;
wire            n21885;
wire      [7:0] n21886;
wire            n21887;
wire      [7:0] n21888;
wire            n21889;
wire      [7:0] n2189;
wire      [7:0] n21890;
wire            n21891;
wire      [7:0] n21892;
wire            n21893;
wire      [7:0] n21894;
wire            n21895;
wire      [7:0] n21896;
wire            n21897;
wire      [7:0] n21898;
wire            n21899;
wire      [7:0] n219;
wire            n2190;
wire      [7:0] n21900;
wire            n21901;
wire      [7:0] n21902;
wire            n21903;
wire      [7:0] n21904;
wire            n21905;
wire      [7:0] n21906;
wire            n21907;
wire      [7:0] n21908;
wire            n21909;
wire      [7:0] n2191;
wire      [7:0] n21910;
wire            n21911;
wire      [7:0] n21912;
wire            n21913;
wire      [7:0] n21914;
wire            n21915;
wire      [7:0] n21916;
wire            n21917;
wire      [7:0] n21918;
wire            n21919;
wire            n2192;
wire      [7:0] n21920;
wire            n21921;
wire      [7:0] n21922;
wire            n21923;
wire      [7:0] n21924;
wire            n21925;
wire      [7:0] n21926;
wire            n21927;
wire      [7:0] n21928;
wire            n21929;
wire      [7:0] n2193;
wire      [7:0] n21930;
wire            n21931;
wire      [7:0] n21932;
wire            n21933;
wire      [7:0] n21934;
wire            n21935;
wire      [7:0] n21936;
wire            n21937;
wire      [7:0] n21938;
wire            n21939;
wire            n2194;
wire      [7:0] n21940;
wire            n21941;
wire      [7:0] n21942;
wire            n21943;
wire      [7:0] n21944;
wire            n21945;
wire      [7:0] n21946;
wire            n21947;
wire      [7:0] n21948;
wire            n21949;
wire      [7:0] n2195;
wire      [7:0] n21950;
wire            n21951;
wire      [7:0] n21952;
wire            n21953;
wire      [7:0] n21954;
wire            n21955;
wire      [7:0] n21956;
wire            n21957;
wire      [7:0] n21958;
wire            n21959;
wire            n2196;
wire      [7:0] n21960;
wire            n21961;
wire      [7:0] n21962;
wire            n21963;
wire      [7:0] n21964;
wire            n21965;
wire      [7:0] n21966;
wire            n21967;
wire      [7:0] n21968;
wire            n21969;
wire      [7:0] n2197;
wire      [7:0] n21970;
wire            n21971;
wire      [7:0] n21972;
wire            n21973;
wire      [7:0] n21974;
wire            n21975;
wire      [7:0] n21976;
wire            n21977;
wire      [7:0] n21978;
wire            n21979;
wire            n2198;
wire      [7:0] n21980;
wire            n21981;
wire      [7:0] n21982;
wire            n21983;
wire      [7:0] n21984;
wire            n21985;
wire      [7:0] n21986;
wire            n21987;
wire      [7:0] n21988;
wire            n21989;
wire      [7:0] n2199;
wire      [7:0] n21990;
wire            n21991;
wire      [7:0] n21992;
wire            n21993;
wire      [7:0] n21994;
wire            n21995;
wire      [7:0] n21996;
wire            n21997;
wire      [7:0] n21998;
wire            n21999;
wire      [7:0] n22;
wire            n2200;
wire      [7:0] n22000;
wire            n22001;
wire      [7:0] n22002;
wire            n22003;
wire      [7:0] n22004;
wire            n22005;
wire      [7:0] n22006;
wire            n22007;
wire      [7:0] n22008;
wire            n22009;
wire      [7:0] n2201;
wire      [7:0] n22010;
wire            n22011;
wire      [7:0] n22012;
wire            n22013;
wire      [7:0] n22014;
wire            n22015;
wire      [7:0] n22016;
wire            n22017;
wire      [7:0] n22018;
wire            n22019;
wire            n2202;
wire      [7:0] n22020;
wire            n22021;
wire      [7:0] n22022;
wire            n22023;
wire      [7:0] n22024;
wire            n22025;
wire      [7:0] n22026;
wire            n22027;
wire      [7:0] n22028;
wire            n22029;
wire      [7:0] n2203;
wire      [7:0] n22030;
wire            n22031;
wire      [7:0] n22032;
wire            n22033;
wire      [7:0] n22034;
wire            n22035;
wire      [7:0] n22036;
wire            n22037;
wire      [7:0] n22038;
wire            n22039;
wire            n2204;
wire      [7:0] n22040;
wire            n22041;
wire      [7:0] n22042;
wire            n22043;
wire      [7:0] n22044;
wire            n22045;
wire      [7:0] n22046;
wire            n22047;
wire      [7:0] n22048;
wire            n22049;
wire      [7:0] n2205;
wire      [7:0] n22050;
wire            n22051;
wire      [7:0] n22052;
wire            n22053;
wire      [7:0] n22054;
wire            n22055;
wire      [7:0] n22056;
wire            n22057;
wire      [7:0] n22058;
wire            n22059;
wire            n2206;
wire      [7:0] n22060;
wire            n22061;
wire      [7:0] n22062;
wire            n22063;
wire      [7:0] n22064;
wire            n22065;
wire      [7:0] n22066;
wire            n22067;
wire      [7:0] n22068;
wire            n22069;
wire      [7:0] n2207;
wire      [7:0] n22070;
wire            n22071;
wire      [7:0] n22072;
wire            n22073;
wire      [7:0] n22074;
wire            n22075;
wire      [7:0] n22076;
wire            n22077;
wire      [7:0] n22078;
wire            n22079;
wire            n2208;
wire      [7:0] n22080;
wire            n22081;
wire      [7:0] n22082;
wire            n22083;
wire      [7:0] n22084;
wire            n22085;
wire      [7:0] n22086;
wire            n22087;
wire      [7:0] n22088;
wire            n22089;
wire      [7:0] n2209;
wire      [7:0] n22090;
wire            n22091;
wire      [7:0] n22092;
wire            n22093;
wire      [7:0] n22094;
wire            n22095;
wire      [7:0] n22096;
wire            n22097;
wire      [7:0] n22098;
wire            n22099;
wire            n221;
wire            n2210;
wire      [7:0] n22100;
wire            n22101;
wire      [7:0] n22102;
wire            n22103;
wire      [7:0] n22104;
wire            n22105;
wire      [7:0] n22106;
wire            n22107;
wire      [7:0] n22108;
wire            n22109;
wire      [7:0] n2211;
wire      [7:0] n22110;
wire            n22111;
wire      [7:0] n22112;
wire            n22113;
wire      [7:0] n22114;
wire            n22115;
wire      [7:0] n22116;
wire            n22117;
wire      [7:0] n22118;
wire            n22119;
wire            n2212;
wire      [7:0] n22120;
wire            n22121;
wire      [7:0] n22122;
wire            n22123;
wire      [7:0] n22124;
wire            n22125;
wire      [7:0] n22126;
wire            n22127;
wire      [7:0] n22128;
wire            n22129;
wire      [7:0] n2213;
wire      [7:0] n22130;
wire            n22131;
wire      [7:0] n22132;
wire            n22133;
wire      [7:0] n22134;
wire            n22135;
wire      [7:0] n22136;
wire            n22137;
wire      [7:0] n22138;
wire            n22139;
wire            n2214;
wire      [7:0] n22140;
wire            n22141;
wire      [7:0] n22142;
wire            n22143;
wire      [7:0] n22144;
wire            n22145;
wire      [7:0] n22146;
wire            n22147;
wire      [7:0] n22148;
wire            n22149;
wire      [7:0] n2215;
wire      [7:0] n22150;
wire            n22151;
wire      [7:0] n22152;
wire            n22153;
wire      [7:0] n22154;
wire            n22155;
wire      [7:0] n22156;
wire            n22157;
wire      [7:0] n22158;
wire            n22159;
wire            n2216;
wire      [7:0] n22160;
wire            n22161;
wire      [7:0] n22162;
wire            n22163;
wire      [7:0] n22164;
wire            n22165;
wire      [7:0] n22166;
wire            n22167;
wire      [7:0] n22168;
wire            n22169;
wire      [7:0] n2217;
wire      [7:0] n22170;
wire            n22171;
wire      [7:0] n22172;
wire            n22173;
wire      [7:0] n22174;
wire            n22175;
wire      [7:0] n22176;
wire            n22177;
wire      [7:0] n22178;
wire            n22179;
wire            n2218;
wire      [7:0] n22180;
wire            n22181;
wire      [7:0] n22182;
wire            n22183;
wire      [7:0] n22184;
wire            n22185;
wire      [7:0] n22186;
wire            n22187;
wire      [7:0] n22188;
wire            n22189;
wire      [7:0] n2219;
wire      [7:0] n22190;
wire            n22191;
wire      [7:0] n22192;
wire            n22193;
wire      [7:0] n22194;
wire            n22195;
wire      [7:0] n22196;
wire            n22197;
wire      [7:0] n22198;
wire            n22199;
wire            n2220;
wire      [7:0] n22200;
wire            n22201;
wire      [7:0] n22202;
wire            n22203;
wire      [7:0] n22204;
wire            n22205;
wire      [7:0] n22206;
wire            n22207;
wire      [7:0] n22208;
wire            n22209;
wire      [7:0] n2221;
wire      [7:0] n22210;
wire            n22211;
wire      [7:0] n22212;
wire            n22213;
wire      [7:0] n22214;
wire            n22215;
wire      [7:0] n22216;
wire            n22217;
wire      [7:0] n22218;
wire            n22219;
wire            n2222;
wire      [7:0] n22220;
wire            n22221;
wire      [7:0] n22222;
wire            n22223;
wire      [7:0] n22224;
wire            n22225;
wire      [7:0] n22226;
wire            n22227;
wire      [7:0] n22228;
wire            n22229;
wire      [7:0] n2223;
wire      [7:0] n22230;
wire            n22231;
wire      [7:0] n22232;
wire            n22233;
wire      [7:0] n22234;
wire            n22235;
wire      [7:0] n22236;
wire            n22237;
wire      [7:0] n22238;
wire            n22239;
wire            n2224;
wire      [7:0] n22240;
wire            n22241;
wire      [7:0] n22242;
wire            n22243;
wire      [7:0] n22244;
wire            n22245;
wire      [7:0] n22246;
wire            n22247;
wire      [7:0] n22248;
wire            n22249;
wire      [7:0] n2225;
wire      [7:0] n22250;
wire            n22251;
wire      [7:0] n22252;
wire            n22253;
wire      [7:0] n22254;
wire            n22255;
wire      [7:0] n22256;
wire            n22257;
wire      [7:0] n22258;
wire            n22259;
wire            n2226;
wire      [7:0] n22260;
wire            n22261;
wire      [7:0] n22262;
wire            n22263;
wire      [7:0] n22264;
wire            n22265;
wire      [7:0] n22266;
wire            n22267;
wire      [7:0] n22268;
wire            n22269;
wire      [7:0] n2227;
wire      [7:0] n22270;
wire            n22271;
wire      [7:0] n22272;
wire            n22273;
wire      [7:0] n22274;
wire            n22275;
wire      [7:0] n22276;
wire            n22277;
wire      [7:0] n22278;
wire            n22279;
wire            n2228;
wire      [7:0] n22280;
wire            n22281;
wire      [7:0] n22282;
wire            n22283;
wire      [7:0] n22284;
wire            n22285;
wire      [7:0] n22286;
wire            n22287;
wire      [7:0] n22288;
wire            n22289;
wire      [7:0] n2229;
wire      [7:0] n22290;
wire            n22291;
wire      [7:0] n22292;
wire            n22293;
wire      [7:0] n22294;
wire            n22295;
wire      [7:0] n22296;
wire            n22297;
wire      [7:0] n22298;
wire            n22299;
wire      [7:0] n223;
wire            n2230;
wire      [7:0] n22300;
wire            n22301;
wire      [7:0] n22302;
wire            n22303;
wire      [7:0] n22304;
wire            n22305;
wire      [7:0] n22306;
wire            n22307;
wire      [7:0] n22308;
wire            n22309;
wire      [7:0] n2231;
wire      [7:0] n22310;
wire            n22311;
wire      [7:0] n22312;
wire            n22313;
wire      [7:0] n22314;
wire            n22315;
wire      [7:0] n22316;
wire            n22317;
wire      [7:0] n22318;
wire            n22319;
wire            n2232;
wire      [7:0] n22320;
wire            n22321;
wire      [7:0] n22322;
wire            n22323;
wire      [7:0] n22324;
wire            n22325;
wire      [7:0] n22326;
wire            n22327;
wire      [7:0] n22328;
wire            n22329;
wire      [7:0] n2233;
wire      [7:0] n22330;
wire            n22331;
wire      [7:0] n22332;
wire            n22333;
wire      [7:0] n22334;
wire            n22335;
wire      [7:0] n22336;
wire            n22337;
wire      [7:0] n22338;
wire            n22339;
wire            n2234;
wire      [7:0] n22340;
wire            n22341;
wire      [7:0] n22342;
wire            n22343;
wire      [7:0] n22344;
wire            n22345;
wire      [7:0] n22346;
wire            n22347;
wire      [7:0] n22348;
wire            n22349;
wire      [7:0] n2235;
wire      [7:0] n22350;
wire            n22351;
wire      [7:0] n22352;
wire            n22353;
wire      [7:0] n22354;
wire            n22355;
wire      [7:0] n22356;
wire            n22357;
wire      [7:0] n22358;
wire            n22359;
wire            n2236;
wire      [7:0] n22360;
wire      [7:0] n22361;
wire      [7:0] n22362;
wire      [7:0] n22363;
wire      [7:0] n22364;
wire      [7:0] n22365;
wire      [7:0] n22366;
wire      [7:0] n22367;
wire      [7:0] n22368;
wire      [7:0] n22369;
wire      [7:0] n2237;
wire      [7:0] n22370;
wire      [7:0] n22371;
wire      [7:0] n22372;
wire      [7:0] n22373;
wire      [7:0] n22374;
wire      [7:0] n22375;
wire      [7:0] n22376;
wire      [7:0] n22377;
wire      [7:0] n22378;
wire      [7:0] n22379;
wire            n2238;
wire      [7:0] n22380;
wire      [7:0] n22381;
wire      [7:0] n22382;
wire      [7:0] n22383;
wire      [7:0] n22384;
wire      [7:0] n22385;
wire      [7:0] n22386;
wire      [7:0] n22387;
wire      [7:0] n22388;
wire      [7:0] n22389;
wire      [7:0] n2239;
wire      [7:0] n22390;
wire      [7:0] n22391;
wire      [7:0] n22392;
wire      [7:0] n22393;
wire      [7:0] n22394;
wire      [7:0] n22395;
wire      [7:0] n22396;
wire      [7:0] n22397;
wire      [7:0] n22398;
wire      [7:0] n22399;
wire            n2240;
wire      [7:0] n22400;
wire      [7:0] n22401;
wire      [7:0] n22402;
wire      [7:0] n22403;
wire      [7:0] n22404;
wire      [7:0] n22405;
wire      [7:0] n22406;
wire      [7:0] n22407;
wire      [7:0] n22408;
wire      [7:0] n22409;
wire      [7:0] n2241;
wire      [7:0] n22410;
wire      [7:0] n22411;
wire      [7:0] n22412;
wire      [7:0] n22413;
wire      [7:0] n22414;
wire      [7:0] n22415;
wire      [7:0] n22416;
wire      [7:0] n22417;
wire      [7:0] n22418;
wire      [7:0] n22419;
wire            n2242;
wire      [7:0] n22420;
wire      [7:0] n22421;
wire      [7:0] n22422;
wire      [7:0] n22423;
wire      [7:0] n22424;
wire      [7:0] n22425;
wire      [7:0] n22426;
wire      [7:0] n22427;
wire      [7:0] n22428;
wire      [7:0] n22429;
wire      [7:0] n2243;
wire      [7:0] n22430;
wire      [7:0] n22431;
wire      [7:0] n22432;
wire      [7:0] n22433;
wire      [7:0] n22434;
wire      [7:0] n22435;
wire      [7:0] n22436;
wire      [7:0] n22437;
wire      [7:0] n22438;
wire      [7:0] n22439;
wire            n2244;
wire      [7:0] n22440;
wire      [7:0] n22441;
wire      [7:0] n22442;
wire      [7:0] n22443;
wire      [7:0] n22444;
wire      [7:0] n22445;
wire      [7:0] n22446;
wire      [7:0] n22447;
wire      [7:0] n22448;
wire      [7:0] n22449;
wire      [7:0] n2245;
wire      [7:0] n22450;
wire      [7:0] n22451;
wire      [7:0] n22452;
wire      [7:0] n22453;
wire      [7:0] n22454;
wire      [7:0] n22455;
wire      [7:0] n22456;
wire      [7:0] n22457;
wire      [7:0] n22458;
wire      [7:0] n22459;
wire            n2246;
wire      [7:0] n22460;
wire      [7:0] n22461;
wire      [7:0] n22462;
wire      [7:0] n22463;
wire      [7:0] n22464;
wire      [7:0] n22465;
wire      [7:0] n22466;
wire      [7:0] n22467;
wire      [7:0] n22468;
wire      [7:0] n22469;
wire      [7:0] n2247;
wire      [7:0] n22470;
wire      [7:0] n22471;
wire      [7:0] n22472;
wire      [7:0] n22473;
wire      [7:0] n22474;
wire      [7:0] n22475;
wire      [7:0] n22476;
wire      [7:0] n22477;
wire      [7:0] n22478;
wire      [7:0] n22479;
wire            n2248;
wire      [7:0] n22480;
wire      [7:0] n22481;
wire      [7:0] n22482;
wire      [7:0] n22483;
wire      [7:0] n22484;
wire      [7:0] n22485;
wire      [7:0] n22486;
wire      [7:0] n22487;
wire      [7:0] n22488;
wire      [7:0] n22489;
wire      [7:0] n2249;
wire      [7:0] n22490;
wire      [7:0] n22491;
wire      [7:0] n22492;
wire      [7:0] n22493;
wire      [7:0] n22494;
wire      [7:0] n22495;
wire      [7:0] n22496;
wire      [7:0] n22497;
wire      [7:0] n22498;
wire      [7:0] n22499;
wire            n225;
wire            n2250;
wire      [7:0] n22500;
wire      [7:0] n22501;
wire      [7:0] n22502;
wire      [7:0] n22503;
wire      [7:0] n22504;
wire      [7:0] n22505;
wire      [7:0] n22506;
wire      [7:0] n22507;
wire      [7:0] n22508;
wire      [7:0] n22509;
wire      [7:0] n2251;
wire      [7:0] n22510;
wire      [7:0] n22511;
wire      [7:0] n22512;
wire      [7:0] n22513;
wire      [7:0] n22514;
wire      [7:0] n22515;
wire      [7:0] n22516;
wire      [7:0] n22517;
wire      [7:0] n22518;
wire      [7:0] n22519;
wire            n2252;
wire      [7:0] n22520;
wire      [7:0] n22521;
wire      [7:0] n22522;
wire      [7:0] n22523;
wire      [7:0] n22524;
wire      [7:0] n22525;
wire      [7:0] n22526;
wire      [7:0] n22527;
wire      [7:0] n22528;
wire      [7:0] n22529;
wire      [7:0] n2253;
wire      [7:0] n22530;
wire      [7:0] n22531;
wire      [7:0] n22532;
wire      [7:0] n22533;
wire      [7:0] n22534;
wire      [7:0] n22535;
wire      [7:0] n22536;
wire      [7:0] n22537;
wire      [7:0] n22538;
wire      [7:0] n22539;
wire            n2254;
wire      [7:0] n22540;
wire      [7:0] n22541;
wire      [7:0] n22542;
wire      [7:0] n22543;
wire      [7:0] n22544;
wire      [7:0] n22545;
wire      [7:0] n22546;
wire      [7:0] n22547;
wire      [7:0] n22548;
wire      [7:0] n22549;
wire      [7:0] n2255;
wire      [7:0] n22550;
wire      [7:0] n22551;
wire      [7:0] n22552;
wire      [7:0] n22553;
wire      [7:0] n22554;
wire      [7:0] n22555;
wire      [7:0] n22556;
wire      [7:0] n22557;
wire      [7:0] n22558;
wire      [7:0] n22559;
wire            n2256;
wire      [7:0] n22560;
wire      [7:0] n22561;
wire      [7:0] n22562;
wire      [7:0] n22563;
wire      [7:0] n22564;
wire      [7:0] n22565;
wire      [7:0] n22566;
wire      [7:0] n22567;
wire      [7:0] n22568;
wire      [7:0] n22569;
wire      [7:0] n2257;
wire      [7:0] n22570;
wire      [7:0] n22571;
wire      [7:0] n22572;
wire      [7:0] n22573;
wire      [7:0] n22574;
wire      [7:0] n22575;
wire      [7:0] n22576;
wire      [7:0] n22577;
wire      [7:0] n22578;
wire      [7:0] n22579;
wire            n2258;
wire      [7:0] n22580;
wire      [7:0] n22581;
wire      [7:0] n22582;
wire      [7:0] n22583;
wire      [7:0] n22584;
wire      [7:0] n22585;
wire      [7:0] n22586;
wire      [7:0] n22587;
wire      [7:0] n22588;
wire      [7:0] n22589;
wire      [7:0] n2259;
wire      [7:0] n22590;
wire      [7:0] n22591;
wire      [7:0] n22592;
wire      [7:0] n22593;
wire      [7:0] n22594;
wire      [7:0] n22595;
wire      [7:0] n22596;
wire      [7:0] n22597;
wire      [7:0] n22598;
wire      [7:0] n22599;
wire            n2260;
wire      [7:0] n22600;
wire      [7:0] n22601;
wire      [7:0] n22602;
wire      [7:0] n22603;
wire      [7:0] n22604;
wire      [7:0] n22605;
wire      [7:0] n22606;
wire      [7:0] n22607;
wire      [7:0] n22608;
wire      [7:0] n22609;
wire      [7:0] n2261;
wire      [7:0] n22610;
wire      [7:0] n22611;
wire      [7:0] n22612;
wire      [7:0] n22613;
wire      [7:0] n22614;
wire      [7:0] n22615;
wire      [7:0] n22616;
wire      [7:0] n22617;
wire      [7:0] n22618;
wire    [103:0] n22619;
wire            n2262;
wire      [7:0] n22620;
wire      [7:0] n22621;
wire            n22622;
wire      [7:0] n22623;
wire            n22624;
wire      [7:0] n22625;
wire            n22626;
wire      [7:0] n22627;
wire            n22628;
wire      [7:0] n22629;
wire      [7:0] n2263;
wire            n22630;
wire      [7:0] n22631;
wire            n22632;
wire      [7:0] n22633;
wire            n22634;
wire      [7:0] n22635;
wire            n22636;
wire      [7:0] n22637;
wire            n22638;
wire      [7:0] n22639;
wire            n2264;
wire            n22640;
wire      [7:0] n22641;
wire            n22642;
wire      [7:0] n22643;
wire            n22644;
wire      [7:0] n22645;
wire            n22646;
wire      [7:0] n22647;
wire            n22648;
wire      [7:0] n22649;
wire      [7:0] n2265;
wire            n22650;
wire      [7:0] n22651;
wire            n22652;
wire      [7:0] n22653;
wire            n22654;
wire      [7:0] n22655;
wire            n22656;
wire      [7:0] n22657;
wire            n22658;
wire      [7:0] n22659;
wire            n2266;
wire            n22660;
wire      [7:0] n22661;
wire            n22662;
wire      [7:0] n22663;
wire            n22664;
wire      [7:0] n22665;
wire            n22666;
wire      [7:0] n22667;
wire            n22668;
wire      [7:0] n22669;
wire      [7:0] n2267;
wire            n22670;
wire      [7:0] n22671;
wire            n22672;
wire      [7:0] n22673;
wire            n22674;
wire      [7:0] n22675;
wire            n22676;
wire      [7:0] n22677;
wire            n22678;
wire      [7:0] n22679;
wire            n2268;
wire            n22680;
wire      [7:0] n22681;
wire            n22682;
wire      [7:0] n22683;
wire            n22684;
wire      [7:0] n22685;
wire            n22686;
wire      [7:0] n22687;
wire            n22688;
wire      [7:0] n22689;
wire      [7:0] n2269;
wire            n22690;
wire      [7:0] n22691;
wire            n22692;
wire      [7:0] n22693;
wire            n22694;
wire      [7:0] n22695;
wire            n22696;
wire      [7:0] n22697;
wire            n22698;
wire      [7:0] n22699;
wire      [7:0] n227;
wire            n2270;
wire            n22700;
wire      [7:0] n22701;
wire            n22702;
wire      [7:0] n22703;
wire            n22704;
wire      [7:0] n22705;
wire            n22706;
wire      [7:0] n22707;
wire            n22708;
wire      [7:0] n22709;
wire      [7:0] n2271;
wire            n22710;
wire      [7:0] n22711;
wire            n22712;
wire      [7:0] n22713;
wire            n22714;
wire      [7:0] n22715;
wire            n22716;
wire      [7:0] n22717;
wire            n22718;
wire      [7:0] n22719;
wire            n2272;
wire            n22720;
wire      [7:0] n22721;
wire            n22722;
wire      [7:0] n22723;
wire            n22724;
wire      [7:0] n22725;
wire            n22726;
wire      [7:0] n22727;
wire            n22728;
wire      [7:0] n22729;
wire      [7:0] n2273;
wire            n22730;
wire      [7:0] n22731;
wire            n22732;
wire      [7:0] n22733;
wire            n22734;
wire      [7:0] n22735;
wire            n22736;
wire      [7:0] n22737;
wire            n22738;
wire      [7:0] n22739;
wire            n2274;
wire            n22740;
wire      [7:0] n22741;
wire            n22742;
wire      [7:0] n22743;
wire            n22744;
wire      [7:0] n22745;
wire            n22746;
wire      [7:0] n22747;
wire            n22748;
wire      [7:0] n22749;
wire      [7:0] n2275;
wire            n22750;
wire      [7:0] n22751;
wire            n22752;
wire      [7:0] n22753;
wire            n22754;
wire      [7:0] n22755;
wire            n22756;
wire      [7:0] n22757;
wire            n22758;
wire      [7:0] n22759;
wire            n2276;
wire            n22760;
wire      [7:0] n22761;
wire            n22762;
wire      [7:0] n22763;
wire            n22764;
wire      [7:0] n22765;
wire            n22766;
wire      [7:0] n22767;
wire            n22768;
wire      [7:0] n22769;
wire      [7:0] n2277;
wire            n22770;
wire      [7:0] n22771;
wire            n22772;
wire      [7:0] n22773;
wire            n22774;
wire      [7:0] n22775;
wire            n22776;
wire      [7:0] n22777;
wire            n22778;
wire      [7:0] n22779;
wire            n2278;
wire            n22780;
wire      [7:0] n22781;
wire            n22782;
wire      [7:0] n22783;
wire            n22784;
wire      [7:0] n22785;
wire            n22786;
wire      [7:0] n22787;
wire            n22788;
wire      [7:0] n22789;
wire      [7:0] n2279;
wire            n22790;
wire      [7:0] n22791;
wire            n22792;
wire      [7:0] n22793;
wire            n22794;
wire      [7:0] n22795;
wire            n22796;
wire      [7:0] n22797;
wire            n22798;
wire      [7:0] n22799;
wire            n2280;
wire            n22800;
wire      [7:0] n22801;
wire            n22802;
wire      [7:0] n22803;
wire            n22804;
wire      [7:0] n22805;
wire            n22806;
wire      [7:0] n22807;
wire            n22808;
wire      [7:0] n22809;
wire      [7:0] n2281;
wire            n22810;
wire      [7:0] n22811;
wire            n22812;
wire      [7:0] n22813;
wire            n22814;
wire      [7:0] n22815;
wire            n22816;
wire      [7:0] n22817;
wire            n22818;
wire      [7:0] n22819;
wire            n2282;
wire            n22820;
wire      [7:0] n22821;
wire            n22822;
wire      [7:0] n22823;
wire            n22824;
wire      [7:0] n22825;
wire            n22826;
wire      [7:0] n22827;
wire            n22828;
wire      [7:0] n22829;
wire      [7:0] n2283;
wire            n22830;
wire      [7:0] n22831;
wire            n22832;
wire      [7:0] n22833;
wire            n22834;
wire      [7:0] n22835;
wire            n22836;
wire      [7:0] n22837;
wire            n22838;
wire      [7:0] n22839;
wire            n2284;
wire            n22840;
wire      [7:0] n22841;
wire            n22842;
wire      [7:0] n22843;
wire            n22844;
wire      [7:0] n22845;
wire            n22846;
wire      [7:0] n22847;
wire            n22848;
wire      [7:0] n22849;
wire      [7:0] n2285;
wire            n22850;
wire      [7:0] n22851;
wire            n22852;
wire      [7:0] n22853;
wire            n22854;
wire      [7:0] n22855;
wire            n22856;
wire      [7:0] n22857;
wire            n22858;
wire      [7:0] n22859;
wire            n2286;
wire            n22860;
wire      [7:0] n22861;
wire            n22862;
wire      [7:0] n22863;
wire            n22864;
wire      [7:0] n22865;
wire            n22866;
wire      [7:0] n22867;
wire            n22868;
wire      [7:0] n22869;
wire      [7:0] n2287;
wire            n22870;
wire      [7:0] n22871;
wire            n22872;
wire      [7:0] n22873;
wire            n22874;
wire      [7:0] n22875;
wire            n22876;
wire      [7:0] n22877;
wire            n22878;
wire      [7:0] n22879;
wire            n2288;
wire            n22880;
wire      [7:0] n22881;
wire            n22882;
wire      [7:0] n22883;
wire            n22884;
wire      [7:0] n22885;
wire            n22886;
wire      [7:0] n22887;
wire            n22888;
wire      [7:0] n22889;
wire      [7:0] n2289;
wire            n22890;
wire      [7:0] n22891;
wire            n22892;
wire      [7:0] n22893;
wire            n22894;
wire      [7:0] n22895;
wire            n22896;
wire      [7:0] n22897;
wire            n22898;
wire      [7:0] n22899;
wire            n229;
wire            n2290;
wire            n22900;
wire      [7:0] n22901;
wire            n22902;
wire      [7:0] n22903;
wire            n22904;
wire      [7:0] n22905;
wire            n22906;
wire      [7:0] n22907;
wire            n22908;
wire      [7:0] n22909;
wire      [7:0] n2291;
wire            n22910;
wire      [7:0] n22911;
wire            n22912;
wire      [7:0] n22913;
wire            n22914;
wire      [7:0] n22915;
wire            n22916;
wire      [7:0] n22917;
wire            n22918;
wire      [7:0] n22919;
wire            n2292;
wire            n22920;
wire      [7:0] n22921;
wire            n22922;
wire      [7:0] n22923;
wire            n22924;
wire      [7:0] n22925;
wire            n22926;
wire      [7:0] n22927;
wire            n22928;
wire      [7:0] n22929;
wire      [7:0] n2293;
wire            n22930;
wire      [7:0] n22931;
wire            n22932;
wire      [7:0] n22933;
wire            n22934;
wire      [7:0] n22935;
wire            n22936;
wire      [7:0] n22937;
wire            n22938;
wire      [7:0] n22939;
wire            n2294;
wire            n22940;
wire      [7:0] n22941;
wire            n22942;
wire      [7:0] n22943;
wire            n22944;
wire      [7:0] n22945;
wire            n22946;
wire      [7:0] n22947;
wire            n22948;
wire      [7:0] n22949;
wire      [7:0] n2295;
wire            n22950;
wire      [7:0] n22951;
wire            n22952;
wire      [7:0] n22953;
wire            n22954;
wire      [7:0] n22955;
wire            n22956;
wire      [7:0] n22957;
wire            n22958;
wire      [7:0] n22959;
wire            n2296;
wire            n22960;
wire      [7:0] n22961;
wire            n22962;
wire      [7:0] n22963;
wire            n22964;
wire      [7:0] n22965;
wire            n22966;
wire      [7:0] n22967;
wire            n22968;
wire      [7:0] n22969;
wire      [7:0] n2297;
wire            n22970;
wire      [7:0] n22971;
wire            n22972;
wire      [7:0] n22973;
wire            n22974;
wire      [7:0] n22975;
wire            n22976;
wire      [7:0] n22977;
wire            n22978;
wire      [7:0] n22979;
wire            n2298;
wire            n22980;
wire      [7:0] n22981;
wire            n22982;
wire      [7:0] n22983;
wire            n22984;
wire      [7:0] n22985;
wire            n22986;
wire      [7:0] n22987;
wire            n22988;
wire      [7:0] n22989;
wire      [7:0] n2299;
wire            n22990;
wire      [7:0] n22991;
wire            n22992;
wire      [7:0] n22993;
wire            n22994;
wire      [7:0] n22995;
wire            n22996;
wire      [7:0] n22997;
wire            n22998;
wire      [7:0] n22999;
wire            n2300;
wire            n23000;
wire      [7:0] n23001;
wire            n23002;
wire      [7:0] n23003;
wire            n23004;
wire      [7:0] n23005;
wire            n23006;
wire      [7:0] n23007;
wire            n23008;
wire      [7:0] n23009;
wire      [7:0] n2301;
wire            n23010;
wire      [7:0] n23011;
wire            n23012;
wire      [7:0] n23013;
wire            n23014;
wire      [7:0] n23015;
wire            n23016;
wire      [7:0] n23017;
wire            n23018;
wire      [7:0] n23019;
wire            n2302;
wire            n23020;
wire      [7:0] n23021;
wire            n23022;
wire      [7:0] n23023;
wire            n23024;
wire      [7:0] n23025;
wire            n23026;
wire      [7:0] n23027;
wire            n23028;
wire      [7:0] n23029;
wire      [7:0] n2303;
wire            n23030;
wire      [7:0] n23031;
wire            n23032;
wire      [7:0] n23033;
wire            n23034;
wire      [7:0] n23035;
wire            n23036;
wire      [7:0] n23037;
wire            n23038;
wire      [7:0] n23039;
wire            n2304;
wire            n23040;
wire      [7:0] n23041;
wire            n23042;
wire      [7:0] n23043;
wire            n23044;
wire      [7:0] n23045;
wire            n23046;
wire      [7:0] n23047;
wire            n23048;
wire      [7:0] n23049;
wire      [7:0] n2305;
wire            n23050;
wire      [7:0] n23051;
wire            n23052;
wire      [7:0] n23053;
wire            n23054;
wire      [7:0] n23055;
wire            n23056;
wire      [7:0] n23057;
wire            n23058;
wire      [7:0] n23059;
wire            n2306;
wire            n23060;
wire      [7:0] n23061;
wire            n23062;
wire      [7:0] n23063;
wire            n23064;
wire      [7:0] n23065;
wire            n23066;
wire      [7:0] n23067;
wire            n23068;
wire      [7:0] n23069;
wire      [7:0] n2307;
wire            n23070;
wire      [7:0] n23071;
wire            n23072;
wire      [7:0] n23073;
wire            n23074;
wire      [7:0] n23075;
wire            n23076;
wire      [7:0] n23077;
wire            n23078;
wire      [7:0] n23079;
wire      [7:0] n2308;
wire            n23080;
wire      [7:0] n23081;
wire            n23082;
wire      [7:0] n23083;
wire            n23084;
wire      [7:0] n23085;
wire            n23086;
wire      [7:0] n23087;
wire            n23088;
wire      [7:0] n23089;
wire      [7:0] n2309;
wire            n23090;
wire      [7:0] n23091;
wire            n23092;
wire      [7:0] n23093;
wire            n23094;
wire      [7:0] n23095;
wire            n23096;
wire      [7:0] n23097;
wire            n23098;
wire      [7:0] n23099;
wire      [7:0] n231;
wire      [7:0] n2310;
wire            n23100;
wire      [7:0] n23101;
wire            n23102;
wire      [7:0] n23103;
wire            n23104;
wire      [7:0] n23105;
wire            n23106;
wire      [7:0] n23107;
wire            n23108;
wire      [7:0] n23109;
wire      [7:0] n2311;
wire            n23110;
wire      [7:0] n23111;
wire            n23112;
wire      [7:0] n23113;
wire            n23114;
wire      [7:0] n23115;
wire            n23116;
wire      [7:0] n23117;
wire            n23118;
wire      [7:0] n23119;
wire      [7:0] n2312;
wire            n23120;
wire      [7:0] n23121;
wire            n23122;
wire      [7:0] n23123;
wire            n23124;
wire      [7:0] n23125;
wire            n23126;
wire      [7:0] n23127;
wire            n23128;
wire      [7:0] n23129;
wire      [7:0] n2313;
wire            n23130;
wire      [7:0] n23131;
wire            n23132;
wire      [7:0] n23133;
wire      [7:0] n23134;
wire      [7:0] n23135;
wire      [7:0] n23136;
wire      [7:0] n23137;
wire      [7:0] n23138;
wire      [7:0] n23139;
wire      [7:0] n2314;
wire      [7:0] n23140;
wire      [7:0] n23141;
wire      [7:0] n23142;
wire      [7:0] n23143;
wire      [7:0] n23144;
wire      [7:0] n23145;
wire      [7:0] n23146;
wire      [7:0] n23147;
wire      [7:0] n23148;
wire      [7:0] n23149;
wire      [7:0] n2315;
wire      [7:0] n23150;
wire      [7:0] n23151;
wire      [7:0] n23152;
wire      [7:0] n23153;
wire      [7:0] n23154;
wire      [7:0] n23155;
wire      [7:0] n23156;
wire      [7:0] n23157;
wire      [7:0] n23158;
wire      [7:0] n23159;
wire      [7:0] n2316;
wire      [7:0] n23160;
wire      [7:0] n23161;
wire      [7:0] n23162;
wire      [7:0] n23163;
wire      [7:0] n23164;
wire      [7:0] n23165;
wire      [7:0] n23166;
wire      [7:0] n23167;
wire      [7:0] n23168;
wire      [7:0] n23169;
wire      [7:0] n2317;
wire      [7:0] n23170;
wire      [7:0] n23171;
wire      [7:0] n23172;
wire      [7:0] n23173;
wire      [7:0] n23174;
wire      [7:0] n23175;
wire      [7:0] n23176;
wire      [7:0] n23177;
wire      [7:0] n23178;
wire      [7:0] n23179;
wire      [7:0] n2318;
wire      [7:0] n23180;
wire      [7:0] n23181;
wire      [7:0] n23182;
wire      [7:0] n23183;
wire      [7:0] n23184;
wire      [7:0] n23185;
wire      [7:0] n23186;
wire      [7:0] n23187;
wire      [7:0] n23188;
wire      [7:0] n23189;
wire      [7:0] n2319;
wire      [7:0] n23190;
wire      [7:0] n23191;
wire      [7:0] n23192;
wire      [7:0] n23193;
wire      [7:0] n23194;
wire      [7:0] n23195;
wire      [7:0] n23196;
wire      [7:0] n23197;
wire      [7:0] n23198;
wire      [7:0] n23199;
wire      [7:0] n2320;
wire      [7:0] n23200;
wire      [7:0] n23201;
wire      [7:0] n23202;
wire      [7:0] n23203;
wire      [7:0] n23204;
wire      [7:0] n23205;
wire      [7:0] n23206;
wire      [7:0] n23207;
wire      [7:0] n23208;
wire      [7:0] n23209;
wire      [7:0] n2321;
wire      [7:0] n23210;
wire      [7:0] n23211;
wire      [7:0] n23212;
wire      [7:0] n23213;
wire      [7:0] n23214;
wire      [7:0] n23215;
wire      [7:0] n23216;
wire      [7:0] n23217;
wire      [7:0] n23218;
wire      [7:0] n23219;
wire      [7:0] n2322;
wire      [7:0] n23220;
wire      [7:0] n23221;
wire      [7:0] n23222;
wire      [7:0] n23223;
wire      [7:0] n23224;
wire      [7:0] n23225;
wire      [7:0] n23226;
wire      [7:0] n23227;
wire      [7:0] n23228;
wire      [7:0] n23229;
wire      [7:0] n2323;
wire      [7:0] n23230;
wire      [7:0] n23231;
wire      [7:0] n23232;
wire      [7:0] n23233;
wire      [7:0] n23234;
wire      [7:0] n23235;
wire      [7:0] n23236;
wire      [7:0] n23237;
wire      [7:0] n23238;
wire      [7:0] n23239;
wire      [7:0] n2324;
wire      [7:0] n23240;
wire      [7:0] n23241;
wire      [7:0] n23242;
wire      [7:0] n23243;
wire      [7:0] n23244;
wire      [7:0] n23245;
wire      [7:0] n23246;
wire      [7:0] n23247;
wire      [7:0] n23248;
wire      [7:0] n23249;
wire      [7:0] n2325;
wire      [7:0] n23250;
wire      [7:0] n23251;
wire      [7:0] n23252;
wire      [7:0] n23253;
wire      [7:0] n23254;
wire      [7:0] n23255;
wire      [7:0] n23256;
wire      [7:0] n23257;
wire      [7:0] n23258;
wire      [7:0] n23259;
wire      [7:0] n2326;
wire      [7:0] n23260;
wire      [7:0] n23261;
wire      [7:0] n23262;
wire      [7:0] n23263;
wire      [7:0] n23264;
wire      [7:0] n23265;
wire      [7:0] n23266;
wire      [7:0] n23267;
wire      [7:0] n23268;
wire      [7:0] n23269;
wire      [7:0] n2327;
wire      [7:0] n23270;
wire      [7:0] n23271;
wire      [7:0] n23272;
wire      [7:0] n23273;
wire      [7:0] n23274;
wire      [7:0] n23275;
wire      [7:0] n23276;
wire      [7:0] n23277;
wire      [7:0] n23278;
wire      [7:0] n23279;
wire      [7:0] n2328;
wire      [7:0] n23280;
wire      [7:0] n23281;
wire      [7:0] n23282;
wire      [7:0] n23283;
wire      [7:0] n23284;
wire      [7:0] n23285;
wire      [7:0] n23286;
wire      [7:0] n23287;
wire      [7:0] n23288;
wire      [7:0] n23289;
wire      [7:0] n2329;
wire      [7:0] n23290;
wire      [7:0] n23291;
wire      [7:0] n23292;
wire      [7:0] n23293;
wire      [7:0] n23294;
wire      [7:0] n23295;
wire      [7:0] n23296;
wire      [7:0] n23297;
wire      [7:0] n23298;
wire      [7:0] n23299;
wire            n233;
wire      [7:0] n2330;
wire      [7:0] n23300;
wire      [7:0] n23301;
wire      [7:0] n23302;
wire      [7:0] n23303;
wire      [7:0] n23304;
wire      [7:0] n23305;
wire      [7:0] n23306;
wire      [7:0] n23307;
wire      [7:0] n23308;
wire      [7:0] n23309;
wire      [7:0] n2331;
wire      [7:0] n23310;
wire      [7:0] n23311;
wire      [7:0] n23312;
wire      [7:0] n23313;
wire      [7:0] n23314;
wire      [7:0] n23315;
wire      [7:0] n23316;
wire      [7:0] n23317;
wire      [7:0] n23318;
wire      [7:0] n23319;
wire      [7:0] n2332;
wire      [7:0] n23320;
wire      [7:0] n23321;
wire      [7:0] n23322;
wire      [7:0] n23323;
wire      [7:0] n23324;
wire      [7:0] n23325;
wire      [7:0] n23326;
wire      [7:0] n23327;
wire      [7:0] n23328;
wire      [7:0] n23329;
wire      [7:0] n2333;
wire      [7:0] n23330;
wire      [7:0] n23331;
wire      [7:0] n23332;
wire      [7:0] n23333;
wire      [7:0] n23334;
wire      [7:0] n23335;
wire      [7:0] n23336;
wire      [7:0] n23337;
wire      [7:0] n23338;
wire      [7:0] n23339;
wire      [7:0] n2334;
wire      [7:0] n23340;
wire      [7:0] n23341;
wire      [7:0] n23342;
wire      [7:0] n23343;
wire      [7:0] n23344;
wire      [7:0] n23345;
wire      [7:0] n23346;
wire      [7:0] n23347;
wire      [7:0] n23348;
wire      [7:0] n23349;
wire      [7:0] n2335;
wire      [7:0] n23350;
wire      [7:0] n23351;
wire      [7:0] n23352;
wire      [7:0] n23353;
wire      [7:0] n23354;
wire      [7:0] n23355;
wire      [7:0] n23356;
wire      [7:0] n23357;
wire      [7:0] n23358;
wire      [7:0] n23359;
wire      [7:0] n2336;
wire      [7:0] n23360;
wire      [7:0] n23361;
wire      [7:0] n23362;
wire      [7:0] n23363;
wire      [7:0] n23364;
wire      [7:0] n23365;
wire      [7:0] n23366;
wire      [7:0] n23367;
wire      [7:0] n23368;
wire      [7:0] n23369;
wire      [7:0] n2337;
wire      [7:0] n23370;
wire      [7:0] n23371;
wire      [7:0] n23372;
wire      [7:0] n23373;
wire      [7:0] n23374;
wire      [7:0] n23375;
wire      [7:0] n23376;
wire      [7:0] n23377;
wire      [7:0] n23378;
wire      [7:0] n23379;
wire      [7:0] n2338;
wire      [7:0] n23380;
wire      [7:0] n23381;
wire      [7:0] n23382;
wire      [7:0] n23383;
wire      [7:0] n23384;
wire      [7:0] n23385;
wire      [7:0] n23386;
wire      [7:0] n23387;
wire      [7:0] n23388;
wire      [7:0] n23389;
wire      [7:0] n2339;
wire      [7:0] n23390;
wire      [7:0] n23391;
wire            n23392;
wire      [7:0] n23393;
wire            n23394;
wire      [7:0] n23395;
wire            n23396;
wire      [7:0] n23397;
wire            n23398;
wire      [7:0] n23399;
wire      [7:0] n2340;
wire            n23400;
wire      [7:0] n23401;
wire            n23402;
wire      [7:0] n23403;
wire            n23404;
wire      [7:0] n23405;
wire            n23406;
wire      [7:0] n23407;
wire            n23408;
wire      [7:0] n23409;
wire      [7:0] n2341;
wire            n23410;
wire      [7:0] n23411;
wire            n23412;
wire      [7:0] n23413;
wire            n23414;
wire      [7:0] n23415;
wire            n23416;
wire      [7:0] n23417;
wire            n23418;
wire      [7:0] n23419;
wire      [7:0] n2342;
wire            n23420;
wire      [7:0] n23421;
wire            n23422;
wire      [7:0] n23423;
wire            n23424;
wire      [7:0] n23425;
wire            n23426;
wire      [7:0] n23427;
wire            n23428;
wire      [7:0] n23429;
wire      [7:0] n2343;
wire            n23430;
wire      [7:0] n23431;
wire            n23432;
wire      [7:0] n23433;
wire            n23434;
wire      [7:0] n23435;
wire            n23436;
wire      [7:0] n23437;
wire            n23438;
wire      [7:0] n23439;
wire      [7:0] n2344;
wire            n23440;
wire      [7:0] n23441;
wire            n23442;
wire      [7:0] n23443;
wire            n23444;
wire      [7:0] n23445;
wire            n23446;
wire      [7:0] n23447;
wire            n23448;
wire      [7:0] n23449;
wire      [7:0] n2345;
wire            n23450;
wire      [7:0] n23451;
wire            n23452;
wire      [7:0] n23453;
wire            n23454;
wire      [7:0] n23455;
wire            n23456;
wire      [7:0] n23457;
wire            n23458;
wire      [7:0] n23459;
wire      [7:0] n2346;
wire            n23460;
wire      [7:0] n23461;
wire            n23462;
wire      [7:0] n23463;
wire            n23464;
wire      [7:0] n23465;
wire            n23466;
wire      [7:0] n23467;
wire            n23468;
wire      [7:0] n23469;
wire      [7:0] n2347;
wire            n23470;
wire      [7:0] n23471;
wire            n23472;
wire      [7:0] n23473;
wire            n23474;
wire      [7:0] n23475;
wire            n23476;
wire      [7:0] n23477;
wire            n23478;
wire      [7:0] n23479;
wire      [7:0] n2348;
wire            n23480;
wire      [7:0] n23481;
wire            n23482;
wire      [7:0] n23483;
wire            n23484;
wire      [7:0] n23485;
wire            n23486;
wire      [7:0] n23487;
wire            n23488;
wire      [7:0] n23489;
wire      [7:0] n2349;
wire            n23490;
wire      [7:0] n23491;
wire            n23492;
wire      [7:0] n23493;
wire            n23494;
wire      [7:0] n23495;
wire            n23496;
wire      [7:0] n23497;
wire            n23498;
wire      [7:0] n23499;
wire      [7:0] n235;
wire      [7:0] n2350;
wire            n23500;
wire      [7:0] n23501;
wire            n23502;
wire      [7:0] n23503;
wire            n23504;
wire      [7:0] n23505;
wire            n23506;
wire      [7:0] n23507;
wire            n23508;
wire      [7:0] n23509;
wire      [7:0] n2351;
wire            n23510;
wire      [7:0] n23511;
wire            n23512;
wire      [7:0] n23513;
wire            n23514;
wire      [7:0] n23515;
wire            n23516;
wire      [7:0] n23517;
wire            n23518;
wire      [7:0] n23519;
wire      [7:0] n2352;
wire            n23520;
wire      [7:0] n23521;
wire            n23522;
wire      [7:0] n23523;
wire            n23524;
wire      [7:0] n23525;
wire            n23526;
wire      [7:0] n23527;
wire            n23528;
wire      [7:0] n23529;
wire      [7:0] n2353;
wire            n23530;
wire      [7:0] n23531;
wire            n23532;
wire      [7:0] n23533;
wire            n23534;
wire      [7:0] n23535;
wire            n23536;
wire      [7:0] n23537;
wire            n23538;
wire      [7:0] n23539;
wire      [7:0] n2354;
wire            n23540;
wire      [7:0] n23541;
wire            n23542;
wire      [7:0] n23543;
wire            n23544;
wire      [7:0] n23545;
wire            n23546;
wire      [7:0] n23547;
wire            n23548;
wire      [7:0] n23549;
wire      [7:0] n2355;
wire            n23550;
wire      [7:0] n23551;
wire            n23552;
wire      [7:0] n23553;
wire            n23554;
wire      [7:0] n23555;
wire            n23556;
wire      [7:0] n23557;
wire            n23558;
wire      [7:0] n23559;
wire      [7:0] n2356;
wire            n23560;
wire      [7:0] n23561;
wire            n23562;
wire      [7:0] n23563;
wire            n23564;
wire      [7:0] n23565;
wire            n23566;
wire      [7:0] n23567;
wire            n23568;
wire      [7:0] n23569;
wire      [7:0] n2357;
wire            n23570;
wire      [7:0] n23571;
wire            n23572;
wire      [7:0] n23573;
wire            n23574;
wire      [7:0] n23575;
wire            n23576;
wire      [7:0] n23577;
wire            n23578;
wire      [7:0] n23579;
wire      [7:0] n2358;
wire            n23580;
wire      [7:0] n23581;
wire            n23582;
wire      [7:0] n23583;
wire            n23584;
wire      [7:0] n23585;
wire            n23586;
wire      [7:0] n23587;
wire            n23588;
wire      [7:0] n23589;
wire      [7:0] n2359;
wire            n23590;
wire      [7:0] n23591;
wire            n23592;
wire      [7:0] n23593;
wire            n23594;
wire      [7:0] n23595;
wire            n23596;
wire      [7:0] n23597;
wire            n23598;
wire      [7:0] n23599;
wire            n236;
wire      [7:0] n2360;
wire            n23600;
wire      [7:0] n23601;
wire            n23602;
wire      [7:0] n23603;
wire            n23604;
wire      [7:0] n23605;
wire            n23606;
wire      [7:0] n23607;
wire            n23608;
wire      [7:0] n23609;
wire      [7:0] n2361;
wire            n23610;
wire      [7:0] n23611;
wire            n23612;
wire      [7:0] n23613;
wire            n23614;
wire      [7:0] n23615;
wire            n23616;
wire      [7:0] n23617;
wire            n23618;
wire      [7:0] n23619;
wire      [7:0] n2362;
wire            n23620;
wire      [7:0] n23621;
wire            n23622;
wire      [7:0] n23623;
wire            n23624;
wire      [7:0] n23625;
wire            n23626;
wire      [7:0] n23627;
wire            n23628;
wire      [7:0] n23629;
wire      [7:0] n2363;
wire            n23630;
wire      [7:0] n23631;
wire            n23632;
wire      [7:0] n23633;
wire            n23634;
wire      [7:0] n23635;
wire            n23636;
wire      [7:0] n23637;
wire            n23638;
wire      [7:0] n23639;
wire      [7:0] n2364;
wire            n23640;
wire      [7:0] n23641;
wire            n23642;
wire      [7:0] n23643;
wire            n23644;
wire      [7:0] n23645;
wire            n23646;
wire      [7:0] n23647;
wire            n23648;
wire      [7:0] n23649;
wire      [7:0] n2365;
wire            n23650;
wire      [7:0] n23651;
wire            n23652;
wire      [7:0] n23653;
wire            n23654;
wire      [7:0] n23655;
wire            n23656;
wire      [7:0] n23657;
wire            n23658;
wire      [7:0] n23659;
wire      [7:0] n2366;
wire            n23660;
wire      [7:0] n23661;
wire            n23662;
wire      [7:0] n23663;
wire            n23664;
wire      [7:0] n23665;
wire            n23666;
wire      [7:0] n23667;
wire            n23668;
wire      [7:0] n23669;
wire      [7:0] n2367;
wire            n23670;
wire      [7:0] n23671;
wire            n23672;
wire      [7:0] n23673;
wire            n23674;
wire      [7:0] n23675;
wire            n23676;
wire      [7:0] n23677;
wire            n23678;
wire      [7:0] n23679;
wire      [7:0] n2368;
wire            n23680;
wire      [7:0] n23681;
wire            n23682;
wire      [7:0] n23683;
wire            n23684;
wire      [7:0] n23685;
wire            n23686;
wire      [7:0] n23687;
wire            n23688;
wire      [7:0] n23689;
wire      [7:0] n2369;
wire            n23690;
wire      [7:0] n23691;
wire            n23692;
wire      [7:0] n23693;
wire            n23694;
wire      [7:0] n23695;
wire            n23696;
wire      [7:0] n23697;
wire            n23698;
wire      [7:0] n23699;
wire      [7:0] n2370;
wire            n23700;
wire      [7:0] n23701;
wire            n23702;
wire      [7:0] n23703;
wire            n23704;
wire      [7:0] n23705;
wire            n23706;
wire      [7:0] n23707;
wire            n23708;
wire      [7:0] n23709;
wire      [7:0] n2371;
wire            n23710;
wire      [7:0] n23711;
wire            n23712;
wire      [7:0] n23713;
wire            n23714;
wire      [7:0] n23715;
wire            n23716;
wire      [7:0] n23717;
wire            n23718;
wire      [7:0] n23719;
wire      [7:0] n2372;
wire            n23720;
wire      [7:0] n23721;
wire            n23722;
wire      [7:0] n23723;
wire            n23724;
wire      [7:0] n23725;
wire            n23726;
wire      [7:0] n23727;
wire            n23728;
wire      [7:0] n23729;
wire      [7:0] n2373;
wire            n23730;
wire      [7:0] n23731;
wire            n23732;
wire      [7:0] n23733;
wire            n23734;
wire      [7:0] n23735;
wire            n23736;
wire      [7:0] n23737;
wire            n23738;
wire      [7:0] n23739;
wire      [7:0] n2374;
wire            n23740;
wire      [7:0] n23741;
wire            n23742;
wire      [7:0] n23743;
wire            n23744;
wire      [7:0] n23745;
wire            n23746;
wire      [7:0] n23747;
wire            n23748;
wire      [7:0] n23749;
wire      [7:0] n2375;
wire            n23750;
wire      [7:0] n23751;
wire            n23752;
wire      [7:0] n23753;
wire            n23754;
wire      [7:0] n23755;
wire            n23756;
wire      [7:0] n23757;
wire            n23758;
wire      [7:0] n23759;
wire      [7:0] n2376;
wire            n23760;
wire      [7:0] n23761;
wire            n23762;
wire      [7:0] n23763;
wire            n23764;
wire      [7:0] n23765;
wire            n23766;
wire      [7:0] n23767;
wire            n23768;
wire      [7:0] n23769;
wire      [7:0] n2377;
wire            n23770;
wire      [7:0] n23771;
wire            n23772;
wire      [7:0] n23773;
wire            n23774;
wire      [7:0] n23775;
wire            n23776;
wire      [7:0] n23777;
wire            n23778;
wire      [7:0] n23779;
wire      [7:0] n2378;
wire            n23780;
wire      [7:0] n23781;
wire            n23782;
wire      [7:0] n23783;
wire            n23784;
wire      [7:0] n23785;
wire            n23786;
wire      [7:0] n23787;
wire            n23788;
wire      [7:0] n23789;
wire      [7:0] n2379;
wire            n23790;
wire      [7:0] n23791;
wire            n23792;
wire      [7:0] n23793;
wire            n23794;
wire      [7:0] n23795;
wire            n23796;
wire      [7:0] n23797;
wire            n23798;
wire      [7:0] n23799;
wire      [7:0] n238;
wire      [7:0] n2380;
wire            n23800;
wire      [7:0] n23801;
wire            n23802;
wire      [7:0] n23803;
wire            n23804;
wire      [7:0] n23805;
wire            n23806;
wire      [7:0] n23807;
wire            n23808;
wire      [7:0] n23809;
wire      [7:0] n2381;
wire            n23810;
wire      [7:0] n23811;
wire            n23812;
wire      [7:0] n23813;
wire            n23814;
wire      [7:0] n23815;
wire            n23816;
wire      [7:0] n23817;
wire            n23818;
wire      [7:0] n23819;
wire      [7:0] n2382;
wire            n23820;
wire      [7:0] n23821;
wire            n23822;
wire      [7:0] n23823;
wire            n23824;
wire      [7:0] n23825;
wire            n23826;
wire      [7:0] n23827;
wire            n23828;
wire      [7:0] n23829;
wire      [7:0] n2383;
wire            n23830;
wire      [7:0] n23831;
wire            n23832;
wire      [7:0] n23833;
wire            n23834;
wire      [7:0] n23835;
wire            n23836;
wire      [7:0] n23837;
wire            n23838;
wire      [7:0] n23839;
wire      [7:0] n2384;
wire            n23840;
wire      [7:0] n23841;
wire            n23842;
wire      [7:0] n23843;
wire            n23844;
wire      [7:0] n23845;
wire            n23846;
wire      [7:0] n23847;
wire            n23848;
wire      [7:0] n23849;
wire      [7:0] n2385;
wire            n23850;
wire      [7:0] n23851;
wire            n23852;
wire      [7:0] n23853;
wire            n23854;
wire      [7:0] n23855;
wire            n23856;
wire      [7:0] n23857;
wire            n23858;
wire      [7:0] n23859;
wire      [7:0] n2386;
wire            n23860;
wire      [7:0] n23861;
wire            n23862;
wire      [7:0] n23863;
wire            n23864;
wire      [7:0] n23865;
wire            n23866;
wire      [7:0] n23867;
wire            n23868;
wire      [7:0] n23869;
wire      [7:0] n2387;
wire            n23870;
wire      [7:0] n23871;
wire            n23872;
wire      [7:0] n23873;
wire            n23874;
wire      [7:0] n23875;
wire            n23876;
wire      [7:0] n23877;
wire            n23878;
wire      [7:0] n23879;
wire      [7:0] n2388;
wire            n23880;
wire      [7:0] n23881;
wire            n23882;
wire      [7:0] n23883;
wire            n23884;
wire      [7:0] n23885;
wire            n23886;
wire      [7:0] n23887;
wire            n23888;
wire      [7:0] n23889;
wire      [7:0] n2389;
wire            n23890;
wire      [7:0] n23891;
wire            n23892;
wire      [7:0] n23893;
wire            n23894;
wire      [7:0] n23895;
wire            n23896;
wire      [7:0] n23897;
wire            n23898;
wire      [7:0] n23899;
wire      [7:0] n2390;
wire            n23900;
wire      [7:0] n23901;
wire            n23902;
wire      [7:0] n23903;
wire      [7:0] n23904;
wire      [7:0] n23905;
wire      [7:0] n23906;
wire      [7:0] n23907;
wire      [7:0] n23908;
wire      [7:0] n23909;
wire      [7:0] n2391;
wire      [7:0] n23910;
wire      [7:0] n23911;
wire      [7:0] n23912;
wire      [7:0] n23913;
wire      [7:0] n23914;
wire      [7:0] n23915;
wire      [7:0] n23916;
wire      [7:0] n23917;
wire      [7:0] n23918;
wire      [7:0] n23919;
wire      [7:0] n2392;
wire      [7:0] n23920;
wire      [7:0] n23921;
wire      [7:0] n23922;
wire      [7:0] n23923;
wire      [7:0] n23924;
wire      [7:0] n23925;
wire      [7:0] n23926;
wire      [7:0] n23927;
wire      [7:0] n23928;
wire      [7:0] n23929;
wire      [7:0] n2393;
wire      [7:0] n23930;
wire      [7:0] n23931;
wire      [7:0] n23932;
wire      [7:0] n23933;
wire      [7:0] n23934;
wire      [7:0] n23935;
wire      [7:0] n23936;
wire      [7:0] n23937;
wire      [7:0] n23938;
wire      [7:0] n23939;
wire      [7:0] n2394;
wire      [7:0] n23940;
wire      [7:0] n23941;
wire      [7:0] n23942;
wire      [7:0] n23943;
wire      [7:0] n23944;
wire      [7:0] n23945;
wire      [7:0] n23946;
wire      [7:0] n23947;
wire      [7:0] n23948;
wire      [7:0] n23949;
wire      [7:0] n2395;
wire      [7:0] n23950;
wire      [7:0] n23951;
wire      [7:0] n23952;
wire      [7:0] n23953;
wire      [7:0] n23954;
wire      [7:0] n23955;
wire      [7:0] n23956;
wire      [7:0] n23957;
wire      [7:0] n23958;
wire      [7:0] n23959;
wire      [7:0] n2396;
wire      [7:0] n23960;
wire      [7:0] n23961;
wire      [7:0] n23962;
wire      [7:0] n23963;
wire      [7:0] n23964;
wire      [7:0] n23965;
wire      [7:0] n23966;
wire      [7:0] n23967;
wire      [7:0] n23968;
wire      [7:0] n23969;
wire      [7:0] n2397;
wire      [7:0] n23970;
wire      [7:0] n23971;
wire      [7:0] n23972;
wire      [7:0] n23973;
wire      [7:0] n23974;
wire      [7:0] n23975;
wire      [7:0] n23976;
wire      [7:0] n23977;
wire      [7:0] n23978;
wire      [7:0] n23979;
wire      [7:0] n2398;
wire      [7:0] n23980;
wire      [7:0] n23981;
wire      [7:0] n23982;
wire      [7:0] n23983;
wire      [7:0] n23984;
wire      [7:0] n23985;
wire      [7:0] n23986;
wire      [7:0] n23987;
wire      [7:0] n23988;
wire      [7:0] n23989;
wire      [7:0] n2399;
wire      [7:0] n23990;
wire      [7:0] n23991;
wire      [7:0] n23992;
wire      [7:0] n23993;
wire      [7:0] n23994;
wire      [7:0] n23995;
wire      [7:0] n23996;
wire      [7:0] n23997;
wire      [7:0] n23998;
wire      [7:0] n23999;
wire            n24;
wire            n240;
wire      [7:0] n2400;
wire      [7:0] n24000;
wire      [7:0] n24001;
wire      [7:0] n24002;
wire      [7:0] n24003;
wire      [7:0] n24004;
wire      [7:0] n24005;
wire      [7:0] n24006;
wire      [7:0] n24007;
wire      [7:0] n24008;
wire      [7:0] n24009;
wire      [7:0] n2401;
wire      [7:0] n24010;
wire      [7:0] n24011;
wire      [7:0] n24012;
wire      [7:0] n24013;
wire      [7:0] n24014;
wire      [7:0] n24015;
wire      [7:0] n24016;
wire      [7:0] n24017;
wire      [7:0] n24018;
wire      [7:0] n24019;
wire      [7:0] n2402;
wire      [7:0] n24020;
wire      [7:0] n24021;
wire      [7:0] n24022;
wire      [7:0] n24023;
wire      [7:0] n24024;
wire      [7:0] n24025;
wire      [7:0] n24026;
wire      [7:0] n24027;
wire      [7:0] n24028;
wire      [7:0] n24029;
wire      [7:0] n2403;
wire      [7:0] n24030;
wire      [7:0] n24031;
wire      [7:0] n24032;
wire      [7:0] n24033;
wire      [7:0] n24034;
wire      [7:0] n24035;
wire      [7:0] n24036;
wire      [7:0] n24037;
wire      [7:0] n24038;
wire      [7:0] n24039;
wire      [7:0] n2404;
wire      [7:0] n24040;
wire      [7:0] n24041;
wire      [7:0] n24042;
wire      [7:0] n24043;
wire      [7:0] n24044;
wire      [7:0] n24045;
wire      [7:0] n24046;
wire      [7:0] n24047;
wire      [7:0] n24048;
wire      [7:0] n24049;
wire      [7:0] n2405;
wire      [7:0] n24050;
wire      [7:0] n24051;
wire      [7:0] n24052;
wire      [7:0] n24053;
wire      [7:0] n24054;
wire      [7:0] n24055;
wire      [7:0] n24056;
wire      [7:0] n24057;
wire      [7:0] n24058;
wire      [7:0] n24059;
wire      [7:0] n2406;
wire      [7:0] n24060;
wire      [7:0] n24061;
wire      [7:0] n24062;
wire      [7:0] n24063;
wire      [7:0] n24064;
wire      [7:0] n24065;
wire      [7:0] n24066;
wire      [7:0] n24067;
wire      [7:0] n24068;
wire      [7:0] n24069;
wire      [7:0] n2407;
wire      [7:0] n24070;
wire      [7:0] n24071;
wire      [7:0] n24072;
wire      [7:0] n24073;
wire      [7:0] n24074;
wire      [7:0] n24075;
wire      [7:0] n24076;
wire      [7:0] n24077;
wire      [7:0] n24078;
wire      [7:0] n24079;
wire      [7:0] n2408;
wire      [7:0] n24080;
wire      [7:0] n24081;
wire      [7:0] n24082;
wire      [7:0] n24083;
wire      [7:0] n24084;
wire      [7:0] n24085;
wire      [7:0] n24086;
wire      [7:0] n24087;
wire      [7:0] n24088;
wire      [7:0] n24089;
wire      [7:0] n2409;
wire      [7:0] n24090;
wire      [7:0] n24091;
wire      [7:0] n24092;
wire      [7:0] n24093;
wire      [7:0] n24094;
wire      [7:0] n24095;
wire      [7:0] n24096;
wire      [7:0] n24097;
wire      [7:0] n24098;
wire      [7:0] n24099;
wire      [7:0] n241;
wire      [7:0] n2410;
wire      [7:0] n24100;
wire      [7:0] n24101;
wire      [7:0] n24102;
wire      [7:0] n24103;
wire      [7:0] n24104;
wire      [7:0] n24105;
wire      [7:0] n24106;
wire      [7:0] n24107;
wire      [7:0] n24108;
wire      [7:0] n24109;
wire      [7:0] n2411;
wire      [7:0] n24110;
wire      [7:0] n24111;
wire      [7:0] n24112;
wire      [7:0] n24113;
wire      [7:0] n24114;
wire      [7:0] n24115;
wire      [7:0] n24116;
wire      [7:0] n24117;
wire      [7:0] n24118;
wire      [7:0] n24119;
wire      [7:0] n2412;
wire      [7:0] n24120;
wire      [7:0] n24121;
wire      [7:0] n24122;
wire      [7:0] n24123;
wire      [7:0] n24124;
wire      [7:0] n24125;
wire      [7:0] n24126;
wire      [7:0] n24127;
wire      [7:0] n24128;
wire      [7:0] n24129;
wire      [7:0] n2413;
wire      [7:0] n24130;
wire      [7:0] n24131;
wire      [7:0] n24132;
wire      [7:0] n24133;
wire      [7:0] n24134;
wire      [7:0] n24135;
wire      [7:0] n24136;
wire      [7:0] n24137;
wire      [7:0] n24138;
wire      [7:0] n24139;
wire      [7:0] n2414;
wire      [7:0] n24140;
wire      [7:0] n24141;
wire      [7:0] n24142;
wire      [7:0] n24143;
wire      [7:0] n24144;
wire      [7:0] n24145;
wire      [7:0] n24146;
wire      [7:0] n24147;
wire      [7:0] n24148;
wire      [7:0] n24149;
wire      [7:0] n2415;
wire      [7:0] n24150;
wire      [7:0] n24151;
wire      [7:0] n24152;
wire      [7:0] n24153;
wire      [7:0] n24154;
wire      [7:0] n24155;
wire      [7:0] n24156;
wire      [7:0] n24157;
wire      [7:0] n24158;
wire      [7:0] n24159;
wire      [7:0] n2416;
wire      [7:0] n24160;
wire      [7:0] n24161;
wire    [111:0] n24162;
wire      [7:0] n24163;
wire      [7:0] n24164;
wire      [7:0] n24165;
wire            n24166;
wire      [7:0] n24167;
wire            n24168;
wire      [7:0] n24169;
wire      [7:0] n2417;
wire            n24170;
wire      [7:0] n24171;
wire            n24172;
wire      [7:0] n24173;
wire            n24174;
wire      [7:0] n24175;
wire            n24176;
wire      [7:0] n24177;
wire            n24178;
wire      [7:0] n24179;
wire      [7:0] n2418;
wire            n24180;
wire      [7:0] n24181;
wire            n24182;
wire      [7:0] n24183;
wire            n24184;
wire      [7:0] n24185;
wire            n24186;
wire      [7:0] n24187;
wire            n24188;
wire      [7:0] n24189;
wire      [7:0] n2419;
wire            n24190;
wire      [7:0] n24191;
wire            n24192;
wire      [7:0] n24193;
wire            n24194;
wire      [7:0] n24195;
wire            n24196;
wire      [7:0] n24197;
wire            n24198;
wire      [7:0] n24199;
wire      [7:0] n2420;
wire            n24200;
wire      [7:0] n24201;
wire            n24202;
wire      [7:0] n24203;
wire            n24204;
wire      [7:0] n24205;
wire            n24206;
wire      [7:0] n24207;
wire            n24208;
wire      [7:0] n24209;
wire      [7:0] n2421;
wire            n24210;
wire      [7:0] n24211;
wire            n24212;
wire      [7:0] n24213;
wire            n24214;
wire      [7:0] n24215;
wire            n24216;
wire      [7:0] n24217;
wire            n24218;
wire      [7:0] n24219;
wire      [7:0] n2422;
wire            n24220;
wire      [7:0] n24221;
wire            n24222;
wire      [7:0] n24223;
wire            n24224;
wire      [7:0] n24225;
wire            n24226;
wire      [7:0] n24227;
wire            n24228;
wire      [7:0] n24229;
wire      [7:0] n2423;
wire            n24230;
wire      [7:0] n24231;
wire            n24232;
wire      [7:0] n24233;
wire            n24234;
wire      [7:0] n24235;
wire            n24236;
wire      [7:0] n24237;
wire            n24238;
wire      [7:0] n24239;
wire      [7:0] n2424;
wire            n24240;
wire      [7:0] n24241;
wire            n24242;
wire      [7:0] n24243;
wire            n24244;
wire      [7:0] n24245;
wire            n24246;
wire      [7:0] n24247;
wire            n24248;
wire      [7:0] n24249;
wire      [7:0] n2425;
wire            n24250;
wire      [7:0] n24251;
wire            n24252;
wire      [7:0] n24253;
wire            n24254;
wire      [7:0] n24255;
wire            n24256;
wire      [7:0] n24257;
wire            n24258;
wire      [7:0] n24259;
wire      [7:0] n2426;
wire            n24260;
wire      [7:0] n24261;
wire            n24262;
wire      [7:0] n24263;
wire            n24264;
wire      [7:0] n24265;
wire            n24266;
wire      [7:0] n24267;
wire            n24268;
wire      [7:0] n24269;
wire      [7:0] n2427;
wire            n24270;
wire      [7:0] n24271;
wire            n24272;
wire      [7:0] n24273;
wire            n24274;
wire      [7:0] n24275;
wire            n24276;
wire      [7:0] n24277;
wire            n24278;
wire      [7:0] n24279;
wire      [7:0] n2428;
wire            n24280;
wire      [7:0] n24281;
wire            n24282;
wire      [7:0] n24283;
wire            n24284;
wire      [7:0] n24285;
wire            n24286;
wire      [7:0] n24287;
wire            n24288;
wire      [7:0] n24289;
wire      [7:0] n2429;
wire            n24290;
wire      [7:0] n24291;
wire            n24292;
wire      [7:0] n24293;
wire            n24294;
wire      [7:0] n24295;
wire            n24296;
wire      [7:0] n24297;
wire            n24298;
wire      [7:0] n24299;
wire            n243;
wire      [7:0] n2430;
wire            n24300;
wire      [7:0] n24301;
wire            n24302;
wire      [7:0] n24303;
wire            n24304;
wire      [7:0] n24305;
wire            n24306;
wire      [7:0] n24307;
wire            n24308;
wire      [7:0] n24309;
wire      [7:0] n2431;
wire            n24310;
wire      [7:0] n24311;
wire            n24312;
wire      [7:0] n24313;
wire            n24314;
wire      [7:0] n24315;
wire            n24316;
wire      [7:0] n24317;
wire            n24318;
wire      [7:0] n24319;
wire      [7:0] n2432;
wire            n24320;
wire      [7:0] n24321;
wire            n24322;
wire      [7:0] n24323;
wire            n24324;
wire      [7:0] n24325;
wire            n24326;
wire      [7:0] n24327;
wire            n24328;
wire      [7:0] n24329;
wire      [7:0] n2433;
wire            n24330;
wire      [7:0] n24331;
wire            n24332;
wire      [7:0] n24333;
wire            n24334;
wire      [7:0] n24335;
wire            n24336;
wire      [7:0] n24337;
wire            n24338;
wire      [7:0] n24339;
wire      [7:0] n2434;
wire            n24340;
wire      [7:0] n24341;
wire            n24342;
wire      [7:0] n24343;
wire            n24344;
wire      [7:0] n24345;
wire            n24346;
wire      [7:0] n24347;
wire            n24348;
wire      [7:0] n24349;
wire      [7:0] n2435;
wire            n24350;
wire      [7:0] n24351;
wire            n24352;
wire      [7:0] n24353;
wire            n24354;
wire      [7:0] n24355;
wire            n24356;
wire      [7:0] n24357;
wire            n24358;
wire      [7:0] n24359;
wire      [7:0] n2436;
wire            n24360;
wire      [7:0] n24361;
wire            n24362;
wire      [7:0] n24363;
wire            n24364;
wire      [7:0] n24365;
wire            n24366;
wire      [7:0] n24367;
wire            n24368;
wire      [7:0] n24369;
wire      [7:0] n2437;
wire            n24370;
wire      [7:0] n24371;
wire            n24372;
wire      [7:0] n24373;
wire            n24374;
wire      [7:0] n24375;
wire            n24376;
wire      [7:0] n24377;
wire            n24378;
wire      [7:0] n24379;
wire      [7:0] n2438;
wire            n24380;
wire      [7:0] n24381;
wire            n24382;
wire      [7:0] n24383;
wire            n24384;
wire      [7:0] n24385;
wire            n24386;
wire      [7:0] n24387;
wire            n24388;
wire      [7:0] n24389;
wire      [7:0] n2439;
wire            n24390;
wire      [7:0] n24391;
wire            n24392;
wire      [7:0] n24393;
wire            n24394;
wire      [7:0] n24395;
wire            n24396;
wire      [7:0] n24397;
wire            n24398;
wire      [7:0] n24399;
wire      [7:0] n2440;
wire            n24400;
wire      [7:0] n24401;
wire            n24402;
wire      [7:0] n24403;
wire            n24404;
wire      [7:0] n24405;
wire            n24406;
wire      [7:0] n24407;
wire            n24408;
wire      [7:0] n24409;
wire      [7:0] n2441;
wire            n24410;
wire      [7:0] n24411;
wire            n24412;
wire      [7:0] n24413;
wire            n24414;
wire      [7:0] n24415;
wire            n24416;
wire      [7:0] n24417;
wire            n24418;
wire      [7:0] n24419;
wire      [7:0] n2442;
wire            n24420;
wire      [7:0] n24421;
wire            n24422;
wire      [7:0] n24423;
wire            n24424;
wire      [7:0] n24425;
wire            n24426;
wire      [7:0] n24427;
wire            n24428;
wire      [7:0] n24429;
wire      [7:0] n2443;
wire            n24430;
wire      [7:0] n24431;
wire            n24432;
wire      [7:0] n24433;
wire            n24434;
wire      [7:0] n24435;
wire            n24436;
wire      [7:0] n24437;
wire            n24438;
wire      [7:0] n24439;
wire      [7:0] n2444;
wire            n24440;
wire      [7:0] n24441;
wire            n24442;
wire      [7:0] n24443;
wire            n24444;
wire      [7:0] n24445;
wire            n24446;
wire      [7:0] n24447;
wire            n24448;
wire      [7:0] n24449;
wire      [7:0] n2445;
wire            n24450;
wire      [7:0] n24451;
wire            n24452;
wire      [7:0] n24453;
wire            n24454;
wire      [7:0] n24455;
wire            n24456;
wire      [7:0] n24457;
wire            n24458;
wire      [7:0] n24459;
wire      [7:0] n2446;
wire            n24460;
wire      [7:0] n24461;
wire            n24462;
wire      [7:0] n24463;
wire            n24464;
wire      [7:0] n24465;
wire            n24466;
wire      [7:0] n24467;
wire            n24468;
wire      [7:0] n24469;
wire      [7:0] n2447;
wire            n24470;
wire      [7:0] n24471;
wire            n24472;
wire      [7:0] n24473;
wire            n24474;
wire      [7:0] n24475;
wire            n24476;
wire      [7:0] n24477;
wire            n24478;
wire      [7:0] n24479;
wire      [7:0] n2448;
wire            n24480;
wire      [7:0] n24481;
wire            n24482;
wire      [7:0] n24483;
wire            n24484;
wire      [7:0] n24485;
wire            n24486;
wire      [7:0] n24487;
wire            n24488;
wire      [7:0] n24489;
wire      [7:0] n2449;
wire            n24490;
wire      [7:0] n24491;
wire            n24492;
wire      [7:0] n24493;
wire            n24494;
wire      [7:0] n24495;
wire            n24496;
wire      [7:0] n24497;
wire            n24498;
wire      [7:0] n24499;
wire      [7:0] n245;
wire      [7:0] n2450;
wire            n24500;
wire      [7:0] n24501;
wire            n24502;
wire      [7:0] n24503;
wire            n24504;
wire      [7:0] n24505;
wire            n24506;
wire      [7:0] n24507;
wire            n24508;
wire      [7:0] n24509;
wire      [7:0] n2451;
wire            n24510;
wire      [7:0] n24511;
wire            n24512;
wire      [7:0] n24513;
wire            n24514;
wire      [7:0] n24515;
wire            n24516;
wire      [7:0] n24517;
wire            n24518;
wire      [7:0] n24519;
wire      [7:0] n2452;
wire            n24520;
wire      [7:0] n24521;
wire            n24522;
wire      [7:0] n24523;
wire            n24524;
wire      [7:0] n24525;
wire            n24526;
wire      [7:0] n24527;
wire            n24528;
wire      [7:0] n24529;
wire      [7:0] n2453;
wire            n24530;
wire      [7:0] n24531;
wire            n24532;
wire      [7:0] n24533;
wire            n24534;
wire      [7:0] n24535;
wire            n24536;
wire      [7:0] n24537;
wire            n24538;
wire      [7:0] n24539;
wire      [7:0] n2454;
wire            n24540;
wire      [7:0] n24541;
wire            n24542;
wire      [7:0] n24543;
wire            n24544;
wire      [7:0] n24545;
wire            n24546;
wire      [7:0] n24547;
wire            n24548;
wire      [7:0] n24549;
wire      [7:0] n2455;
wire            n24550;
wire      [7:0] n24551;
wire            n24552;
wire      [7:0] n24553;
wire            n24554;
wire      [7:0] n24555;
wire            n24556;
wire      [7:0] n24557;
wire            n24558;
wire      [7:0] n24559;
wire      [7:0] n2456;
wire            n24560;
wire      [7:0] n24561;
wire            n24562;
wire      [7:0] n24563;
wire            n24564;
wire      [7:0] n24565;
wire            n24566;
wire      [7:0] n24567;
wire            n24568;
wire      [7:0] n24569;
wire      [7:0] n2457;
wire            n24570;
wire      [7:0] n24571;
wire            n24572;
wire      [7:0] n24573;
wire            n24574;
wire      [7:0] n24575;
wire            n24576;
wire      [7:0] n24577;
wire            n24578;
wire      [7:0] n24579;
wire      [7:0] n2458;
wire            n24580;
wire      [7:0] n24581;
wire            n24582;
wire      [7:0] n24583;
wire            n24584;
wire      [7:0] n24585;
wire            n24586;
wire      [7:0] n24587;
wire            n24588;
wire      [7:0] n24589;
wire      [7:0] n2459;
wire            n24590;
wire      [7:0] n24591;
wire            n24592;
wire      [7:0] n24593;
wire            n24594;
wire      [7:0] n24595;
wire            n24596;
wire      [7:0] n24597;
wire            n24598;
wire      [7:0] n24599;
wire      [7:0] n2460;
wire            n24600;
wire      [7:0] n24601;
wire            n24602;
wire      [7:0] n24603;
wire            n24604;
wire      [7:0] n24605;
wire            n24606;
wire      [7:0] n24607;
wire            n24608;
wire      [7:0] n24609;
wire      [7:0] n2461;
wire            n24610;
wire      [7:0] n24611;
wire            n24612;
wire      [7:0] n24613;
wire            n24614;
wire      [7:0] n24615;
wire            n24616;
wire      [7:0] n24617;
wire            n24618;
wire      [7:0] n24619;
wire      [7:0] n2462;
wire            n24620;
wire      [7:0] n24621;
wire            n24622;
wire      [7:0] n24623;
wire            n24624;
wire      [7:0] n24625;
wire            n24626;
wire      [7:0] n24627;
wire            n24628;
wire      [7:0] n24629;
wire      [7:0] n2463;
wire            n24630;
wire      [7:0] n24631;
wire            n24632;
wire      [7:0] n24633;
wire            n24634;
wire      [7:0] n24635;
wire            n24636;
wire      [7:0] n24637;
wire            n24638;
wire      [7:0] n24639;
wire      [7:0] n2464;
wire            n24640;
wire      [7:0] n24641;
wire            n24642;
wire      [7:0] n24643;
wire            n24644;
wire      [7:0] n24645;
wire            n24646;
wire      [7:0] n24647;
wire            n24648;
wire      [7:0] n24649;
wire      [7:0] n2465;
wire            n24650;
wire      [7:0] n24651;
wire            n24652;
wire      [7:0] n24653;
wire            n24654;
wire      [7:0] n24655;
wire            n24656;
wire      [7:0] n24657;
wire            n24658;
wire      [7:0] n24659;
wire      [7:0] n2466;
wire            n24660;
wire      [7:0] n24661;
wire            n24662;
wire      [7:0] n24663;
wire            n24664;
wire      [7:0] n24665;
wire            n24666;
wire      [7:0] n24667;
wire            n24668;
wire      [7:0] n24669;
wire      [7:0] n2467;
wire            n24670;
wire      [7:0] n24671;
wire            n24672;
wire      [7:0] n24673;
wire            n24674;
wire      [7:0] n24675;
wire            n24676;
wire      [7:0] n24677;
wire      [7:0] n24678;
wire      [7:0] n24679;
wire      [7:0] n2468;
wire      [7:0] n24680;
wire      [7:0] n24681;
wire      [7:0] n24682;
wire      [7:0] n24683;
wire      [7:0] n24684;
wire      [7:0] n24685;
wire      [7:0] n24686;
wire      [7:0] n24687;
wire      [7:0] n24688;
wire      [7:0] n24689;
wire      [7:0] n2469;
wire      [7:0] n24690;
wire      [7:0] n24691;
wire      [7:0] n24692;
wire      [7:0] n24693;
wire      [7:0] n24694;
wire      [7:0] n24695;
wire      [7:0] n24696;
wire      [7:0] n24697;
wire      [7:0] n24698;
wire      [7:0] n24699;
wire            n247;
wire      [7:0] n2470;
wire      [7:0] n24700;
wire      [7:0] n24701;
wire      [7:0] n24702;
wire      [7:0] n24703;
wire      [7:0] n24704;
wire      [7:0] n24705;
wire      [7:0] n24706;
wire      [7:0] n24707;
wire      [7:0] n24708;
wire      [7:0] n24709;
wire      [7:0] n2471;
wire      [7:0] n24710;
wire      [7:0] n24711;
wire      [7:0] n24712;
wire      [7:0] n24713;
wire      [7:0] n24714;
wire      [7:0] n24715;
wire      [7:0] n24716;
wire      [7:0] n24717;
wire      [7:0] n24718;
wire      [7:0] n24719;
wire      [7:0] n2472;
wire      [7:0] n24720;
wire      [7:0] n24721;
wire      [7:0] n24722;
wire      [7:0] n24723;
wire      [7:0] n24724;
wire      [7:0] n24725;
wire      [7:0] n24726;
wire      [7:0] n24727;
wire      [7:0] n24728;
wire      [7:0] n24729;
wire      [7:0] n2473;
wire      [7:0] n24730;
wire      [7:0] n24731;
wire      [7:0] n24732;
wire      [7:0] n24733;
wire      [7:0] n24734;
wire      [7:0] n24735;
wire      [7:0] n24736;
wire      [7:0] n24737;
wire      [7:0] n24738;
wire      [7:0] n24739;
wire      [7:0] n2474;
wire      [7:0] n24740;
wire      [7:0] n24741;
wire      [7:0] n24742;
wire      [7:0] n24743;
wire      [7:0] n24744;
wire      [7:0] n24745;
wire      [7:0] n24746;
wire      [7:0] n24747;
wire      [7:0] n24748;
wire      [7:0] n24749;
wire      [7:0] n2475;
wire      [7:0] n24750;
wire      [7:0] n24751;
wire      [7:0] n24752;
wire      [7:0] n24753;
wire      [7:0] n24754;
wire      [7:0] n24755;
wire      [7:0] n24756;
wire      [7:0] n24757;
wire      [7:0] n24758;
wire      [7:0] n24759;
wire      [7:0] n2476;
wire      [7:0] n24760;
wire      [7:0] n24761;
wire      [7:0] n24762;
wire      [7:0] n24763;
wire      [7:0] n24764;
wire      [7:0] n24765;
wire      [7:0] n24766;
wire      [7:0] n24767;
wire      [7:0] n24768;
wire      [7:0] n24769;
wire      [7:0] n2477;
wire      [7:0] n24770;
wire      [7:0] n24771;
wire      [7:0] n24772;
wire      [7:0] n24773;
wire      [7:0] n24774;
wire      [7:0] n24775;
wire      [7:0] n24776;
wire      [7:0] n24777;
wire      [7:0] n24778;
wire      [7:0] n24779;
wire      [7:0] n2478;
wire      [7:0] n24780;
wire      [7:0] n24781;
wire      [7:0] n24782;
wire      [7:0] n24783;
wire      [7:0] n24784;
wire      [7:0] n24785;
wire      [7:0] n24786;
wire      [7:0] n24787;
wire      [7:0] n24788;
wire      [7:0] n24789;
wire      [7:0] n2479;
wire      [7:0] n24790;
wire      [7:0] n24791;
wire      [7:0] n24792;
wire      [7:0] n24793;
wire      [7:0] n24794;
wire      [7:0] n24795;
wire      [7:0] n24796;
wire      [7:0] n24797;
wire      [7:0] n24798;
wire      [7:0] n24799;
wire      [7:0] n2480;
wire      [7:0] n24800;
wire      [7:0] n24801;
wire      [7:0] n24802;
wire      [7:0] n24803;
wire      [7:0] n24804;
wire      [7:0] n24805;
wire      [7:0] n24806;
wire      [7:0] n24807;
wire      [7:0] n24808;
wire      [7:0] n24809;
wire      [7:0] n2481;
wire      [7:0] n24810;
wire      [7:0] n24811;
wire      [7:0] n24812;
wire      [7:0] n24813;
wire      [7:0] n24814;
wire      [7:0] n24815;
wire      [7:0] n24816;
wire      [7:0] n24817;
wire      [7:0] n24818;
wire      [7:0] n24819;
wire      [7:0] n2482;
wire      [7:0] n24820;
wire      [7:0] n24821;
wire      [7:0] n24822;
wire      [7:0] n24823;
wire      [7:0] n24824;
wire      [7:0] n24825;
wire      [7:0] n24826;
wire      [7:0] n24827;
wire      [7:0] n24828;
wire      [7:0] n24829;
wire      [7:0] n2483;
wire      [7:0] n24830;
wire      [7:0] n24831;
wire      [7:0] n24832;
wire      [7:0] n24833;
wire      [7:0] n24834;
wire      [7:0] n24835;
wire      [7:0] n24836;
wire      [7:0] n24837;
wire      [7:0] n24838;
wire      [7:0] n24839;
wire      [7:0] n2484;
wire      [7:0] n24840;
wire      [7:0] n24841;
wire      [7:0] n24842;
wire      [7:0] n24843;
wire      [7:0] n24844;
wire      [7:0] n24845;
wire      [7:0] n24846;
wire      [7:0] n24847;
wire      [7:0] n24848;
wire      [7:0] n24849;
wire      [7:0] n2485;
wire      [7:0] n24850;
wire      [7:0] n24851;
wire      [7:0] n24852;
wire      [7:0] n24853;
wire      [7:0] n24854;
wire      [7:0] n24855;
wire      [7:0] n24856;
wire      [7:0] n24857;
wire      [7:0] n24858;
wire      [7:0] n24859;
wire      [7:0] n2486;
wire      [7:0] n24860;
wire      [7:0] n24861;
wire      [7:0] n24862;
wire      [7:0] n24863;
wire      [7:0] n24864;
wire      [7:0] n24865;
wire      [7:0] n24866;
wire      [7:0] n24867;
wire      [7:0] n24868;
wire      [7:0] n24869;
wire      [7:0] n2487;
wire      [7:0] n24870;
wire      [7:0] n24871;
wire      [7:0] n24872;
wire      [7:0] n24873;
wire      [7:0] n24874;
wire      [7:0] n24875;
wire      [7:0] n24876;
wire      [7:0] n24877;
wire      [7:0] n24878;
wire      [7:0] n24879;
wire      [7:0] n2488;
wire      [7:0] n24880;
wire      [7:0] n24881;
wire      [7:0] n24882;
wire      [7:0] n24883;
wire      [7:0] n24884;
wire      [7:0] n24885;
wire      [7:0] n24886;
wire      [7:0] n24887;
wire      [7:0] n24888;
wire      [7:0] n24889;
wire      [7:0] n2489;
wire      [7:0] n24890;
wire      [7:0] n24891;
wire      [7:0] n24892;
wire      [7:0] n24893;
wire      [7:0] n24894;
wire      [7:0] n24895;
wire      [7:0] n24896;
wire      [7:0] n24897;
wire      [7:0] n24898;
wire      [7:0] n24899;
wire      [7:0] n249;
wire      [7:0] n2490;
wire      [7:0] n24900;
wire      [7:0] n24901;
wire      [7:0] n24902;
wire      [7:0] n24903;
wire      [7:0] n24904;
wire      [7:0] n24905;
wire      [7:0] n24906;
wire      [7:0] n24907;
wire      [7:0] n24908;
wire      [7:0] n24909;
wire      [7:0] n2491;
wire      [7:0] n24910;
wire      [7:0] n24911;
wire      [7:0] n24912;
wire      [7:0] n24913;
wire      [7:0] n24914;
wire      [7:0] n24915;
wire      [7:0] n24916;
wire      [7:0] n24917;
wire      [7:0] n24918;
wire      [7:0] n24919;
wire      [7:0] n2492;
wire      [7:0] n24920;
wire      [7:0] n24921;
wire      [7:0] n24922;
wire      [7:0] n24923;
wire      [7:0] n24924;
wire      [7:0] n24925;
wire      [7:0] n24926;
wire      [7:0] n24927;
wire      [7:0] n24928;
wire      [7:0] n24929;
wire      [7:0] n2493;
wire      [7:0] n24930;
wire      [7:0] n24931;
wire      [7:0] n24932;
wire      [7:0] n24933;
wire      [7:0] n24934;
wire      [7:0] n24935;
wire      [7:0] n24936;
wire    [119:0] n24937;
wire      [7:0] n24938;
wire      [7:0] n24939;
wire      [7:0] n2494;
wire      [7:0] n24940;
wire      [7:0] n24941;
wire      [7:0] n24942;
wire      [7:0] n24943;
wire    [127:0] n24944;
wire    [127:0] n24945;
wire      [7:0] n2495;
wire      [7:0] n2496;
wire      [7:0] n2497;
wire      [7:0] n2498;
wire      [7:0] n2499;
wire      [7:0] n2500;
wire      [7:0] n2501;
wire      [7:0] n2502;
wire      [7:0] n2503;
wire      [7:0] n2504;
wire      [7:0] n2505;
wire      [7:0] n2506;
wire      [7:0] n2507;
wire      [7:0] n2508;
wire      [7:0] n2509;
wire            n251;
wire      [7:0] n2510;
wire      [7:0] n2511;
wire      [7:0] n2512;
wire      [7:0] n2513;
wire      [7:0] n2514;
wire      [7:0] n2515;
wire      [7:0] n2516;
wire      [7:0] n2517;
wire      [7:0] n2518;
wire      [7:0] n2519;
wire      [7:0] n2520;
wire      [7:0] n2521;
wire      [7:0] n2522;
wire      [7:0] n2523;
wire      [7:0] n2524;
wire      [7:0] n2525;
wire      [7:0] n2526;
wire      [7:0] n2527;
wire      [7:0] n2528;
wire      [7:0] n2529;
wire      [7:0] n253;
wire      [7:0] n2530;
wire      [7:0] n2531;
wire      [7:0] n2532;
wire      [7:0] n2533;
wire      [7:0] n2534;
wire      [7:0] n2535;
wire      [7:0] n2536;
wire      [7:0] n2537;
wire      [7:0] n2538;
wire      [7:0] n2539;
wire      [7:0] n2540;
wire      [7:0] n2541;
wire      [7:0] n2542;
wire      [7:0] n2543;
wire      [7:0] n2544;
wire      [7:0] n2545;
wire      [7:0] n2546;
wire      [7:0] n2547;
wire      [7:0] n2548;
wire      [7:0] n2549;
wire            n255;
wire      [7:0] n2550;
wire      [7:0] n2551;
wire      [7:0] n2552;
wire      [7:0] n2553;
wire      [7:0] n2554;
wire      [7:0] n2555;
wire      [7:0] n2556;
wire      [7:0] n2557;
wire      [7:0] n2558;
wire      [7:0] n2559;
wire      [7:0] n256;
wire      [7:0] n2560;
wire      [7:0] n2561;
wire      [7:0] n2562;
wire      [7:0] n2563;
wire      [7:0] n2564;
wire            n2565;
wire      [7:0] n2566;
wire            n2567;
wire      [7:0] n2568;
wire            n2569;
wire      [7:0] n2570;
wire            n2571;
wire      [7:0] n2572;
wire            n2573;
wire      [7:0] n2574;
wire            n2575;
wire      [7:0] n2576;
wire            n2577;
wire      [7:0] n2578;
wire            n2579;
wire            n258;
wire      [7:0] n2580;
wire            n2581;
wire      [7:0] n2582;
wire            n2583;
wire      [7:0] n2584;
wire            n2585;
wire      [7:0] n2586;
wire            n2587;
wire      [7:0] n2588;
wire            n2589;
wire      [7:0] n259;
wire      [7:0] n2590;
wire            n2591;
wire      [7:0] n2592;
wire            n2593;
wire      [7:0] n2594;
wire            n2595;
wire      [7:0] n2596;
wire            n2597;
wire      [7:0] n2598;
wire            n2599;
wire      [7:0] n26;
wire      [7:0] n2600;
wire            n2601;
wire      [7:0] n2602;
wire            n2603;
wire      [7:0] n2604;
wire            n2605;
wire      [7:0] n2606;
wire            n2607;
wire      [7:0] n2608;
wire            n2609;
wire            n261;
wire      [7:0] n2610;
wire            n2611;
wire      [7:0] n2612;
wire            n2613;
wire      [7:0] n2614;
wire            n2615;
wire      [7:0] n2616;
wire            n2617;
wire      [7:0] n2618;
wire            n2619;
wire      [7:0] n262;
wire      [7:0] n2620;
wire            n2621;
wire      [7:0] n2622;
wire            n2623;
wire      [7:0] n2624;
wire            n2625;
wire      [7:0] n2626;
wire            n2627;
wire      [7:0] n2628;
wire            n2629;
wire      [7:0] n2630;
wire            n2631;
wire      [7:0] n2632;
wire            n2633;
wire      [7:0] n2634;
wire            n2635;
wire      [7:0] n2636;
wire            n2637;
wire      [7:0] n2638;
wire            n2639;
wire            n264;
wire      [7:0] n2640;
wire            n2641;
wire      [7:0] n2642;
wire            n2643;
wire      [7:0] n2644;
wire            n2645;
wire      [7:0] n2646;
wire            n2647;
wire      [7:0] n2648;
wire            n2649;
wire      [7:0] n265;
wire      [7:0] n2650;
wire            n2651;
wire      [7:0] n2652;
wire            n2653;
wire      [7:0] n2654;
wire            n2655;
wire      [7:0] n2656;
wire            n2657;
wire      [7:0] n2658;
wire            n2659;
wire      [7:0] n2660;
wire            n2661;
wire      [7:0] n2662;
wire            n2663;
wire      [7:0] n2664;
wire            n2665;
wire      [7:0] n2666;
wire            n2667;
wire      [7:0] n2668;
wire            n2669;
wire            n267;
wire      [7:0] n2670;
wire            n2671;
wire      [7:0] n2672;
wire            n2673;
wire      [7:0] n2674;
wire            n2675;
wire      [7:0] n2676;
wire            n2677;
wire      [7:0] n2678;
wire            n2679;
wire      [7:0] n2680;
wire            n2681;
wire      [7:0] n2682;
wire            n2683;
wire      [7:0] n2684;
wire            n2685;
wire      [7:0] n2686;
wire            n2687;
wire      [7:0] n2688;
wire            n2689;
wire      [7:0] n269;
wire      [7:0] n2690;
wire            n2691;
wire      [7:0] n2692;
wire            n2693;
wire      [7:0] n2694;
wire            n2695;
wire      [7:0] n2696;
wire            n2697;
wire      [7:0] n2698;
wire            n2699;
wire      [7:0] n2700;
wire            n2701;
wire      [7:0] n2702;
wire            n2703;
wire      [7:0] n2704;
wire            n2705;
wire      [7:0] n2706;
wire            n2707;
wire      [7:0] n2708;
wire            n2709;
wire            n271;
wire      [7:0] n2710;
wire            n2711;
wire      [7:0] n2712;
wire            n2713;
wire      [7:0] n2714;
wire            n2715;
wire      [7:0] n2716;
wire            n2717;
wire      [7:0] n2718;
wire            n2719;
wire      [7:0] n272;
wire      [7:0] n2720;
wire            n2721;
wire      [7:0] n2722;
wire            n2723;
wire      [7:0] n2724;
wire            n2725;
wire      [7:0] n2726;
wire            n2727;
wire      [7:0] n2728;
wire            n2729;
wire      [7:0] n2730;
wire            n2731;
wire      [7:0] n2732;
wire            n2733;
wire      [7:0] n2734;
wire            n2735;
wire      [7:0] n2736;
wire            n2737;
wire      [7:0] n2738;
wire            n2739;
wire            n274;
wire      [7:0] n2740;
wire            n2741;
wire      [7:0] n2742;
wire            n2743;
wire      [7:0] n2744;
wire            n2745;
wire      [7:0] n2746;
wire            n2747;
wire      [7:0] n2748;
wire            n2749;
wire      [7:0] n2750;
wire            n2751;
wire      [7:0] n2752;
wire            n2753;
wire      [7:0] n2754;
wire            n2755;
wire      [7:0] n2756;
wire            n2757;
wire      [7:0] n2758;
wire            n2759;
wire      [7:0] n276;
wire      [7:0] n2760;
wire            n2761;
wire      [7:0] n2762;
wire            n2763;
wire      [7:0] n2764;
wire            n2765;
wire      [7:0] n2766;
wire            n2767;
wire      [7:0] n2768;
wire            n2769;
wire      [7:0] n2770;
wire            n2771;
wire      [7:0] n2772;
wire            n2773;
wire      [7:0] n2774;
wire            n2775;
wire      [7:0] n2776;
wire            n2777;
wire      [7:0] n2778;
wire            n2779;
wire            n278;
wire      [7:0] n2780;
wire            n2781;
wire      [7:0] n2782;
wire            n2783;
wire      [7:0] n2784;
wire            n2785;
wire      [7:0] n2786;
wire            n2787;
wire      [7:0] n2788;
wire            n2789;
wire      [7:0] n2790;
wire            n2791;
wire      [7:0] n2792;
wire            n2793;
wire      [7:0] n2794;
wire            n2795;
wire      [7:0] n2796;
wire            n2797;
wire      [7:0] n2798;
wire            n2799;
wire            n28;
wire      [7:0] n280;
wire      [7:0] n2800;
wire            n2801;
wire      [7:0] n2802;
wire            n2803;
wire      [7:0] n2804;
wire            n2805;
wire      [7:0] n2806;
wire            n2807;
wire      [7:0] n2808;
wire            n2809;
wire      [7:0] n2810;
wire            n2811;
wire      [7:0] n2812;
wire            n2813;
wire      [7:0] n2814;
wire            n2815;
wire      [7:0] n2816;
wire            n2817;
wire      [7:0] n2818;
wire            n2819;
wire            n282;
wire      [7:0] n2820;
wire            n2821;
wire      [7:0] n2822;
wire            n2823;
wire      [7:0] n2824;
wire            n2825;
wire      [7:0] n2826;
wire            n2827;
wire      [7:0] n2828;
wire            n2829;
wire      [7:0] n2830;
wire            n2831;
wire      [7:0] n2832;
wire            n2833;
wire      [7:0] n2834;
wire            n2835;
wire      [7:0] n2836;
wire            n2837;
wire      [7:0] n2838;
wire            n2839;
wire      [7:0] n284;
wire      [7:0] n2840;
wire            n2841;
wire      [7:0] n2842;
wire            n2843;
wire      [7:0] n2844;
wire            n2845;
wire      [7:0] n2846;
wire            n2847;
wire      [7:0] n2848;
wire            n2849;
wire      [7:0] n2850;
wire            n2851;
wire      [7:0] n2852;
wire            n2853;
wire      [7:0] n2854;
wire            n2855;
wire      [7:0] n2856;
wire            n2857;
wire      [7:0] n2858;
wire            n2859;
wire            n286;
wire      [7:0] n2860;
wire            n2861;
wire      [7:0] n2862;
wire            n2863;
wire      [7:0] n2864;
wire            n2865;
wire      [7:0] n2866;
wire            n2867;
wire      [7:0] n2868;
wire            n2869;
wire      [7:0] n2870;
wire            n2871;
wire      [7:0] n2872;
wire            n2873;
wire      [7:0] n2874;
wire            n2875;
wire      [7:0] n2876;
wire            n2877;
wire      [7:0] n2878;
wire            n2879;
wire      [7:0] n288;
wire      [7:0] n2880;
wire            n2881;
wire      [7:0] n2882;
wire            n2883;
wire      [7:0] n2884;
wire            n2885;
wire      [7:0] n2886;
wire            n2887;
wire      [7:0] n2888;
wire            n2889;
wire      [7:0] n2890;
wire            n2891;
wire      [7:0] n2892;
wire            n2893;
wire      [7:0] n2894;
wire            n2895;
wire      [7:0] n2896;
wire            n2897;
wire      [7:0] n2898;
wire            n2899;
wire            n290;
wire      [7:0] n2900;
wire            n2901;
wire      [7:0] n2902;
wire            n2903;
wire      [7:0] n2904;
wire            n2905;
wire      [7:0] n2906;
wire            n2907;
wire      [7:0] n2908;
wire            n2909;
wire      [7:0] n291;
wire      [7:0] n2910;
wire            n2911;
wire      [7:0] n2912;
wire            n2913;
wire      [7:0] n2914;
wire            n2915;
wire      [7:0] n2916;
wire            n2917;
wire      [7:0] n2918;
wire            n2919;
wire      [7:0] n2920;
wire            n2921;
wire      [7:0] n2922;
wire            n2923;
wire      [7:0] n2924;
wire            n2925;
wire      [7:0] n2926;
wire            n2927;
wire      [7:0] n2928;
wire            n2929;
wire            n293;
wire      [7:0] n2930;
wire            n2931;
wire      [7:0] n2932;
wire            n2933;
wire      [7:0] n2934;
wire            n2935;
wire      [7:0] n2936;
wire            n2937;
wire      [7:0] n2938;
wire            n2939;
wire      [7:0] n2940;
wire            n2941;
wire      [7:0] n2942;
wire            n2943;
wire      [7:0] n2944;
wire            n2945;
wire      [7:0] n2946;
wire            n2947;
wire      [7:0] n2948;
wire            n2949;
wire      [7:0] n295;
wire      [7:0] n2950;
wire            n2951;
wire      [7:0] n2952;
wire            n2953;
wire      [7:0] n2954;
wire            n2955;
wire      [7:0] n2956;
wire            n2957;
wire      [7:0] n2958;
wire            n2959;
wire            n296;
wire      [7:0] n2960;
wire            n2961;
wire      [7:0] n2962;
wire            n2963;
wire      [7:0] n2964;
wire            n2965;
wire      [7:0] n2966;
wire            n2967;
wire      [7:0] n2968;
wire            n2969;
wire      [7:0] n2970;
wire            n2971;
wire      [7:0] n2972;
wire            n2973;
wire      [7:0] n2974;
wire            n2975;
wire      [7:0] n2976;
wire            n2977;
wire      [7:0] n2978;
wire            n2979;
wire      [7:0] n298;
wire      [7:0] n2980;
wire            n2981;
wire      [7:0] n2982;
wire            n2983;
wire      [7:0] n2984;
wire            n2985;
wire      [7:0] n2986;
wire            n2987;
wire      [7:0] n2988;
wire            n2989;
wire      [7:0] n2990;
wire            n2991;
wire      [7:0] n2992;
wire            n2993;
wire      [7:0] n2994;
wire            n2995;
wire      [7:0] n2996;
wire            n2997;
wire      [7:0] n2998;
wire            n2999;
wire      [7:0] n30;
wire            n300;
wire      [7:0] n3000;
wire            n3001;
wire      [7:0] n3002;
wire            n3003;
wire      [7:0] n3004;
wire            n3005;
wire      [7:0] n3006;
wire            n3007;
wire      [7:0] n3008;
wire            n3009;
wire      [7:0] n301;
wire      [7:0] n3010;
wire            n3011;
wire      [7:0] n3012;
wire            n3013;
wire      [7:0] n3014;
wire            n3015;
wire      [7:0] n3016;
wire            n3017;
wire      [7:0] n3018;
wire            n3019;
wire      [7:0] n3020;
wire            n3021;
wire      [7:0] n3022;
wire            n3023;
wire      [7:0] n3024;
wire            n3025;
wire      [7:0] n3026;
wire            n3027;
wire      [7:0] n3028;
wire            n3029;
wire            n303;
wire      [7:0] n3030;
wire            n3031;
wire      [7:0] n3032;
wire            n3033;
wire      [7:0] n3034;
wire            n3035;
wire      [7:0] n3036;
wire            n3037;
wire      [7:0] n3038;
wire            n3039;
wire      [7:0] n304;
wire      [7:0] n3040;
wire            n3041;
wire      [7:0] n3042;
wire            n3043;
wire      [7:0] n3044;
wire            n3045;
wire      [7:0] n3046;
wire            n3047;
wire      [7:0] n3048;
wire            n3049;
wire            n305;
wire      [7:0] n3050;
wire            n3051;
wire      [7:0] n3052;
wire            n3053;
wire      [7:0] n3054;
wire            n3055;
wire      [7:0] n3056;
wire            n3057;
wire      [7:0] n3058;
wire            n3059;
wire      [7:0] n306;
wire      [7:0] n3060;
wire            n3061;
wire      [7:0] n3062;
wire            n3063;
wire      [7:0] n3064;
wire            n3065;
wire      [7:0] n3066;
wire            n3067;
wire      [7:0] n3068;
wire            n3069;
wire      [7:0] n3070;
wire            n3071;
wire      [7:0] n3072;
wire            n3073;
wire      [7:0] n3074;
wire            n3075;
wire      [7:0] n3076;
wire      [7:0] n3077;
wire      [7:0] n3078;
wire      [7:0] n3079;
wire            n308;
wire      [7:0] n3080;
wire      [7:0] n3081;
wire      [7:0] n3082;
wire      [7:0] n3083;
wire      [7:0] n3084;
wire      [7:0] n3085;
wire      [7:0] n3086;
wire      [7:0] n3087;
wire      [7:0] n3088;
wire      [7:0] n3089;
wire      [7:0] n3090;
wire      [7:0] n3091;
wire      [7:0] n3092;
wire      [7:0] n3093;
wire      [7:0] n3094;
wire      [7:0] n3095;
wire      [7:0] n3096;
wire      [7:0] n3097;
wire      [7:0] n3098;
wire      [7:0] n3099;
wire      [7:0] n310;
wire      [7:0] n3100;
wire      [7:0] n3101;
wire      [7:0] n3102;
wire      [7:0] n3103;
wire      [7:0] n3104;
wire      [7:0] n3105;
wire      [7:0] n3106;
wire      [7:0] n3107;
wire      [7:0] n3108;
wire      [7:0] n3109;
wire            n311;
wire      [7:0] n3110;
wire      [7:0] n3111;
wire      [7:0] n3112;
wire      [7:0] n3113;
wire      [7:0] n3114;
wire      [7:0] n3115;
wire      [7:0] n3116;
wire      [7:0] n3117;
wire      [7:0] n3118;
wire      [7:0] n3119;
wire      [7:0] n3120;
wire      [7:0] n3121;
wire      [7:0] n3122;
wire      [7:0] n3123;
wire      [7:0] n3124;
wire      [7:0] n3125;
wire      [7:0] n3126;
wire      [7:0] n3127;
wire      [7:0] n3128;
wire      [7:0] n3129;
wire      [7:0] n313;
wire      [7:0] n3130;
wire      [7:0] n3131;
wire      [7:0] n3132;
wire      [7:0] n3133;
wire      [7:0] n3134;
wire      [7:0] n3135;
wire      [7:0] n3136;
wire      [7:0] n3137;
wire      [7:0] n3138;
wire      [7:0] n3139;
wire      [7:0] n3140;
wire      [7:0] n3141;
wire      [7:0] n3142;
wire      [7:0] n3143;
wire      [7:0] n3144;
wire      [7:0] n3145;
wire      [7:0] n3146;
wire      [7:0] n3147;
wire      [7:0] n3148;
wire      [7:0] n3149;
wire            n315;
wire      [7:0] n3150;
wire      [7:0] n3151;
wire      [7:0] n3152;
wire      [7:0] n3153;
wire      [7:0] n3154;
wire      [7:0] n3155;
wire      [7:0] n3156;
wire      [7:0] n3157;
wire      [7:0] n3158;
wire      [7:0] n3159;
wire      [7:0] n316;
wire      [7:0] n3160;
wire      [7:0] n3161;
wire      [7:0] n3162;
wire      [7:0] n3163;
wire      [7:0] n3164;
wire      [7:0] n3165;
wire      [7:0] n3166;
wire      [7:0] n3167;
wire      [7:0] n3168;
wire      [7:0] n3169;
wire            n317;
wire      [7:0] n3170;
wire      [7:0] n3171;
wire      [7:0] n3172;
wire      [7:0] n3173;
wire      [7:0] n3174;
wire      [7:0] n3175;
wire      [7:0] n3176;
wire      [7:0] n3177;
wire      [7:0] n3178;
wire      [7:0] n3179;
wire      [7:0] n3180;
wire      [7:0] n3181;
wire      [7:0] n3182;
wire      [7:0] n3183;
wire      [7:0] n3184;
wire      [7:0] n3185;
wire      [7:0] n3186;
wire      [7:0] n3187;
wire      [7:0] n3188;
wire      [7:0] n3189;
wire      [7:0] n319;
wire      [7:0] n3190;
wire      [7:0] n3191;
wire      [7:0] n3192;
wire      [7:0] n3193;
wire      [7:0] n3194;
wire      [7:0] n3195;
wire      [7:0] n3196;
wire      [7:0] n3197;
wire      [7:0] n3198;
wire      [7:0] n3199;
wire            n32;
wire            n320;
wire      [7:0] n3200;
wire      [7:0] n3201;
wire      [7:0] n3202;
wire      [7:0] n3203;
wire      [7:0] n3204;
wire      [7:0] n3205;
wire      [7:0] n3206;
wire      [7:0] n3207;
wire      [7:0] n3208;
wire      [7:0] n3209;
wire      [7:0] n321;
wire      [7:0] n3210;
wire      [7:0] n3211;
wire      [7:0] n3212;
wire      [7:0] n3213;
wire      [7:0] n3214;
wire      [7:0] n3215;
wire      [7:0] n3216;
wire      [7:0] n3217;
wire      [7:0] n3218;
wire      [7:0] n3219;
wire            n322;
wire      [7:0] n3220;
wire      [7:0] n3221;
wire      [7:0] n3222;
wire      [7:0] n3223;
wire      [7:0] n3224;
wire      [7:0] n3225;
wire      [7:0] n3226;
wire      [7:0] n3227;
wire      [7:0] n3228;
wire      [7:0] n3229;
wire      [7:0] n3230;
wire      [7:0] n3231;
wire      [7:0] n3232;
wire      [7:0] n3233;
wire      [7:0] n3234;
wire      [7:0] n3235;
wire      [7:0] n3236;
wire      [7:0] n3237;
wire      [7:0] n3238;
wire      [7:0] n3239;
wire      [7:0] n324;
wire      [7:0] n3240;
wire      [7:0] n3241;
wire      [7:0] n3242;
wire      [7:0] n3243;
wire      [7:0] n3244;
wire      [7:0] n3245;
wire      [7:0] n3246;
wire      [7:0] n3247;
wire      [7:0] n3248;
wire      [7:0] n3249;
wire      [7:0] n3250;
wire      [7:0] n3251;
wire      [7:0] n3252;
wire      [7:0] n3253;
wire      [7:0] n3254;
wire      [7:0] n3255;
wire      [7:0] n3256;
wire      [7:0] n3257;
wire      [7:0] n3258;
wire      [7:0] n3259;
wire            n326;
wire      [7:0] n3260;
wire      [7:0] n3261;
wire      [7:0] n3262;
wire      [7:0] n3263;
wire      [7:0] n3264;
wire      [7:0] n3265;
wire      [7:0] n3266;
wire      [7:0] n3267;
wire      [7:0] n3268;
wire      [7:0] n3269;
wire      [7:0] n327;
wire      [7:0] n3270;
wire      [7:0] n3271;
wire      [7:0] n3272;
wire      [7:0] n3273;
wire      [7:0] n3274;
wire      [7:0] n3275;
wire      [7:0] n3276;
wire      [7:0] n3277;
wire      [7:0] n3278;
wire      [7:0] n3279;
wire      [7:0] n3280;
wire      [7:0] n3281;
wire      [7:0] n3282;
wire      [7:0] n3283;
wire      [7:0] n3284;
wire      [7:0] n3285;
wire      [7:0] n3286;
wire      [7:0] n3287;
wire      [7:0] n3288;
wire      [7:0] n3289;
wire            n329;
wire      [7:0] n3290;
wire      [7:0] n3291;
wire      [7:0] n3292;
wire      [7:0] n3293;
wire      [7:0] n3294;
wire      [7:0] n3295;
wire      [7:0] n3296;
wire      [7:0] n3297;
wire      [7:0] n3298;
wire      [7:0] n3299;
wire      [7:0] n3300;
wire      [7:0] n3301;
wire      [7:0] n3302;
wire      [7:0] n3303;
wire      [7:0] n3304;
wire      [7:0] n3305;
wire      [7:0] n3306;
wire      [7:0] n3307;
wire      [7:0] n3308;
wire      [7:0] n3309;
wire      [7:0] n331;
wire      [7:0] n3310;
wire      [7:0] n3311;
wire      [7:0] n3312;
wire      [7:0] n3313;
wire      [7:0] n3314;
wire      [7:0] n3315;
wire      [7:0] n3316;
wire      [7:0] n3317;
wire      [7:0] n3318;
wire      [7:0] n3319;
wire            n332;
wire      [7:0] n3320;
wire      [7:0] n3321;
wire      [7:0] n3322;
wire      [7:0] n3323;
wire      [7:0] n3324;
wire      [7:0] n3325;
wire      [7:0] n3326;
wire      [7:0] n3327;
wire      [7:0] n3328;
wire      [7:0] n3329;
wire      [7:0] n3330;
wire      [7:0] n3331;
wire      [7:0] n3332;
wire      [7:0] n3333;
wire            n3334;
wire      [7:0] n3335;
wire            n3336;
wire      [7:0] n3337;
wire            n3338;
wire      [7:0] n3339;
wire      [7:0] n334;
wire            n3340;
wire      [7:0] n3341;
wire            n3342;
wire      [7:0] n3343;
wire            n3344;
wire      [7:0] n3345;
wire            n3346;
wire      [7:0] n3347;
wire            n3348;
wire      [7:0] n3349;
wire            n3350;
wire      [7:0] n3351;
wire            n3352;
wire      [7:0] n3353;
wire            n3354;
wire      [7:0] n3355;
wire            n3356;
wire      [7:0] n3357;
wire            n3358;
wire      [7:0] n3359;
wire            n336;
wire            n3360;
wire      [7:0] n3361;
wire            n3362;
wire      [7:0] n3363;
wire            n3364;
wire      [7:0] n3365;
wire            n3366;
wire      [7:0] n3367;
wire            n3368;
wire      [7:0] n3369;
wire            n3370;
wire      [7:0] n3371;
wire            n3372;
wire      [7:0] n3373;
wire            n3374;
wire      [7:0] n3375;
wire            n3376;
wire      [7:0] n3377;
wire            n3378;
wire      [7:0] n3379;
wire      [7:0] n338;
wire            n3380;
wire      [7:0] n3381;
wire            n3382;
wire      [7:0] n3383;
wire            n3384;
wire      [7:0] n3385;
wire            n3386;
wire      [7:0] n3387;
wire            n3388;
wire      [7:0] n3389;
wire            n3390;
wire      [7:0] n3391;
wire            n3392;
wire      [7:0] n3393;
wire            n3394;
wire      [7:0] n3395;
wire            n3396;
wire      [7:0] n3397;
wire            n3398;
wire      [7:0] n3399;
wire      [7:0] n34;
wire            n340;
wire            n3400;
wire      [7:0] n3401;
wire            n3402;
wire      [7:0] n3403;
wire            n3404;
wire      [7:0] n3405;
wire            n3406;
wire      [7:0] n3407;
wire            n3408;
wire      [7:0] n3409;
wire            n3410;
wire      [7:0] n3411;
wire            n3412;
wire      [7:0] n3413;
wire            n3414;
wire      [7:0] n3415;
wire            n3416;
wire      [7:0] n3417;
wire            n3418;
wire      [7:0] n3419;
wire      [7:0] n342;
wire            n3420;
wire      [7:0] n3421;
wire            n3422;
wire      [7:0] n3423;
wire            n3424;
wire      [7:0] n3425;
wire            n3426;
wire      [7:0] n3427;
wire            n3428;
wire      [7:0] n3429;
wire            n3430;
wire      [7:0] n3431;
wire            n3432;
wire      [7:0] n3433;
wire            n3434;
wire      [7:0] n3435;
wire            n3436;
wire      [7:0] n3437;
wire            n3438;
wire      [7:0] n3439;
wire            n344;
wire            n3440;
wire      [7:0] n3441;
wire            n3442;
wire      [7:0] n3443;
wire            n3444;
wire      [7:0] n3445;
wire            n3446;
wire      [7:0] n3447;
wire            n3448;
wire      [7:0] n3449;
wire            n3450;
wire      [7:0] n3451;
wire            n3452;
wire      [7:0] n3453;
wire            n3454;
wire      [7:0] n3455;
wire            n3456;
wire      [7:0] n3457;
wire            n3458;
wire      [7:0] n3459;
wire      [7:0] n346;
wire            n3460;
wire      [7:0] n3461;
wire            n3462;
wire      [7:0] n3463;
wire            n3464;
wire      [7:0] n3465;
wire            n3466;
wire      [7:0] n3467;
wire            n3468;
wire      [7:0] n3469;
wire            n347;
wire            n3470;
wire      [7:0] n3471;
wire            n3472;
wire      [7:0] n3473;
wire            n3474;
wire      [7:0] n3475;
wire            n3476;
wire      [7:0] n3477;
wire            n3478;
wire      [7:0] n3479;
wire            n3480;
wire      [7:0] n3481;
wire            n3482;
wire      [7:0] n3483;
wire            n3484;
wire      [7:0] n3485;
wire            n3486;
wire      [7:0] n3487;
wire            n3488;
wire      [7:0] n3489;
wire      [7:0] n349;
wire            n3490;
wire      [7:0] n3491;
wire            n3492;
wire      [7:0] n3493;
wire            n3494;
wire      [7:0] n3495;
wire            n3496;
wire      [7:0] n3497;
wire            n3498;
wire      [7:0] n3499;
wire            n3500;
wire      [7:0] n3501;
wire            n3502;
wire      [7:0] n3503;
wire            n3504;
wire      [7:0] n3505;
wire            n3506;
wire      [7:0] n3507;
wire            n3508;
wire      [7:0] n3509;
wire            n351;
wire            n3510;
wire      [7:0] n3511;
wire            n3512;
wire      [7:0] n3513;
wire            n3514;
wire      [7:0] n3515;
wire            n3516;
wire      [7:0] n3517;
wire            n3518;
wire      [7:0] n3519;
wire      [7:0] n352;
wire            n3520;
wire      [7:0] n3521;
wire            n3522;
wire      [7:0] n3523;
wire            n3524;
wire      [7:0] n3525;
wire            n3526;
wire      [7:0] n3527;
wire            n3528;
wire      [7:0] n3529;
wire            n353;
wire            n3530;
wire      [7:0] n3531;
wire            n3532;
wire      [7:0] n3533;
wire            n3534;
wire      [7:0] n3535;
wire            n3536;
wire      [7:0] n3537;
wire            n3538;
wire      [7:0] n3539;
wire      [7:0] n354;
wire            n3540;
wire      [7:0] n3541;
wire            n3542;
wire      [7:0] n3543;
wire            n3544;
wire      [7:0] n3545;
wire            n3546;
wire      [7:0] n3547;
wire            n3548;
wire      [7:0] n3549;
wire            n3550;
wire      [7:0] n3551;
wire            n3552;
wire      [7:0] n3553;
wire            n3554;
wire      [7:0] n3555;
wire            n3556;
wire      [7:0] n3557;
wire            n3558;
wire      [7:0] n3559;
wire            n356;
wire            n3560;
wire      [7:0] n3561;
wire            n3562;
wire      [7:0] n3563;
wire            n3564;
wire      [7:0] n3565;
wire            n3566;
wire      [7:0] n3567;
wire            n3568;
wire      [7:0] n3569;
wire            n3570;
wire      [7:0] n3571;
wire            n3572;
wire      [7:0] n3573;
wire            n3574;
wire      [7:0] n3575;
wire            n3576;
wire      [7:0] n3577;
wire            n3578;
wire      [7:0] n3579;
wire      [7:0] n358;
wire            n3580;
wire      [7:0] n3581;
wire            n3582;
wire      [7:0] n3583;
wire            n3584;
wire      [7:0] n3585;
wire            n3586;
wire      [7:0] n3587;
wire            n3588;
wire      [7:0] n3589;
wire            n3590;
wire      [7:0] n3591;
wire            n3592;
wire      [7:0] n3593;
wire            n3594;
wire      [7:0] n3595;
wire            n3596;
wire      [7:0] n3597;
wire            n3598;
wire      [7:0] n3599;
wire            n36;
wire            n360;
wire            n3600;
wire      [7:0] n3601;
wire            n3602;
wire      [7:0] n3603;
wire            n3604;
wire      [7:0] n3605;
wire            n3606;
wire      [7:0] n3607;
wire            n3608;
wire      [7:0] n3609;
wire      [7:0] n361;
wire            n3610;
wire      [7:0] n3611;
wire            n3612;
wire      [7:0] n3613;
wire            n3614;
wire      [7:0] n3615;
wire            n3616;
wire      [7:0] n3617;
wire            n3618;
wire      [7:0] n3619;
wire            n362;
wire            n3620;
wire      [7:0] n3621;
wire            n3622;
wire      [7:0] n3623;
wire            n3624;
wire      [7:0] n3625;
wire            n3626;
wire      [7:0] n3627;
wire            n3628;
wire      [7:0] n3629;
wire      [7:0] n363;
wire            n3630;
wire      [7:0] n3631;
wire            n3632;
wire      [7:0] n3633;
wire            n3634;
wire      [7:0] n3635;
wire            n3636;
wire      [7:0] n3637;
wire            n3638;
wire      [7:0] n3639;
wire            n3640;
wire      [7:0] n3641;
wire            n3642;
wire      [7:0] n3643;
wire            n3644;
wire      [7:0] n3645;
wire            n3646;
wire      [7:0] n3647;
wire            n3648;
wire      [7:0] n3649;
wire            n365;
wire            n3650;
wire      [7:0] n3651;
wire            n3652;
wire      [7:0] n3653;
wire            n3654;
wire      [7:0] n3655;
wire            n3656;
wire      [7:0] n3657;
wire            n3658;
wire      [7:0] n3659;
wire            n3660;
wire      [7:0] n3661;
wire            n3662;
wire      [7:0] n3663;
wire            n3664;
wire      [7:0] n3665;
wire            n3666;
wire      [7:0] n3667;
wire            n3668;
wire      [7:0] n3669;
wire      [7:0] n367;
wire            n3670;
wire      [7:0] n3671;
wire            n3672;
wire      [7:0] n3673;
wire            n3674;
wire      [7:0] n3675;
wire            n3676;
wire      [7:0] n3677;
wire            n3678;
wire      [7:0] n3679;
wire            n3680;
wire      [7:0] n3681;
wire            n3682;
wire      [7:0] n3683;
wire            n3684;
wire      [7:0] n3685;
wire            n3686;
wire      [7:0] n3687;
wire            n3688;
wire      [7:0] n3689;
wire            n369;
wire            n3690;
wire      [7:0] n3691;
wire            n3692;
wire      [7:0] n3693;
wire            n3694;
wire      [7:0] n3695;
wire            n3696;
wire      [7:0] n3697;
wire            n3698;
wire      [7:0] n3699;
wire            n3700;
wire      [7:0] n3701;
wire            n3702;
wire      [7:0] n3703;
wire            n3704;
wire      [7:0] n3705;
wire            n3706;
wire      [7:0] n3707;
wire            n3708;
wire      [7:0] n3709;
wire      [7:0] n371;
wire            n3710;
wire      [7:0] n3711;
wire            n3712;
wire      [7:0] n3713;
wire            n3714;
wire      [7:0] n3715;
wire            n3716;
wire      [7:0] n3717;
wire            n3718;
wire      [7:0] n3719;
wire            n372;
wire            n3720;
wire      [7:0] n3721;
wire            n3722;
wire      [7:0] n3723;
wire            n3724;
wire      [7:0] n3725;
wire            n3726;
wire      [7:0] n3727;
wire            n3728;
wire      [7:0] n3729;
wire      [7:0] n373;
wire            n3730;
wire      [7:0] n3731;
wire            n3732;
wire      [7:0] n3733;
wire            n3734;
wire      [7:0] n3735;
wire            n3736;
wire      [7:0] n3737;
wire            n3738;
wire      [7:0] n3739;
wire            n3740;
wire      [7:0] n3741;
wire            n3742;
wire      [7:0] n3743;
wire            n3744;
wire      [7:0] n3745;
wire            n3746;
wire      [7:0] n3747;
wire            n3748;
wire      [7:0] n3749;
wire            n375;
wire            n3750;
wire      [7:0] n3751;
wire            n3752;
wire      [7:0] n3753;
wire            n3754;
wire      [7:0] n3755;
wire            n3756;
wire      [7:0] n3757;
wire            n3758;
wire      [7:0] n3759;
wire            n3760;
wire      [7:0] n3761;
wire            n3762;
wire      [7:0] n3763;
wire            n3764;
wire      [7:0] n3765;
wire            n3766;
wire      [7:0] n3767;
wire            n3768;
wire      [7:0] n3769;
wire      [7:0] n377;
wire            n3770;
wire      [7:0] n3771;
wire            n3772;
wire      [7:0] n3773;
wire            n3774;
wire      [7:0] n3775;
wire            n3776;
wire      [7:0] n3777;
wire            n3778;
wire      [7:0] n3779;
wire            n378;
wire            n3780;
wire      [7:0] n3781;
wire            n3782;
wire      [7:0] n3783;
wire            n3784;
wire      [7:0] n3785;
wire            n3786;
wire      [7:0] n3787;
wire            n3788;
wire      [7:0] n3789;
wire            n3790;
wire      [7:0] n3791;
wire            n3792;
wire      [7:0] n3793;
wire            n3794;
wire      [7:0] n3795;
wire            n3796;
wire      [7:0] n3797;
wire            n3798;
wire      [7:0] n3799;
wire      [7:0] n38;
wire      [7:0] n380;
wire            n3800;
wire      [7:0] n3801;
wire            n3802;
wire      [7:0] n3803;
wire            n3804;
wire      [7:0] n3805;
wire            n3806;
wire      [7:0] n3807;
wire            n3808;
wire      [7:0] n3809;
wire            n381;
wire            n3810;
wire      [7:0] n3811;
wire            n3812;
wire      [7:0] n3813;
wire            n3814;
wire      [7:0] n3815;
wire            n3816;
wire      [7:0] n3817;
wire            n3818;
wire      [7:0] n3819;
wire            n3820;
wire      [7:0] n3821;
wire            n3822;
wire      [7:0] n3823;
wire            n3824;
wire      [7:0] n3825;
wire            n3826;
wire      [7:0] n3827;
wire            n3828;
wire      [7:0] n3829;
wire      [7:0] n383;
wire            n3830;
wire      [7:0] n3831;
wire            n3832;
wire      [7:0] n3833;
wire            n3834;
wire      [7:0] n3835;
wire            n3836;
wire      [7:0] n3837;
wire            n3838;
wire      [7:0] n3839;
wire            n3840;
wire      [7:0] n3841;
wire            n3842;
wire      [7:0] n3843;
wire            n3844;
wire      [7:0] n3845;
wire      [7:0] n3846;
wire      [7:0] n3847;
wire      [7:0] n3848;
wire      [7:0] n3849;
wire            n385;
wire      [7:0] n3850;
wire      [7:0] n3851;
wire      [7:0] n3852;
wire      [7:0] n3853;
wire      [7:0] n3854;
wire      [7:0] n3855;
wire      [7:0] n3856;
wire      [7:0] n3857;
wire      [7:0] n3858;
wire      [7:0] n3859;
wire      [7:0] n3860;
wire      [7:0] n3861;
wire      [7:0] n3862;
wire      [7:0] n3863;
wire      [7:0] n3864;
wire      [7:0] n3865;
wire      [7:0] n3866;
wire      [7:0] n3867;
wire      [7:0] n3868;
wire      [7:0] n3869;
wire      [7:0] n387;
wire      [7:0] n3870;
wire      [7:0] n3871;
wire      [7:0] n3872;
wire      [7:0] n3873;
wire      [7:0] n3874;
wire      [7:0] n3875;
wire      [7:0] n3876;
wire      [7:0] n3877;
wire      [7:0] n3878;
wire      [7:0] n3879;
wire      [7:0] n3880;
wire      [7:0] n3881;
wire      [7:0] n3882;
wire      [7:0] n3883;
wire      [7:0] n3884;
wire      [7:0] n3885;
wire      [7:0] n3886;
wire      [7:0] n3887;
wire      [7:0] n3888;
wire      [7:0] n3889;
wire            n389;
wire      [7:0] n3890;
wire      [7:0] n3891;
wire      [7:0] n3892;
wire      [7:0] n3893;
wire      [7:0] n3894;
wire      [7:0] n3895;
wire      [7:0] n3896;
wire      [7:0] n3897;
wire      [7:0] n3898;
wire      [7:0] n3899;
wire      [7:0] n3900;
wire      [7:0] n3901;
wire      [7:0] n3902;
wire      [7:0] n3903;
wire      [7:0] n3904;
wire      [7:0] n3905;
wire      [7:0] n3906;
wire      [7:0] n3907;
wire      [7:0] n3908;
wire      [7:0] n3909;
wire      [7:0] n391;
wire      [7:0] n3910;
wire      [7:0] n3911;
wire      [7:0] n3912;
wire      [7:0] n3913;
wire      [7:0] n3914;
wire      [7:0] n3915;
wire      [7:0] n3916;
wire      [7:0] n3917;
wire      [7:0] n3918;
wire      [7:0] n3919;
wire      [7:0] n3920;
wire      [7:0] n3921;
wire      [7:0] n3922;
wire      [7:0] n3923;
wire      [7:0] n3924;
wire      [7:0] n3925;
wire      [7:0] n3926;
wire      [7:0] n3927;
wire      [7:0] n3928;
wire      [7:0] n3929;
wire            n393;
wire      [7:0] n3930;
wire      [7:0] n3931;
wire      [7:0] n3932;
wire      [7:0] n3933;
wire      [7:0] n3934;
wire      [7:0] n3935;
wire      [7:0] n3936;
wire      [7:0] n3937;
wire      [7:0] n3938;
wire      [7:0] n3939;
wire      [7:0] n394;
wire      [7:0] n3940;
wire      [7:0] n3941;
wire      [7:0] n3942;
wire      [7:0] n3943;
wire      [7:0] n3944;
wire      [7:0] n3945;
wire      [7:0] n3946;
wire      [7:0] n3947;
wire      [7:0] n3948;
wire      [7:0] n3949;
wire            n395;
wire      [7:0] n3950;
wire      [7:0] n3951;
wire      [7:0] n3952;
wire      [7:0] n3953;
wire      [7:0] n3954;
wire      [7:0] n3955;
wire      [7:0] n3956;
wire      [7:0] n3957;
wire      [7:0] n3958;
wire      [7:0] n3959;
wire      [7:0] n396;
wire      [7:0] n3960;
wire      [7:0] n3961;
wire      [7:0] n3962;
wire      [7:0] n3963;
wire      [7:0] n3964;
wire      [7:0] n3965;
wire      [7:0] n3966;
wire      [7:0] n3967;
wire      [7:0] n3968;
wire      [7:0] n3969;
wire      [7:0] n3970;
wire      [7:0] n3971;
wire      [7:0] n3972;
wire      [7:0] n3973;
wire      [7:0] n3974;
wire      [7:0] n3975;
wire      [7:0] n3976;
wire      [7:0] n3977;
wire      [7:0] n3978;
wire      [7:0] n3979;
wire            n398;
wire      [7:0] n3980;
wire      [7:0] n3981;
wire      [7:0] n3982;
wire      [7:0] n3983;
wire      [7:0] n3984;
wire      [7:0] n3985;
wire      [7:0] n3986;
wire      [7:0] n3987;
wire      [7:0] n3988;
wire      [7:0] n3989;
wire      [7:0] n3990;
wire      [7:0] n3991;
wire      [7:0] n3992;
wire      [7:0] n3993;
wire      [7:0] n3994;
wire      [7:0] n3995;
wire      [7:0] n3996;
wire      [7:0] n3997;
wire      [7:0] n3998;
wire      [7:0] n3999;
wire            n4;
wire            n40;
wire      [7:0] n400;
wire      [7:0] n4000;
wire      [7:0] n4001;
wire      [7:0] n4002;
wire      [7:0] n4003;
wire      [7:0] n4004;
wire      [7:0] n4005;
wire      [7:0] n4006;
wire      [7:0] n4007;
wire      [7:0] n4008;
wire      [7:0] n4009;
wire            n401;
wire      [7:0] n4010;
wire      [7:0] n4011;
wire      [7:0] n4012;
wire      [7:0] n4013;
wire      [7:0] n4014;
wire      [7:0] n4015;
wire      [7:0] n4016;
wire      [7:0] n4017;
wire      [7:0] n4018;
wire      [7:0] n4019;
wire      [7:0] n402;
wire      [7:0] n4020;
wire      [7:0] n4021;
wire      [7:0] n4022;
wire      [7:0] n4023;
wire      [7:0] n4024;
wire      [7:0] n4025;
wire      [7:0] n4026;
wire      [7:0] n4027;
wire      [7:0] n4028;
wire      [7:0] n4029;
wire      [7:0] n4030;
wire      [7:0] n4031;
wire      [7:0] n4032;
wire      [7:0] n4033;
wire      [7:0] n4034;
wire      [7:0] n4035;
wire      [7:0] n4036;
wire      [7:0] n4037;
wire      [7:0] n4038;
wire      [7:0] n4039;
wire            n404;
wire      [7:0] n4040;
wire      [7:0] n4041;
wire      [7:0] n4042;
wire      [7:0] n4043;
wire      [7:0] n4044;
wire      [7:0] n4045;
wire      [7:0] n4046;
wire      [7:0] n4047;
wire      [7:0] n4048;
wire      [7:0] n4049;
wire      [7:0] n405;
wire      [7:0] n4050;
wire      [7:0] n4051;
wire      [7:0] n4052;
wire      [7:0] n4053;
wire      [7:0] n4054;
wire      [7:0] n4055;
wire      [7:0] n4056;
wire      [7:0] n4057;
wire      [7:0] n4058;
wire      [7:0] n4059;
wire      [7:0] n4060;
wire      [7:0] n4061;
wire      [7:0] n4062;
wire      [7:0] n4063;
wire      [7:0] n4064;
wire      [7:0] n4065;
wire      [7:0] n4066;
wire      [7:0] n4067;
wire      [7:0] n4068;
wire      [7:0] n4069;
wire            n407;
wire      [7:0] n4070;
wire      [7:0] n4071;
wire      [7:0] n4072;
wire      [7:0] n4073;
wire      [7:0] n4074;
wire      [7:0] n4075;
wire      [7:0] n4076;
wire      [7:0] n4077;
wire      [7:0] n4078;
wire      [7:0] n4079;
wire      [7:0] n4080;
wire      [7:0] n4081;
wire      [7:0] n4082;
wire      [7:0] n4083;
wire      [7:0] n4084;
wire      [7:0] n4085;
wire      [7:0] n4086;
wire      [7:0] n4087;
wire      [7:0] n4088;
wire      [7:0] n4089;
wire      [7:0] n409;
wire      [7:0] n4090;
wire      [7:0] n4091;
wire      [7:0] n4092;
wire      [7:0] n4093;
wire      [7:0] n4094;
wire      [7:0] n4095;
wire      [7:0] n4096;
wire      [7:0] n4097;
wire      [7:0] n4098;
wire      [7:0] n4099;
wire      [7:0] n4100;
wire      [7:0] n4101;
wire      [7:0] n4102;
wire      [7:0] n4103;
wire      [7:0] n4104;
wire            n4105;
wire      [7:0] n4106;
wire            n4107;
wire      [7:0] n4108;
wire            n4109;
wire            n411;
wire      [7:0] n4110;
wire            n4111;
wire      [7:0] n4112;
wire            n4113;
wire      [7:0] n4114;
wire            n4115;
wire      [7:0] n4116;
wire            n4117;
wire      [7:0] n4118;
wire            n4119;
wire      [7:0] n412;
wire      [7:0] n4120;
wire            n4121;
wire      [7:0] n4122;
wire            n4123;
wire      [7:0] n4124;
wire            n4125;
wire      [7:0] n4126;
wire            n4127;
wire      [7:0] n4128;
wire            n4129;
wire            n413;
wire      [7:0] n4130;
wire            n4131;
wire      [7:0] n4132;
wire            n4133;
wire      [7:0] n4134;
wire            n4135;
wire      [7:0] n4136;
wire            n4137;
wire      [7:0] n4138;
wire            n4139;
wire      [7:0] n414;
wire      [7:0] n4140;
wire            n4141;
wire      [7:0] n4142;
wire            n4143;
wire      [7:0] n4144;
wire            n4145;
wire      [7:0] n4146;
wire            n4147;
wire      [7:0] n4148;
wire            n4149;
wire            n415;
wire      [7:0] n4150;
wire            n4151;
wire      [7:0] n4152;
wire            n4153;
wire      [7:0] n4154;
wire            n4155;
wire      [7:0] n4156;
wire            n4157;
wire      [7:0] n4158;
wire            n4159;
wire      [7:0] n4160;
wire            n4161;
wire      [7:0] n4162;
wire            n4163;
wire      [7:0] n4164;
wire            n4165;
wire      [7:0] n4166;
wire            n4167;
wire      [7:0] n4168;
wire            n4169;
wire      [7:0] n417;
wire      [7:0] n4170;
wire            n4171;
wire      [7:0] n4172;
wire            n4173;
wire      [7:0] n4174;
wire            n4175;
wire      [7:0] n4176;
wire            n4177;
wire      [7:0] n4178;
wire            n4179;
wire      [7:0] n4180;
wire            n4181;
wire      [7:0] n4182;
wire            n4183;
wire      [7:0] n4184;
wire            n4185;
wire      [7:0] n4186;
wire            n4187;
wire      [7:0] n4188;
wire            n4189;
wire            n419;
wire      [7:0] n4190;
wire            n4191;
wire      [7:0] n4192;
wire            n4193;
wire      [7:0] n4194;
wire            n4195;
wire      [7:0] n4196;
wire            n4197;
wire      [7:0] n4198;
wire            n4199;
wire      [7:0] n42;
wire      [7:0] n420;
wire      [7:0] n4200;
wire            n4201;
wire      [7:0] n4202;
wire            n4203;
wire      [7:0] n4204;
wire            n4205;
wire      [7:0] n4206;
wire            n4207;
wire      [7:0] n4208;
wire            n4209;
wire      [7:0] n4210;
wire            n4211;
wire      [7:0] n4212;
wire            n4213;
wire      [7:0] n4214;
wire            n4215;
wire      [7:0] n4216;
wire            n4217;
wire      [7:0] n4218;
wire            n4219;
wire            n422;
wire      [7:0] n4220;
wire            n4221;
wire      [7:0] n4222;
wire            n4223;
wire      [7:0] n4224;
wire            n4225;
wire      [7:0] n4226;
wire            n4227;
wire      [7:0] n4228;
wire            n4229;
wire      [7:0] n4230;
wire            n4231;
wire      [7:0] n4232;
wire            n4233;
wire      [7:0] n4234;
wire            n4235;
wire      [7:0] n4236;
wire            n4237;
wire      [7:0] n4238;
wire            n4239;
wire      [7:0] n424;
wire      [7:0] n4240;
wire            n4241;
wire      [7:0] n4242;
wire            n4243;
wire      [7:0] n4244;
wire            n4245;
wire      [7:0] n4246;
wire            n4247;
wire      [7:0] n4248;
wire            n4249;
wire      [7:0] n4250;
wire            n4251;
wire      [7:0] n4252;
wire            n4253;
wire      [7:0] n4254;
wire            n4255;
wire      [7:0] n4256;
wire            n4257;
wire      [7:0] n4258;
wire            n4259;
wire            n426;
wire      [7:0] n4260;
wire            n4261;
wire      [7:0] n4262;
wire            n4263;
wire      [7:0] n4264;
wire            n4265;
wire      [7:0] n4266;
wire            n4267;
wire      [7:0] n4268;
wire            n4269;
wire      [7:0] n427;
wire      [7:0] n4270;
wire            n4271;
wire      [7:0] n4272;
wire            n4273;
wire      [7:0] n4274;
wire            n4275;
wire      [7:0] n4276;
wire            n4277;
wire      [7:0] n4278;
wire            n4279;
wire            n428;
wire      [7:0] n4280;
wire            n4281;
wire      [7:0] n4282;
wire            n4283;
wire      [7:0] n4284;
wire            n4285;
wire      [7:0] n4286;
wire            n4287;
wire      [7:0] n4288;
wire            n4289;
wire      [7:0] n4290;
wire            n4291;
wire      [7:0] n4292;
wire            n4293;
wire      [7:0] n4294;
wire            n4295;
wire      [7:0] n4296;
wire            n4297;
wire      [7:0] n4298;
wire            n4299;
wire      [7:0] n430;
wire      [7:0] n4300;
wire            n4301;
wire      [7:0] n4302;
wire            n4303;
wire      [7:0] n4304;
wire            n4305;
wire      [7:0] n4306;
wire            n4307;
wire      [7:0] n4308;
wire            n4309;
wire      [7:0] n4310;
wire            n4311;
wire      [7:0] n4312;
wire            n4313;
wire      [7:0] n4314;
wire            n4315;
wire      [7:0] n4316;
wire            n4317;
wire      [7:0] n4318;
wire            n4319;
wire            n432;
wire      [7:0] n4320;
wire            n4321;
wire      [7:0] n4322;
wire            n4323;
wire      [7:0] n4324;
wire            n4325;
wire      [7:0] n4326;
wire            n4327;
wire      [7:0] n4328;
wire            n4329;
wire      [7:0] n433;
wire      [7:0] n4330;
wire            n4331;
wire      [7:0] n4332;
wire            n4333;
wire      [7:0] n4334;
wire            n4335;
wire      [7:0] n4336;
wire            n4337;
wire      [7:0] n4338;
wire            n4339;
wire      [7:0] n4340;
wire            n4341;
wire      [7:0] n4342;
wire            n4343;
wire      [7:0] n4344;
wire            n4345;
wire      [7:0] n4346;
wire            n4347;
wire      [7:0] n4348;
wire            n4349;
wire            n435;
wire      [7:0] n4350;
wire            n4351;
wire      [7:0] n4352;
wire            n4353;
wire      [7:0] n4354;
wire            n4355;
wire      [7:0] n4356;
wire            n4357;
wire      [7:0] n4358;
wire            n4359;
wire      [7:0] n4360;
wire            n4361;
wire      [7:0] n4362;
wire            n4363;
wire      [7:0] n4364;
wire            n4365;
wire      [7:0] n4366;
wire            n4367;
wire      [7:0] n4368;
wire            n4369;
wire      [7:0] n437;
wire      [7:0] n4370;
wire            n4371;
wire      [7:0] n4372;
wire            n4373;
wire      [7:0] n4374;
wire            n4375;
wire      [7:0] n4376;
wire            n4377;
wire      [7:0] n4378;
wire            n4379;
wire            n438;
wire      [7:0] n4380;
wire            n4381;
wire      [7:0] n4382;
wire            n4383;
wire      [7:0] n4384;
wire            n4385;
wire      [7:0] n4386;
wire            n4387;
wire      [7:0] n4388;
wire            n4389;
wire      [7:0] n439;
wire      [7:0] n4390;
wire            n4391;
wire      [7:0] n4392;
wire            n4393;
wire      [7:0] n4394;
wire            n4395;
wire      [7:0] n4396;
wire            n4397;
wire      [7:0] n4398;
wire            n4399;
wire            n44;
wire      [7:0] n4400;
wire            n4401;
wire      [7:0] n4402;
wire            n4403;
wire      [7:0] n4404;
wire            n4405;
wire      [7:0] n4406;
wire            n4407;
wire      [7:0] n4408;
wire            n4409;
wire            n441;
wire      [7:0] n4410;
wire            n4411;
wire      [7:0] n4412;
wire            n4413;
wire      [7:0] n4414;
wire            n4415;
wire      [7:0] n4416;
wire            n4417;
wire      [7:0] n4418;
wire            n4419;
wire      [7:0] n442;
wire      [7:0] n4420;
wire            n4421;
wire      [7:0] n4422;
wire            n4423;
wire      [7:0] n4424;
wire            n4425;
wire      [7:0] n4426;
wire            n4427;
wire      [7:0] n4428;
wire            n4429;
wire            n443;
wire      [7:0] n4430;
wire            n4431;
wire      [7:0] n4432;
wire            n4433;
wire      [7:0] n4434;
wire            n4435;
wire      [7:0] n4436;
wire            n4437;
wire      [7:0] n4438;
wire            n4439;
wire      [7:0] n4440;
wire            n4441;
wire      [7:0] n4442;
wire            n4443;
wire      [7:0] n4444;
wire            n4445;
wire      [7:0] n4446;
wire            n4447;
wire      [7:0] n4448;
wire            n4449;
wire      [7:0] n445;
wire      [7:0] n4450;
wire            n4451;
wire      [7:0] n4452;
wire            n4453;
wire      [7:0] n4454;
wire            n4455;
wire      [7:0] n4456;
wire            n4457;
wire      [7:0] n4458;
wire            n4459;
wire      [7:0] n4460;
wire            n4461;
wire      [7:0] n4462;
wire            n4463;
wire      [7:0] n4464;
wire            n4465;
wire      [7:0] n4466;
wire            n4467;
wire      [7:0] n4468;
wire            n4469;
wire            n447;
wire      [7:0] n4470;
wire            n4471;
wire      [7:0] n4472;
wire            n4473;
wire      [7:0] n4474;
wire            n4475;
wire      [7:0] n4476;
wire            n4477;
wire      [7:0] n4478;
wire            n4479;
wire      [7:0] n4480;
wire            n4481;
wire      [7:0] n4482;
wire            n4483;
wire      [7:0] n4484;
wire            n4485;
wire      [7:0] n4486;
wire            n4487;
wire      [7:0] n4488;
wire            n4489;
wire      [7:0] n449;
wire      [7:0] n4490;
wire            n4491;
wire      [7:0] n4492;
wire            n4493;
wire      [7:0] n4494;
wire            n4495;
wire      [7:0] n4496;
wire            n4497;
wire      [7:0] n4498;
wire            n4499;
wire      [7:0] n4500;
wire            n4501;
wire      [7:0] n4502;
wire            n4503;
wire      [7:0] n4504;
wire            n4505;
wire      [7:0] n4506;
wire            n4507;
wire      [7:0] n4508;
wire            n4509;
wire            n451;
wire      [7:0] n4510;
wire            n4511;
wire      [7:0] n4512;
wire            n4513;
wire      [7:0] n4514;
wire            n4515;
wire      [7:0] n4516;
wire            n4517;
wire      [7:0] n4518;
wire            n4519;
wire      [7:0] n452;
wire      [7:0] n4520;
wire            n4521;
wire      [7:0] n4522;
wire            n4523;
wire      [7:0] n4524;
wire            n4525;
wire      [7:0] n4526;
wire            n4527;
wire      [7:0] n4528;
wire            n4529;
wire      [7:0] n4530;
wire            n4531;
wire      [7:0] n4532;
wire            n4533;
wire      [7:0] n4534;
wire            n4535;
wire      [7:0] n4536;
wire            n4537;
wire      [7:0] n4538;
wire            n4539;
wire            n454;
wire      [7:0] n4540;
wire            n4541;
wire      [7:0] n4542;
wire            n4543;
wire      [7:0] n4544;
wire            n4545;
wire      [7:0] n4546;
wire            n4547;
wire      [7:0] n4548;
wire            n4549;
wire      [7:0] n455;
wire      [7:0] n4550;
wire            n4551;
wire      [7:0] n4552;
wire            n4553;
wire      [7:0] n4554;
wire            n4555;
wire      [7:0] n4556;
wire            n4557;
wire      [7:0] n4558;
wire            n4559;
wire      [7:0] n4560;
wire            n4561;
wire      [7:0] n4562;
wire            n4563;
wire      [7:0] n4564;
wire            n4565;
wire      [7:0] n4566;
wire            n4567;
wire      [7:0] n4568;
wire            n4569;
wire            n457;
wire      [7:0] n4570;
wire            n4571;
wire      [7:0] n4572;
wire            n4573;
wire      [7:0] n4574;
wire            n4575;
wire      [7:0] n4576;
wire            n4577;
wire      [7:0] n4578;
wire            n4579;
wire      [7:0] n458;
wire      [7:0] n4580;
wire            n4581;
wire      [7:0] n4582;
wire            n4583;
wire      [7:0] n4584;
wire            n4585;
wire      [7:0] n4586;
wire            n4587;
wire      [7:0] n4588;
wire            n4589;
wire      [7:0] n4590;
wire            n4591;
wire      [7:0] n4592;
wire            n4593;
wire      [7:0] n4594;
wire            n4595;
wire      [7:0] n4596;
wire            n4597;
wire      [7:0] n4598;
wire            n4599;
wire      [7:0] n46;
wire            n460;
wire      [7:0] n4600;
wire            n4601;
wire      [7:0] n4602;
wire            n4603;
wire      [7:0] n4604;
wire            n4605;
wire      [7:0] n4606;
wire            n4607;
wire      [7:0] n4608;
wire            n4609;
wire      [7:0] n461;
wire      [7:0] n4610;
wire            n4611;
wire      [7:0] n4612;
wire            n4613;
wire      [7:0] n4614;
wire            n4615;
wire      [7:0] n4616;
wire      [7:0] n4617;
wire      [7:0] n4618;
wire      [7:0] n4619;
wire            n462;
wire      [7:0] n4620;
wire      [7:0] n4621;
wire      [7:0] n4622;
wire      [7:0] n4623;
wire      [7:0] n4624;
wire      [7:0] n4625;
wire      [7:0] n4626;
wire      [7:0] n4627;
wire      [7:0] n4628;
wire      [7:0] n4629;
wire      [7:0] n4630;
wire      [7:0] n4631;
wire      [7:0] n4632;
wire      [7:0] n4633;
wire      [7:0] n4634;
wire      [7:0] n4635;
wire      [7:0] n4636;
wire      [7:0] n4637;
wire      [7:0] n4638;
wire      [7:0] n4639;
wire      [7:0] n464;
wire      [7:0] n4640;
wire      [7:0] n4641;
wire      [7:0] n4642;
wire      [7:0] n4643;
wire      [7:0] n4644;
wire      [7:0] n4645;
wire      [7:0] n4646;
wire      [7:0] n4647;
wire      [7:0] n4648;
wire      [7:0] n4649;
wire            n465;
wire      [7:0] n4650;
wire      [7:0] n4651;
wire      [7:0] n4652;
wire      [7:0] n4653;
wire      [7:0] n4654;
wire      [7:0] n4655;
wire      [7:0] n4656;
wire      [7:0] n4657;
wire      [7:0] n4658;
wire      [7:0] n4659;
wire      [7:0] n4660;
wire      [7:0] n4661;
wire      [7:0] n4662;
wire      [7:0] n4663;
wire      [7:0] n4664;
wire      [7:0] n4665;
wire      [7:0] n4666;
wire      [7:0] n4667;
wire      [7:0] n4668;
wire      [7:0] n4669;
wire      [7:0] n467;
wire      [7:0] n4670;
wire      [7:0] n4671;
wire      [7:0] n4672;
wire      [7:0] n4673;
wire      [7:0] n4674;
wire      [7:0] n4675;
wire      [7:0] n4676;
wire      [7:0] n4677;
wire      [7:0] n4678;
wire      [7:0] n4679;
wire            n468;
wire      [7:0] n4680;
wire      [7:0] n4681;
wire      [7:0] n4682;
wire      [7:0] n4683;
wire      [7:0] n4684;
wire      [7:0] n4685;
wire      [7:0] n4686;
wire      [7:0] n4687;
wire      [7:0] n4688;
wire      [7:0] n4689;
wire      [7:0] n469;
wire      [7:0] n4690;
wire      [7:0] n4691;
wire      [7:0] n4692;
wire      [7:0] n4693;
wire      [7:0] n4694;
wire      [7:0] n4695;
wire      [7:0] n4696;
wire      [7:0] n4697;
wire      [7:0] n4698;
wire      [7:0] n4699;
wire      [7:0] n4700;
wire      [7:0] n4701;
wire      [7:0] n4702;
wire      [7:0] n4703;
wire      [7:0] n4704;
wire      [7:0] n4705;
wire      [7:0] n4706;
wire      [7:0] n4707;
wire      [7:0] n4708;
wire      [7:0] n4709;
wire            n471;
wire      [7:0] n4710;
wire      [7:0] n4711;
wire      [7:0] n4712;
wire      [7:0] n4713;
wire      [7:0] n4714;
wire      [7:0] n4715;
wire      [7:0] n4716;
wire      [7:0] n4717;
wire      [7:0] n4718;
wire      [7:0] n4719;
wire      [7:0] n4720;
wire      [7:0] n4721;
wire      [7:0] n4722;
wire      [7:0] n4723;
wire      [7:0] n4724;
wire      [7:0] n4725;
wire      [7:0] n4726;
wire      [7:0] n4727;
wire      [7:0] n4728;
wire      [7:0] n4729;
wire      [7:0] n473;
wire      [7:0] n4730;
wire      [7:0] n4731;
wire      [7:0] n4732;
wire      [7:0] n4733;
wire      [7:0] n4734;
wire      [7:0] n4735;
wire      [7:0] n4736;
wire      [7:0] n4737;
wire      [7:0] n4738;
wire      [7:0] n4739;
wire      [7:0] n4740;
wire      [7:0] n4741;
wire      [7:0] n4742;
wire      [7:0] n4743;
wire      [7:0] n4744;
wire      [7:0] n4745;
wire      [7:0] n4746;
wire      [7:0] n4747;
wire      [7:0] n4748;
wire      [7:0] n4749;
wire            n475;
wire      [7:0] n4750;
wire      [7:0] n4751;
wire      [7:0] n4752;
wire      [7:0] n4753;
wire      [7:0] n4754;
wire      [7:0] n4755;
wire      [7:0] n4756;
wire      [7:0] n4757;
wire      [7:0] n4758;
wire      [7:0] n4759;
wire      [7:0] n4760;
wire      [7:0] n4761;
wire      [7:0] n4762;
wire      [7:0] n4763;
wire      [7:0] n4764;
wire      [7:0] n4765;
wire      [7:0] n4766;
wire      [7:0] n4767;
wire      [7:0] n4768;
wire      [7:0] n4769;
wire      [7:0] n477;
wire      [7:0] n4770;
wire      [7:0] n4771;
wire      [7:0] n4772;
wire      [7:0] n4773;
wire      [7:0] n4774;
wire      [7:0] n4775;
wire      [7:0] n4776;
wire      [7:0] n4777;
wire      [7:0] n4778;
wire      [7:0] n4779;
wire            n478;
wire      [7:0] n4780;
wire      [7:0] n4781;
wire      [7:0] n4782;
wire      [7:0] n4783;
wire      [7:0] n4784;
wire      [7:0] n4785;
wire      [7:0] n4786;
wire      [7:0] n4787;
wire      [7:0] n4788;
wire      [7:0] n4789;
wire      [7:0] n479;
wire      [7:0] n4790;
wire      [7:0] n4791;
wire      [7:0] n4792;
wire      [7:0] n4793;
wire      [7:0] n4794;
wire      [7:0] n4795;
wire      [7:0] n4796;
wire      [7:0] n4797;
wire      [7:0] n4798;
wire      [7:0] n4799;
wire            n48;
wire      [7:0] n4800;
wire      [7:0] n4801;
wire      [7:0] n4802;
wire      [7:0] n4803;
wire      [7:0] n4804;
wire      [7:0] n4805;
wire      [7:0] n4806;
wire      [7:0] n4807;
wire      [7:0] n4808;
wire      [7:0] n4809;
wire            n481;
wire      [7:0] n4810;
wire      [7:0] n4811;
wire      [7:0] n4812;
wire      [7:0] n4813;
wire      [7:0] n4814;
wire      [7:0] n4815;
wire      [7:0] n4816;
wire      [7:0] n4817;
wire      [7:0] n4818;
wire      [7:0] n4819;
wire      [7:0] n4820;
wire      [7:0] n4821;
wire      [7:0] n4822;
wire      [7:0] n4823;
wire      [7:0] n4824;
wire      [7:0] n4825;
wire      [7:0] n4826;
wire      [7:0] n4827;
wire      [7:0] n4828;
wire      [7:0] n4829;
wire      [7:0] n483;
wire      [7:0] n4830;
wire      [7:0] n4831;
wire      [7:0] n4832;
wire      [7:0] n4833;
wire      [7:0] n4834;
wire      [7:0] n4835;
wire      [7:0] n4836;
wire      [7:0] n4837;
wire      [7:0] n4838;
wire      [7:0] n4839;
wire      [7:0] n4840;
wire      [7:0] n4841;
wire      [7:0] n4842;
wire      [7:0] n4843;
wire      [7:0] n4844;
wire      [7:0] n4845;
wire      [7:0] n4846;
wire      [7:0] n4847;
wire      [7:0] n4848;
wire      [7:0] n4849;
wire            n485;
wire      [7:0] n4850;
wire      [7:0] n4851;
wire      [7:0] n4852;
wire      [7:0] n4853;
wire      [7:0] n4854;
wire      [7:0] n4855;
wire      [7:0] n4856;
wire      [7:0] n4857;
wire      [7:0] n4858;
wire      [7:0] n4859;
wire      [7:0] n4860;
wire      [7:0] n4861;
wire      [7:0] n4862;
wire      [7:0] n4863;
wire      [7:0] n4864;
wire      [7:0] n4865;
wire      [7:0] n4866;
wire      [7:0] n4867;
wire      [7:0] n4868;
wire      [7:0] n4869;
wire      [7:0] n487;
wire      [7:0] n4870;
wire      [7:0] n4871;
wire      [7:0] n4872;
wire      [7:0] n4873;
wire      [7:0] n4874;
wire            n4875;
wire      [7:0] n4876;
wire            n4877;
wire      [7:0] n4878;
wire            n4879;
wire            n488;
wire      [7:0] n4880;
wire            n4881;
wire      [7:0] n4882;
wire            n4883;
wire      [7:0] n4884;
wire            n4885;
wire      [7:0] n4886;
wire            n4887;
wire      [7:0] n4888;
wire            n4889;
wire      [7:0] n4890;
wire            n4891;
wire      [7:0] n4892;
wire            n4893;
wire      [7:0] n4894;
wire            n4895;
wire      [7:0] n4896;
wire            n4897;
wire      [7:0] n4898;
wire            n4899;
wire      [7:0] n490;
wire      [7:0] n4900;
wire            n4901;
wire      [7:0] n4902;
wire            n4903;
wire      [7:0] n4904;
wire            n4905;
wire      [7:0] n4906;
wire            n4907;
wire      [7:0] n4908;
wire            n4909;
wire            n491;
wire      [7:0] n4910;
wire            n4911;
wire      [7:0] n4912;
wire            n4913;
wire      [7:0] n4914;
wire            n4915;
wire      [7:0] n4916;
wire            n4917;
wire      [7:0] n4918;
wire            n4919;
wire      [7:0] n4920;
wire            n4921;
wire      [7:0] n4922;
wire            n4923;
wire      [7:0] n4924;
wire            n4925;
wire      [7:0] n4926;
wire            n4927;
wire      [7:0] n4928;
wire            n4929;
wire      [7:0] n493;
wire      [7:0] n4930;
wire            n4931;
wire      [7:0] n4932;
wire            n4933;
wire      [7:0] n4934;
wire            n4935;
wire      [7:0] n4936;
wire            n4937;
wire      [7:0] n4938;
wire            n4939;
wire      [7:0] n4940;
wire            n4941;
wire      [7:0] n4942;
wire            n4943;
wire      [7:0] n4944;
wire            n4945;
wire      [7:0] n4946;
wire            n4947;
wire      [7:0] n4948;
wire            n4949;
wire            n495;
wire      [7:0] n4950;
wire            n4951;
wire      [7:0] n4952;
wire            n4953;
wire      [7:0] n4954;
wire            n4955;
wire      [7:0] n4956;
wire            n4957;
wire      [7:0] n4958;
wire            n4959;
wire      [7:0] n496;
wire      [7:0] n4960;
wire            n4961;
wire      [7:0] n4962;
wire            n4963;
wire      [7:0] n4964;
wire            n4965;
wire      [7:0] n4966;
wire            n4967;
wire      [7:0] n4968;
wire            n4969;
wire            n497;
wire      [7:0] n4970;
wire            n4971;
wire      [7:0] n4972;
wire            n4973;
wire      [7:0] n4974;
wire            n4975;
wire      [7:0] n4976;
wire            n4977;
wire      [7:0] n4978;
wire            n4979;
wire      [7:0] n4980;
wire            n4981;
wire      [7:0] n4982;
wire            n4983;
wire      [7:0] n4984;
wire            n4985;
wire      [7:0] n4986;
wire            n4987;
wire      [7:0] n4988;
wire            n4989;
wire      [7:0] n499;
wire      [7:0] n4990;
wire            n4991;
wire      [7:0] n4992;
wire            n4993;
wire      [7:0] n4994;
wire            n4995;
wire      [7:0] n4996;
wire            n4997;
wire      [7:0] n4998;
wire            n4999;
wire      [7:0] n50;
wire            n500;
wire      [7:0] n5000;
wire            n5001;
wire      [7:0] n5002;
wire            n5003;
wire      [7:0] n5004;
wire            n5005;
wire      [7:0] n5006;
wire            n5007;
wire      [7:0] n5008;
wire            n5009;
wire      [7:0] n501;
wire      [7:0] n5010;
wire            n5011;
wire      [7:0] n5012;
wire            n5013;
wire      [7:0] n5014;
wire            n5015;
wire      [7:0] n5016;
wire            n5017;
wire      [7:0] n5018;
wire            n5019;
wire            n502;
wire      [7:0] n5020;
wire            n5021;
wire      [7:0] n5022;
wire            n5023;
wire      [7:0] n5024;
wire            n5025;
wire      [7:0] n5026;
wire            n5027;
wire      [7:0] n5028;
wire            n5029;
wire      [7:0] n5030;
wire            n5031;
wire      [7:0] n5032;
wire            n5033;
wire      [7:0] n5034;
wire            n5035;
wire      [7:0] n5036;
wire            n5037;
wire      [7:0] n5038;
wire            n5039;
wire      [7:0] n504;
wire      [7:0] n5040;
wire            n5041;
wire      [7:0] n5042;
wire            n5043;
wire      [7:0] n5044;
wire            n5045;
wire      [7:0] n5046;
wire            n5047;
wire      [7:0] n5048;
wire            n5049;
wire            n505;
wire      [7:0] n5050;
wire            n5051;
wire      [7:0] n5052;
wire            n5053;
wire      [7:0] n5054;
wire            n5055;
wire      [7:0] n5056;
wire            n5057;
wire      [7:0] n5058;
wire            n5059;
wire      [7:0] n5060;
wire            n5061;
wire      [7:0] n5062;
wire            n5063;
wire      [7:0] n5064;
wire            n5065;
wire      [7:0] n5066;
wire            n5067;
wire      [7:0] n5068;
wire            n5069;
wire      [7:0] n507;
wire      [7:0] n5070;
wire            n5071;
wire      [7:0] n5072;
wire            n5073;
wire      [7:0] n5074;
wire            n5075;
wire      [7:0] n5076;
wire            n5077;
wire      [7:0] n5078;
wire            n5079;
wire            n508;
wire      [7:0] n5080;
wire            n5081;
wire      [7:0] n5082;
wire            n5083;
wire      [7:0] n5084;
wire            n5085;
wire      [7:0] n5086;
wire            n5087;
wire      [7:0] n5088;
wire            n5089;
wire      [7:0] n509;
wire      [7:0] n5090;
wire            n5091;
wire      [7:0] n5092;
wire            n5093;
wire      [7:0] n5094;
wire            n5095;
wire      [7:0] n5096;
wire            n5097;
wire      [7:0] n5098;
wire            n5099;
wire      [7:0] n5100;
wire            n5101;
wire      [7:0] n5102;
wire            n5103;
wire      [7:0] n5104;
wire            n5105;
wire      [7:0] n5106;
wire            n5107;
wire      [7:0] n5108;
wire            n5109;
wire            n511;
wire      [7:0] n5110;
wire            n5111;
wire      [7:0] n5112;
wire            n5113;
wire      [7:0] n5114;
wire            n5115;
wire      [7:0] n5116;
wire            n5117;
wire      [7:0] n5118;
wire            n5119;
wire      [7:0] n512;
wire      [7:0] n5120;
wire            n5121;
wire      [7:0] n5122;
wire            n5123;
wire      [7:0] n5124;
wire            n5125;
wire      [7:0] n5126;
wire            n5127;
wire      [7:0] n5128;
wire            n5129;
wire            n513;
wire      [7:0] n5130;
wire            n5131;
wire      [7:0] n5132;
wire            n5133;
wire      [7:0] n5134;
wire            n5135;
wire      [7:0] n5136;
wire            n5137;
wire      [7:0] n5138;
wire            n5139;
wire      [7:0] n514;
wire      [7:0] n5140;
wire            n5141;
wire      [7:0] n5142;
wire            n5143;
wire      [7:0] n5144;
wire            n5145;
wire      [7:0] n5146;
wire            n5147;
wire      [7:0] n5148;
wire            n5149;
wire            n515;
wire      [7:0] n5150;
wire            n5151;
wire      [7:0] n5152;
wire            n5153;
wire      [7:0] n5154;
wire            n5155;
wire      [7:0] n5156;
wire            n5157;
wire      [7:0] n5158;
wire            n5159;
wire      [7:0] n5160;
wire            n5161;
wire      [7:0] n5162;
wire            n5163;
wire      [7:0] n5164;
wire            n5165;
wire      [7:0] n5166;
wire            n5167;
wire      [7:0] n5168;
wire            n5169;
wire      [7:0] n517;
wire      [7:0] n5170;
wire            n5171;
wire      [7:0] n5172;
wire            n5173;
wire      [7:0] n5174;
wire            n5175;
wire      [7:0] n5176;
wire            n5177;
wire      [7:0] n5178;
wire            n5179;
wire            n518;
wire      [7:0] n5180;
wire            n5181;
wire      [7:0] n5182;
wire            n5183;
wire      [7:0] n5184;
wire            n5185;
wire      [7:0] n5186;
wire            n5187;
wire      [7:0] n5188;
wire            n5189;
wire      [7:0] n519;
wire      [7:0] n5190;
wire            n5191;
wire      [7:0] n5192;
wire            n5193;
wire      [7:0] n5194;
wire            n5195;
wire      [7:0] n5196;
wire            n5197;
wire      [7:0] n5198;
wire            n5199;
wire            n52;
wire      [7:0] n5200;
wire            n5201;
wire      [7:0] n5202;
wire            n5203;
wire      [7:0] n5204;
wire            n5205;
wire      [7:0] n5206;
wire            n5207;
wire      [7:0] n5208;
wire            n5209;
wire            n521;
wire      [7:0] n5210;
wire            n5211;
wire      [7:0] n5212;
wire            n5213;
wire      [7:0] n5214;
wire            n5215;
wire      [7:0] n5216;
wire            n5217;
wire      [7:0] n5218;
wire            n5219;
wire      [7:0] n522;
wire      [7:0] n5220;
wire            n5221;
wire      [7:0] n5222;
wire            n5223;
wire      [7:0] n5224;
wire            n5225;
wire      [7:0] n5226;
wire            n5227;
wire      [7:0] n5228;
wire            n5229;
wire      [7:0] n5230;
wire            n5231;
wire      [7:0] n5232;
wire            n5233;
wire      [7:0] n5234;
wire            n5235;
wire      [7:0] n5236;
wire            n5237;
wire      [7:0] n5238;
wire            n5239;
wire            n524;
wire      [7:0] n5240;
wire            n5241;
wire      [7:0] n5242;
wire            n5243;
wire      [7:0] n5244;
wire            n5245;
wire      [7:0] n5246;
wire            n5247;
wire      [7:0] n5248;
wire            n5249;
wire      [7:0] n5250;
wire            n5251;
wire      [7:0] n5252;
wire            n5253;
wire      [7:0] n5254;
wire            n5255;
wire      [7:0] n5256;
wire            n5257;
wire      [7:0] n5258;
wire            n5259;
wire      [7:0] n526;
wire      [7:0] n5260;
wire            n5261;
wire      [7:0] n5262;
wire            n5263;
wire      [7:0] n5264;
wire            n5265;
wire      [7:0] n5266;
wire            n5267;
wire      [7:0] n5268;
wire            n5269;
wire      [7:0] n5270;
wire            n5271;
wire      [7:0] n5272;
wire            n5273;
wire      [7:0] n5274;
wire            n5275;
wire      [7:0] n5276;
wire            n5277;
wire      [7:0] n5278;
wire            n5279;
wire            n528;
wire      [7:0] n5280;
wire            n5281;
wire      [7:0] n5282;
wire            n5283;
wire      [7:0] n5284;
wire            n5285;
wire      [7:0] n5286;
wire            n5287;
wire      [7:0] n5288;
wire            n5289;
wire      [7:0] n529;
wire      [7:0] n5290;
wire            n5291;
wire      [7:0] n5292;
wire            n5293;
wire      [7:0] n5294;
wire            n5295;
wire      [7:0] n5296;
wire            n5297;
wire      [7:0] n5298;
wire            n5299;
wire            n530;
wire      [7:0] n5300;
wire            n5301;
wire      [7:0] n5302;
wire            n5303;
wire      [7:0] n5304;
wire            n5305;
wire      [7:0] n5306;
wire            n5307;
wire      [7:0] n5308;
wire            n5309;
wire      [7:0] n531;
wire      [7:0] n5310;
wire            n5311;
wire      [7:0] n5312;
wire            n5313;
wire      [7:0] n5314;
wire            n5315;
wire      [7:0] n5316;
wire            n5317;
wire      [7:0] n5318;
wire            n5319;
wire            n532;
wire      [7:0] n5320;
wire            n5321;
wire      [7:0] n5322;
wire            n5323;
wire      [7:0] n5324;
wire            n5325;
wire      [7:0] n5326;
wire            n5327;
wire      [7:0] n5328;
wire            n5329;
wire      [7:0] n533;
wire      [7:0] n5330;
wire            n5331;
wire      [7:0] n5332;
wire            n5333;
wire      [7:0] n5334;
wire            n5335;
wire      [7:0] n5336;
wire            n5337;
wire      [7:0] n5338;
wire            n5339;
wire            n534;
wire      [7:0] n5340;
wire            n5341;
wire      [7:0] n5342;
wire            n5343;
wire      [7:0] n5344;
wire            n5345;
wire      [7:0] n5346;
wire            n5347;
wire      [7:0] n5348;
wire            n5349;
wire      [7:0] n535;
wire      [7:0] n5350;
wire            n5351;
wire      [7:0] n5352;
wire            n5353;
wire      [7:0] n5354;
wire            n5355;
wire      [7:0] n5356;
wire            n5357;
wire      [7:0] n5358;
wire            n5359;
wire      [7:0] n5360;
wire            n5361;
wire      [7:0] n5362;
wire            n5363;
wire      [7:0] n5364;
wire            n5365;
wire      [7:0] n5366;
wire            n5367;
wire      [7:0] n5368;
wire            n5369;
wire            n537;
wire      [7:0] n5370;
wire            n5371;
wire      [7:0] n5372;
wire            n5373;
wire      [7:0] n5374;
wire            n5375;
wire      [7:0] n5376;
wire            n5377;
wire      [7:0] n5378;
wire            n5379;
wire      [7:0] n5380;
wire            n5381;
wire      [7:0] n5382;
wire            n5383;
wire      [7:0] n5384;
wire            n5385;
wire      [7:0] n5386;
wire      [7:0] n5387;
wire      [7:0] n5388;
wire      [7:0] n5389;
wire      [7:0] n539;
wire      [7:0] n5390;
wire      [7:0] n5391;
wire      [7:0] n5392;
wire      [7:0] n5393;
wire      [7:0] n5394;
wire      [7:0] n5395;
wire      [7:0] n5396;
wire      [7:0] n5397;
wire      [7:0] n5398;
wire      [7:0] n5399;
wire      [7:0] n54;
wire            n540;
wire      [7:0] n5400;
wire      [7:0] n5401;
wire      [7:0] n5402;
wire      [7:0] n5403;
wire      [7:0] n5404;
wire      [7:0] n5405;
wire      [7:0] n5406;
wire      [7:0] n5407;
wire      [7:0] n5408;
wire      [7:0] n5409;
wire      [7:0] n541;
wire      [7:0] n5410;
wire      [7:0] n5411;
wire      [7:0] n5412;
wire      [7:0] n5413;
wire      [7:0] n5414;
wire      [7:0] n5415;
wire      [7:0] n5416;
wire      [7:0] n5417;
wire      [7:0] n5418;
wire      [7:0] n5419;
wire      [7:0] n5420;
wire      [7:0] n5421;
wire      [7:0] n5422;
wire      [7:0] n5423;
wire      [7:0] n5424;
wire      [7:0] n5425;
wire      [7:0] n5426;
wire      [7:0] n5427;
wire      [7:0] n5428;
wire      [7:0] n5429;
wire            n543;
wire      [7:0] n5430;
wire      [7:0] n5431;
wire      [7:0] n5432;
wire      [7:0] n5433;
wire      [7:0] n5434;
wire      [7:0] n5435;
wire      [7:0] n5436;
wire      [7:0] n5437;
wire      [7:0] n5438;
wire      [7:0] n5439;
wire      [7:0] n544;
wire      [7:0] n5440;
wire      [7:0] n5441;
wire      [7:0] n5442;
wire      [7:0] n5443;
wire      [7:0] n5444;
wire      [7:0] n5445;
wire      [7:0] n5446;
wire      [7:0] n5447;
wire      [7:0] n5448;
wire      [7:0] n5449;
wire      [7:0] n5450;
wire      [7:0] n5451;
wire      [7:0] n5452;
wire      [7:0] n5453;
wire      [7:0] n5454;
wire      [7:0] n5455;
wire      [7:0] n5456;
wire      [7:0] n5457;
wire      [7:0] n5458;
wire      [7:0] n5459;
wire            n546;
wire      [7:0] n5460;
wire      [7:0] n5461;
wire      [7:0] n5462;
wire      [7:0] n5463;
wire      [7:0] n5464;
wire      [7:0] n5465;
wire      [7:0] n5466;
wire      [7:0] n5467;
wire      [7:0] n5468;
wire      [7:0] n5469;
wire      [7:0] n547;
wire      [7:0] n5470;
wire      [7:0] n5471;
wire      [7:0] n5472;
wire      [7:0] n5473;
wire      [7:0] n5474;
wire      [7:0] n5475;
wire      [7:0] n5476;
wire      [7:0] n5477;
wire      [7:0] n5478;
wire      [7:0] n5479;
wire      [7:0] n5480;
wire      [7:0] n5481;
wire      [7:0] n5482;
wire      [7:0] n5483;
wire      [7:0] n5484;
wire      [7:0] n5485;
wire      [7:0] n5486;
wire      [7:0] n5487;
wire      [7:0] n5488;
wire      [7:0] n5489;
wire            n549;
wire      [7:0] n5490;
wire      [7:0] n5491;
wire      [7:0] n5492;
wire      [7:0] n5493;
wire      [7:0] n5494;
wire      [7:0] n5495;
wire      [7:0] n5496;
wire      [7:0] n5497;
wire      [7:0] n5498;
wire      [7:0] n5499;
wire      [7:0] n550;
wire      [7:0] n5500;
wire      [7:0] n5501;
wire      [7:0] n5502;
wire      [7:0] n5503;
wire      [7:0] n5504;
wire      [7:0] n5505;
wire      [7:0] n5506;
wire      [7:0] n5507;
wire      [7:0] n5508;
wire      [7:0] n5509;
wire            n551;
wire      [7:0] n5510;
wire      [7:0] n5511;
wire      [7:0] n5512;
wire      [7:0] n5513;
wire      [7:0] n5514;
wire      [7:0] n5515;
wire      [7:0] n5516;
wire      [7:0] n5517;
wire      [7:0] n5518;
wire      [7:0] n5519;
wire      [7:0] n552;
wire      [7:0] n5520;
wire      [7:0] n5521;
wire      [7:0] n5522;
wire      [7:0] n5523;
wire      [7:0] n5524;
wire      [7:0] n5525;
wire      [7:0] n5526;
wire      [7:0] n5527;
wire      [7:0] n5528;
wire      [7:0] n5529;
wire            n553;
wire      [7:0] n5530;
wire      [7:0] n5531;
wire      [7:0] n5532;
wire      [7:0] n5533;
wire      [7:0] n5534;
wire      [7:0] n5535;
wire      [7:0] n5536;
wire      [7:0] n5537;
wire      [7:0] n5538;
wire      [7:0] n5539;
wire      [7:0] n554;
wire      [7:0] n5540;
wire      [7:0] n5541;
wire      [7:0] n5542;
wire      [7:0] n5543;
wire      [7:0] n5544;
wire      [7:0] n5545;
wire      [7:0] n5546;
wire      [7:0] n5547;
wire      [7:0] n5548;
wire      [7:0] n5549;
wire      [7:0] n5550;
wire      [7:0] n5551;
wire      [7:0] n5552;
wire      [7:0] n5553;
wire      [7:0] n5554;
wire      [7:0] n5555;
wire      [7:0] n5556;
wire      [7:0] n5557;
wire      [7:0] n5558;
wire      [7:0] n5559;
wire            n556;
wire      [7:0] n5560;
wire      [7:0] n5561;
wire      [7:0] n5562;
wire      [7:0] n5563;
wire      [7:0] n5564;
wire      [7:0] n5565;
wire      [7:0] n5566;
wire      [7:0] n5567;
wire      [7:0] n5568;
wire      [7:0] n5569;
wire      [7:0] n557;
wire      [7:0] n5570;
wire      [7:0] n5571;
wire      [7:0] n5572;
wire      [7:0] n5573;
wire      [7:0] n5574;
wire      [7:0] n5575;
wire      [7:0] n5576;
wire      [7:0] n5577;
wire      [7:0] n5578;
wire      [7:0] n5579;
wire            n558;
wire      [7:0] n5580;
wire      [7:0] n5581;
wire      [7:0] n5582;
wire      [7:0] n5583;
wire      [7:0] n5584;
wire      [7:0] n5585;
wire      [7:0] n5586;
wire      [7:0] n5587;
wire      [7:0] n5588;
wire      [7:0] n5589;
wire      [7:0] n559;
wire      [7:0] n5590;
wire      [7:0] n5591;
wire      [7:0] n5592;
wire      [7:0] n5593;
wire      [7:0] n5594;
wire      [7:0] n5595;
wire      [7:0] n5596;
wire      [7:0] n5597;
wire      [7:0] n5598;
wire      [7:0] n5599;
wire            n56;
wire            n560;
wire      [7:0] n5600;
wire      [7:0] n5601;
wire      [7:0] n5602;
wire      [7:0] n5603;
wire      [7:0] n5604;
wire      [7:0] n5605;
wire      [7:0] n5606;
wire      [7:0] n5607;
wire      [7:0] n5608;
wire      [7:0] n5609;
wire      [7:0] n561;
wire      [7:0] n5610;
wire      [7:0] n5611;
wire      [7:0] n5612;
wire      [7:0] n5613;
wire      [7:0] n5614;
wire      [7:0] n5615;
wire      [7:0] n5616;
wire      [7:0] n5617;
wire      [7:0] n5618;
wire      [7:0] n5619;
wire      [7:0] n5620;
wire      [7:0] n5621;
wire      [7:0] n5622;
wire      [7:0] n5623;
wire      [7:0] n5624;
wire      [7:0] n5625;
wire      [7:0] n5626;
wire      [7:0] n5627;
wire      [7:0] n5628;
wire      [7:0] n5629;
wire            n563;
wire      [7:0] n5630;
wire      [7:0] n5631;
wire      [7:0] n5632;
wire      [7:0] n5633;
wire      [7:0] n5634;
wire      [7:0] n5635;
wire      [7:0] n5636;
wire      [7:0] n5637;
wire      [7:0] n5638;
wire      [7:0] n5639;
wire      [7:0] n564;
wire      [7:0] n5640;
wire      [7:0] n5641;
wire      [7:0] n5642;
wire      [7:0] n5643;
wire      [7:0] n5644;
wire      [7:0] n5645;
wire     [15:0] n5646;
wire      [7:0] n5647;
wire      [7:0] n5648;
wire      [7:0] n5649;
wire            n565;
wire      [7:0] n5650;
wire            n5651;
wire      [7:0] n5652;
wire            n5653;
wire      [7:0] n5654;
wire            n5655;
wire      [7:0] n5656;
wire            n5657;
wire      [7:0] n5658;
wire            n5659;
wire      [7:0] n566;
wire      [7:0] n5660;
wire            n5661;
wire      [7:0] n5662;
wire            n5663;
wire      [7:0] n5664;
wire            n5665;
wire      [7:0] n5666;
wire            n5667;
wire      [7:0] n5668;
wire            n5669;
wire      [7:0] n5670;
wire            n5671;
wire      [7:0] n5672;
wire            n5673;
wire      [7:0] n5674;
wire            n5675;
wire      [7:0] n5676;
wire            n5677;
wire      [7:0] n5678;
wire            n5679;
wire            n568;
wire      [7:0] n5680;
wire            n5681;
wire      [7:0] n5682;
wire            n5683;
wire      [7:0] n5684;
wire            n5685;
wire      [7:0] n5686;
wire            n5687;
wire      [7:0] n5688;
wire            n5689;
wire      [7:0] n569;
wire      [7:0] n5690;
wire            n5691;
wire      [7:0] n5692;
wire            n5693;
wire      [7:0] n5694;
wire            n5695;
wire      [7:0] n5696;
wire            n5697;
wire      [7:0] n5698;
wire            n5699;
wire            n570;
wire      [7:0] n5700;
wire            n5701;
wire      [7:0] n5702;
wire            n5703;
wire      [7:0] n5704;
wire            n5705;
wire      [7:0] n5706;
wire            n5707;
wire      [7:0] n5708;
wire            n5709;
wire      [7:0] n571;
wire      [7:0] n5710;
wire            n5711;
wire      [7:0] n5712;
wire            n5713;
wire      [7:0] n5714;
wire            n5715;
wire      [7:0] n5716;
wire            n5717;
wire      [7:0] n5718;
wire            n5719;
wire            n572;
wire      [7:0] n5720;
wire            n5721;
wire      [7:0] n5722;
wire            n5723;
wire      [7:0] n5724;
wire            n5725;
wire      [7:0] n5726;
wire            n5727;
wire      [7:0] n5728;
wire            n5729;
wire      [7:0] n5730;
wire            n5731;
wire      [7:0] n5732;
wire            n5733;
wire      [7:0] n5734;
wire            n5735;
wire      [7:0] n5736;
wire            n5737;
wire      [7:0] n5738;
wire            n5739;
wire      [7:0] n574;
wire      [7:0] n5740;
wire            n5741;
wire      [7:0] n5742;
wire            n5743;
wire      [7:0] n5744;
wire            n5745;
wire      [7:0] n5746;
wire            n5747;
wire      [7:0] n5748;
wire            n5749;
wire      [7:0] n5750;
wire            n5751;
wire      [7:0] n5752;
wire            n5753;
wire      [7:0] n5754;
wire            n5755;
wire      [7:0] n5756;
wire            n5757;
wire      [7:0] n5758;
wire            n5759;
wire            n576;
wire      [7:0] n5760;
wire            n5761;
wire      [7:0] n5762;
wire            n5763;
wire      [7:0] n5764;
wire            n5765;
wire      [7:0] n5766;
wire            n5767;
wire      [7:0] n5768;
wire            n5769;
wire      [7:0] n577;
wire      [7:0] n5770;
wire            n5771;
wire      [7:0] n5772;
wire            n5773;
wire      [7:0] n5774;
wire            n5775;
wire      [7:0] n5776;
wire            n5777;
wire      [7:0] n5778;
wire            n5779;
wire      [7:0] n5780;
wire            n5781;
wire      [7:0] n5782;
wire            n5783;
wire      [7:0] n5784;
wire            n5785;
wire      [7:0] n5786;
wire            n5787;
wire      [7:0] n5788;
wire            n5789;
wire            n579;
wire      [7:0] n5790;
wire            n5791;
wire      [7:0] n5792;
wire            n5793;
wire      [7:0] n5794;
wire            n5795;
wire      [7:0] n5796;
wire            n5797;
wire      [7:0] n5798;
wire            n5799;
wire      [7:0] n58;
wire      [7:0] n5800;
wire            n5801;
wire      [7:0] n5802;
wire            n5803;
wire      [7:0] n5804;
wire            n5805;
wire      [7:0] n5806;
wire            n5807;
wire      [7:0] n5808;
wire            n5809;
wire      [7:0] n581;
wire      [7:0] n5810;
wire            n5811;
wire      [7:0] n5812;
wire            n5813;
wire      [7:0] n5814;
wire            n5815;
wire      [7:0] n5816;
wire            n5817;
wire      [7:0] n5818;
wire            n5819;
wire      [7:0] n5820;
wire            n5821;
wire      [7:0] n5822;
wire            n5823;
wire      [7:0] n5824;
wire            n5825;
wire      [7:0] n5826;
wire            n5827;
wire      [7:0] n5828;
wire            n5829;
wire            n583;
wire      [7:0] n5830;
wire            n5831;
wire      [7:0] n5832;
wire            n5833;
wire      [7:0] n5834;
wire            n5835;
wire      [7:0] n5836;
wire            n5837;
wire      [7:0] n5838;
wire            n5839;
wire      [7:0] n584;
wire      [7:0] n5840;
wire            n5841;
wire      [7:0] n5842;
wire            n5843;
wire      [7:0] n5844;
wire            n5845;
wire      [7:0] n5846;
wire            n5847;
wire      [7:0] n5848;
wire            n5849;
wire            n585;
wire      [7:0] n5850;
wire            n5851;
wire      [7:0] n5852;
wire            n5853;
wire      [7:0] n5854;
wire            n5855;
wire      [7:0] n5856;
wire            n5857;
wire      [7:0] n5858;
wire            n5859;
wire      [7:0] n586;
wire      [7:0] n5860;
wire            n5861;
wire      [7:0] n5862;
wire            n5863;
wire      [7:0] n5864;
wire            n5865;
wire      [7:0] n5866;
wire            n5867;
wire      [7:0] n5868;
wire            n5869;
wire            n587;
wire      [7:0] n5870;
wire            n5871;
wire      [7:0] n5872;
wire            n5873;
wire      [7:0] n5874;
wire            n5875;
wire      [7:0] n5876;
wire            n5877;
wire      [7:0] n5878;
wire            n5879;
wire      [7:0] n5880;
wire            n5881;
wire      [7:0] n5882;
wire            n5883;
wire      [7:0] n5884;
wire            n5885;
wire      [7:0] n5886;
wire            n5887;
wire      [7:0] n5888;
wire            n5889;
wire      [7:0] n589;
wire      [7:0] n5890;
wire            n5891;
wire      [7:0] n5892;
wire            n5893;
wire      [7:0] n5894;
wire            n5895;
wire      [7:0] n5896;
wire            n5897;
wire      [7:0] n5898;
wire            n5899;
wire      [7:0] n5900;
wire            n5901;
wire      [7:0] n5902;
wire            n5903;
wire      [7:0] n5904;
wire            n5905;
wire      [7:0] n5906;
wire            n5907;
wire      [7:0] n5908;
wire            n5909;
wire            n591;
wire      [7:0] n5910;
wire            n5911;
wire      [7:0] n5912;
wire            n5913;
wire      [7:0] n5914;
wire            n5915;
wire      [7:0] n5916;
wire            n5917;
wire      [7:0] n5918;
wire            n5919;
wire      [7:0] n592;
wire      [7:0] n5920;
wire            n5921;
wire      [7:0] n5922;
wire            n5923;
wire      [7:0] n5924;
wire            n5925;
wire      [7:0] n5926;
wire            n5927;
wire      [7:0] n5928;
wire            n5929;
wire      [7:0] n5930;
wire            n5931;
wire      [7:0] n5932;
wire            n5933;
wire      [7:0] n5934;
wire            n5935;
wire      [7:0] n5936;
wire            n5937;
wire      [7:0] n5938;
wire            n5939;
wire            n594;
wire      [7:0] n5940;
wire            n5941;
wire      [7:0] n5942;
wire            n5943;
wire      [7:0] n5944;
wire            n5945;
wire      [7:0] n5946;
wire            n5947;
wire      [7:0] n5948;
wire            n5949;
wire      [7:0] n595;
wire      [7:0] n5950;
wire            n5951;
wire      [7:0] n5952;
wire            n5953;
wire      [7:0] n5954;
wire            n5955;
wire      [7:0] n5956;
wire            n5957;
wire      [7:0] n5958;
wire            n5959;
wire      [7:0] n5960;
wire            n5961;
wire      [7:0] n5962;
wire            n5963;
wire      [7:0] n5964;
wire            n5965;
wire      [7:0] n5966;
wire            n5967;
wire      [7:0] n5968;
wire            n5969;
wire            n597;
wire      [7:0] n5970;
wire            n5971;
wire      [7:0] n5972;
wire            n5973;
wire      [7:0] n5974;
wire            n5975;
wire      [7:0] n5976;
wire            n5977;
wire      [7:0] n5978;
wire            n5979;
wire      [7:0] n598;
wire      [7:0] n5980;
wire            n5981;
wire      [7:0] n5982;
wire            n5983;
wire      [7:0] n5984;
wire            n5985;
wire      [7:0] n5986;
wire            n5987;
wire      [7:0] n5988;
wire            n5989;
wire            n599;
wire      [7:0] n5990;
wire            n5991;
wire      [7:0] n5992;
wire            n5993;
wire      [7:0] n5994;
wire            n5995;
wire      [7:0] n5996;
wire            n5997;
wire      [7:0] n5998;
wire            n5999;
wire      [7:0] n6;
wire            n60;
wire      [7:0] n600;
wire      [7:0] n6000;
wire            n6001;
wire      [7:0] n6002;
wire            n6003;
wire      [7:0] n6004;
wire            n6005;
wire      [7:0] n6006;
wire            n6007;
wire      [7:0] n6008;
wire            n6009;
wire            n601;
wire      [7:0] n6010;
wire            n6011;
wire      [7:0] n6012;
wire            n6013;
wire      [7:0] n6014;
wire            n6015;
wire      [7:0] n6016;
wire            n6017;
wire      [7:0] n6018;
wire            n6019;
wire      [7:0] n602;
wire      [7:0] n6020;
wire            n6021;
wire      [7:0] n6022;
wire            n6023;
wire      [7:0] n6024;
wire            n6025;
wire      [7:0] n6026;
wire            n6027;
wire      [7:0] n6028;
wire            n6029;
wire            n603;
wire      [7:0] n6030;
wire            n6031;
wire      [7:0] n6032;
wire            n6033;
wire      [7:0] n6034;
wire            n6035;
wire      [7:0] n6036;
wire            n6037;
wire      [7:0] n6038;
wire            n6039;
wire      [7:0] n604;
wire      [7:0] n6040;
wire            n6041;
wire      [7:0] n6042;
wire            n6043;
wire      [7:0] n6044;
wire            n6045;
wire      [7:0] n6046;
wire            n6047;
wire      [7:0] n6048;
wire            n6049;
wire            n605;
wire      [7:0] n6050;
wire            n6051;
wire      [7:0] n6052;
wire            n6053;
wire      [7:0] n6054;
wire            n6055;
wire      [7:0] n6056;
wire            n6057;
wire      [7:0] n6058;
wire            n6059;
wire      [7:0] n606;
wire      [7:0] n6060;
wire            n6061;
wire      [7:0] n6062;
wire            n6063;
wire      [7:0] n6064;
wire            n6065;
wire      [7:0] n6066;
wire            n6067;
wire      [7:0] n6068;
wire            n6069;
wire            n607;
wire      [7:0] n6070;
wire            n6071;
wire      [7:0] n6072;
wire            n6073;
wire      [7:0] n6074;
wire            n6075;
wire      [7:0] n6076;
wire            n6077;
wire      [7:0] n6078;
wire            n6079;
wire      [7:0] n608;
wire      [7:0] n6080;
wire            n6081;
wire      [7:0] n6082;
wire            n6083;
wire      [7:0] n6084;
wire            n6085;
wire      [7:0] n6086;
wire            n6087;
wire      [7:0] n6088;
wire            n6089;
wire      [7:0] n6090;
wire            n6091;
wire      [7:0] n6092;
wire            n6093;
wire      [7:0] n6094;
wire            n6095;
wire      [7:0] n6096;
wire            n6097;
wire      [7:0] n6098;
wire            n6099;
wire            n610;
wire      [7:0] n6100;
wire            n6101;
wire      [7:0] n6102;
wire            n6103;
wire      [7:0] n6104;
wire            n6105;
wire      [7:0] n6106;
wire            n6107;
wire      [7:0] n6108;
wire            n6109;
wire      [7:0] n611;
wire      [7:0] n6110;
wire            n6111;
wire      [7:0] n6112;
wire            n6113;
wire      [7:0] n6114;
wire            n6115;
wire      [7:0] n6116;
wire            n6117;
wire      [7:0] n6118;
wire            n6119;
wire      [7:0] n6120;
wire            n6121;
wire      [7:0] n6122;
wire            n6123;
wire      [7:0] n6124;
wire            n6125;
wire      [7:0] n6126;
wire            n6127;
wire      [7:0] n6128;
wire            n6129;
wire            n613;
wire      [7:0] n6130;
wire            n6131;
wire      [7:0] n6132;
wire            n6133;
wire      [7:0] n6134;
wire            n6135;
wire      [7:0] n6136;
wire            n6137;
wire      [7:0] n6138;
wire            n6139;
wire      [7:0] n614;
wire      [7:0] n6140;
wire            n6141;
wire      [7:0] n6142;
wire            n6143;
wire      [7:0] n6144;
wire            n6145;
wire      [7:0] n6146;
wire            n6147;
wire      [7:0] n6148;
wire            n6149;
wire            n615;
wire      [7:0] n6150;
wire            n6151;
wire      [7:0] n6152;
wire            n6153;
wire      [7:0] n6154;
wire            n6155;
wire      [7:0] n6156;
wire            n6157;
wire      [7:0] n6158;
wire            n6159;
wire      [7:0] n6160;
wire            n6161;
wire      [7:0] n6162;
wire      [7:0] n6163;
wire      [7:0] n6164;
wire      [7:0] n6165;
wire      [7:0] n6166;
wire      [7:0] n6167;
wire      [7:0] n6168;
wire      [7:0] n6169;
wire      [7:0] n617;
wire      [7:0] n6170;
wire      [7:0] n6171;
wire      [7:0] n6172;
wire      [7:0] n6173;
wire      [7:0] n6174;
wire      [7:0] n6175;
wire      [7:0] n6176;
wire      [7:0] n6177;
wire      [7:0] n6178;
wire      [7:0] n6179;
wire            n618;
wire      [7:0] n6180;
wire      [7:0] n6181;
wire      [7:0] n6182;
wire      [7:0] n6183;
wire      [7:0] n6184;
wire      [7:0] n6185;
wire      [7:0] n6186;
wire      [7:0] n6187;
wire      [7:0] n6188;
wire      [7:0] n6189;
wire      [7:0] n6190;
wire      [7:0] n6191;
wire      [7:0] n6192;
wire      [7:0] n6193;
wire      [7:0] n6194;
wire      [7:0] n6195;
wire      [7:0] n6196;
wire      [7:0] n6197;
wire      [7:0] n6198;
wire      [7:0] n6199;
wire      [7:0] n62;
wire      [7:0] n620;
wire      [7:0] n6200;
wire      [7:0] n6201;
wire      [7:0] n6202;
wire      [7:0] n6203;
wire      [7:0] n6204;
wire      [7:0] n6205;
wire      [7:0] n6206;
wire      [7:0] n6207;
wire      [7:0] n6208;
wire      [7:0] n6209;
wire            n621;
wire      [7:0] n6210;
wire      [7:0] n6211;
wire      [7:0] n6212;
wire      [7:0] n6213;
wire      [7:0] n6214;
wire      [7:0] n6215;
wire      [7:0] n6216;
wire      [7:0] n6217;
wire      [7:0] n6218;
wire      [7:0] n6219;
wire      [7:0] n622;
wire      [7:0] n6220;
wire      [7:0] n6221;
wire      [7:0] n6222;
wire      [7:0] n6223;
wire      [7:0] n6224;
wire      [7:0] n6225;
wire      [7:0] n6226;
wire      [7:0] n6227;
wire      [7:0] n6228;
wire      [7:0] n6229;
wire      [7:0] n6230;
wire      [7:0] n6231;
wire      [7:0] n6232;
wire      [7:0] n6233;
wire      [7:0] n6234;
wire      [7:0] n6235;
wire      [7:0] n6236;
wire      [7:0] n6237;
wire      [7:0] n6238;
wire      [7:0] n6239;
wire            n624;
wire      [7:0] n6240;
wire      [7:0] n6241;
wire      [7:0] n6242;
wire      [7:0] n6243;
wire      [7:0] n6244;
wire      [7:0] n6245;
wire      [7:0] n6246;
wire      [7:0] n6247;
wire      [7:0] n6248;
wire      [7:0] n6249;
wire      [7:0] n6250;
wire      [7:0] n6251;
wire      [7:0] n6252;
wire      [7:0] n6253;
wire      [7:0] n6254;
wire      [7:0] n6255;
wire      [7:0] n6256;
wire      [7:0] n6257;
wire      [7:0] n6258;
wire      [7:0] n6259;
wire      [7:0] n626;
wire      [7:0] n6260;
wire      [7:0] n6261;
wire      [7:0] n6262;
wire      [7:0] n6263;
wire      [7:0] n6264;
wire      [7:0] n6265;
wire      [7:0] n6266;
wire      [7:0] n6267;
wire      [7:0] n6268;
wire      [7:0] n6269;
wire            n627;
wire      [7:0] n6270;
wire      [7:0] n6271;
wire      [7:0] n6272;
wire      [7:0] n6273;
wire      [7:0] n6274;
wire      [7:0] n6275;
wire      [7:0] n6276;
wire      [7:0] n6277;
wire      [7:0] n6278;
wire      [7:0] n6279;
wire      [7:0] n6280;
wire      [7:0] n6281;
wire      [7:0] n6282;
wire      [7:0] n6283;
wire      [7:0] n6284;
wire      [7:0] n6285;
wire      [7:0] n6286;
wire      [7:0] n6287;
wire      [7:0] n6288;
wire      [7:0] n6289;
wire      [7:0] n629;
wire      [7:0] n6290;
wire      [7:0] n6291;
wire      [7:0] n6292;
wire      [7:0] n6293;
wire      [7:0] n6294;
wire      [7:0] n6295;
wire      [7:0] n6296;
wire      [7:0] n6297;
wire      [7:0] n6298;
wire      [7:0] n6299;
wire            n630;
wire      [7:0] n6300;
wire      [7:0] n6301;
wire      [7:0] n6302;
wire      [7:0] n6303;
wire      [7:0] n6304;
wire      [7:0] n6305;
wire      [7:0] n6306;
wire      [7:0] n6307;
wire      [7:0] n6308;
wire      [7:0] n6309;
wire      [7:0] n631;
wire      [7:0] n6310;
wire      [7:0] n6311;
wire      [7:0] n6312;
wire      [7:0] n6313;
wire      [7:0] n6314;
wire      [7:0] n6315;
wire      [7:0] n6316;
wire      [7:0] n6317;
wire      [7:0] n6318;
wire      [7:0] n6319;
wire            n632;
wire      [7:0] n6320;
wire      [7:0] n6321;
wire      [7:0] n6322;
wire      [7:0] n6323;
wire      [7:0] n6324;
wire      [7:0] n6325;
wire      [7:0] n6326;
wire      [7:0] n6327;
wire      [7:0] n6328;
wire      [7:0] n6329;
wire      [7:0] n633;
wire      [7:0] n6330;
wire      [7:0] n6331;
wire      [7:0] n6332;
wire      [7:0] n6333;
wire      [7:0] n6334;
wire      [7:0] n6335;
wire      [7:0] n6336;
wire      [7:0] n6337;
wire      [7:0] n6338;
wire      [7:0] n6339;
wire      [7:0] n6340;
wire      [7:0] n6341;
wire      [7:0] n6342;
wire      [7:0] n6343;
wire      [7:0] n6344;
wire      [7:0] n6345;
wire      [7:0] n6346;
wire      [7:0] n6347;
wire      [7:0] n6348;
wire      [7:0] n6349;
wire            n635;
wire      [7:0] n6350;
wire      [7:0] n6351;
wire      [7:0] n6352;
wire      [7:0] n6353;
wire      [7:0] n6354;
wire      [7:0] n6355;
wire      [7:0] n6356;
wire      [7:0] n6357;
wire      [7:0] n6358;
wire      [7:0] n6359;
wire      [7:0] n636;
wire      [7:0] n6360;
wire      [7:0] n6361;
wire      [7:0] n6362;
wire      [7:0] n6363;
wire      [7:0] n6364;
wire      [7:0] n6365;
wire      [7:0] n6366;
wire      [7:0] n6367;
wire      [7:0] n6368;
wire      [7:0] n6369;
wire            n637;
wire      [7:0] n6370;
wire      [7:0] n6371;
wire      [7:0] n6372;
wire      [7:0] n6373;
wire      [7:0] n6374;
wire      [7:0] n6375;
wire      [7:0] n6376;
wire      [7:0] n6377;
wire      [7:0] n6378;
wire      [7:0] n6379;
wire      [7:0] n638;
wire      [7:0] n6380;
wire      [7:0] n6381;
wire      [7:0] n6382;
wire      [7:0] n6383;
wire      [7:0] n6384;
wire      [7:0] n6385;
wire      [7:0] n6386;
wire      [7:0] n6387;
wire      [7:0] n6388;
wire      [7:0] n6389;
wire            n639;
wire      [7:0] n6390;
wire      [7:0] n6391;
wire      [7:0] n6392;
wire      [7:0] n6393;
wire      [7:0] n6394;
wire      [7:0] n6395;
wire      [7:0] n6396;
wire      [7:0] n6397;
wire      [7:0] n6398;
wire      [7:0] n6399;
wire            n64;
wire      [7:0] n640;
wire      [7:0] n6400;
wire      [7:0] n6401;
wire      [7:0] n6402;
wire      [7:0] n6403;
wire      [7:0] n6404;
wire      [7:0] n6405;
wire      [7:0] n6406;
wire      [7:0] n6407;
wire      [7:0] n6408;
wire      [7:0] n6409;
wire            n641;
wire      [7:0] n6410;
wire      [7:0] n6411;
wire      [7:0] n6412;
wire      [7:0] n6413;
wire      [7:0] n6414;
wire      [7:0] n6415;
wire      [7:0] n6416;
wire      [7:0] n6417;
wire      [7:0] n6418;
wire      [7:0] n6419;
wire      [7:0] n6420;
wire     [23:0] n6421;
wire      [7:0] n6422;
wire      [7:0] n6423;
wire      [7:0] n6424;
wire      [7:0] n6425;
wire      [7:0] n6426;
wire      [7:0] n6427;
wire     [31:0] n6428;
wire      [7:0] n6429;
wire      [7:0] n643;
wire            n6430;
wire      [7:0] n6431;
wire            n6432;
wire      [7:0] n6433;
wire            n6434;
wire      [7:0] n6435;
wire            n6436;
wire      [7:0] n6437;
wire            n6438;
wire      [7:0] n6439;
wire            n644;
wire            n6440;
wire      [7:0] n6441;
wire            n6442;
wire      [7:0] n6443;
wire            n6444;
wire      [7:0] n6445;
wire            n6446;
wire      [7:0] n6447;
wire            n6448;
wire      [7:0] n6449;
wire            n6450;
wire      [7:0] n6451;
wire            n6452;
wire      [7:0] n6453;
wire            n6454;
wire      [7:0] n6455;
wire            n6456;
wire      [7:0] n6457;
wire            n6458;
wire      [7:0] n6459;
wire      [7:0] n646;
wire            n6460;
wire      [7:0] n6461;
wire            n6462;
wire      [7:0] n6463;
wire            n6464;
wire      [7:0] n6465;
wire            n6466;
wire      [7:0] n6467;
wire            n6468;
wire      [7:0] n6469;
wire            n647;
wire            n6470;
wire      [7:0] n6471;
wire            n6472;
wire      [7:0] n6473;
wire            n6474;
wire      [7:0] n6475;
wire            n6476;
wire      [7:0] n6477;
wire            n6478;
wire      [7:0] n6479;
wire            n6480;
wire      [7:0] n6481;
wire            n6482;
wire      [7:0] n6483;
wire            n6484;
wire      [7:0] n6485;
wire            n6486;
wire      [7:0] n6487;
wire            n6488;
wire      [7:0] n6489;
wire      [7:0] n649;
wire            n6490;
wire      [7:0] n6491;
wire            n6492;
wire      [7:0] n6493;
wire            n6494;
wire      [7:0] n6495;
wire            n6496;
wire      [7:0] n6497;
wire            n6498;
wire      [7:0] n6499;
wire            n6500;
wire      [7:0] n6501;
wire            n6502;
wire      [7:0] n6503;
wire            n6504;
wire      [7:0] n6505;
wire            n6506;
wire      [7:0] n6507;
wire            n6508;
wire      [7:0] n6509;
wire            n651;
wire            n6510;
wire      [7:0] n6511;
wire            n6512;
wire      [7:0] n6513;
wire            n6514;
wire      [7:0] n6515;
wire            n6516;
wire      [7:0] n6517;
wire            n6518;
wire      [7:0] n6519;
wire            n6520;
wire      [7:0] n6521;
wire            n6522;
wire      [7:0] n6523;
wire            n6524;
wire      [7:0] n6525;
wire            n6526;
wire      [7:0] n6527;
wire            n6528;
wire      [7:0] n6529;
wire      [7:0] n653;
wire            n6530;
wire      [7:0] n6531;
wire            n6532;
wire      [7:0] n6533;
wire            n6534;
wire      [7:0] n6535;
wire            n6536;
wire      [7:0] n6537;
wire            n6538;
wire      [7:0] n6539;
wire            n654;
wire            n6540;
wire      [7:0] n6541;
wire            n6542;
wire      [7:0] n6543;
wire            n6544;
wire      [7:0] n6545;
wire            n6546;
wire      [7:0] n6547;
wire            n6548;
wire      [7:0] n6549;
wire            n6550;
wire      [7:0] n6551;
wire            n6552;
wire      [7:0] n6553;
wire            n6554;
wire      [7:0] n6555;
wire            n6556;
wire      [7:0] n6557;
wire            n6558;
wire      [7:0] n6559;
wire      [7:0] n656;
wire            n6560;
wire      [7:0] n6561;
wire            n6562;
wire      [7:0] n6563;
wire            n6564;
wire      [7:0] n6565;
wire            n6566;
wire      [7:0] n6567;
wire            n6568;
wire      [7:0] n6569;
wire            n657;
wire            n6570;
wire      [7:0] n6571;
wire            n6572;
wire      [7:0] n6573;
wire            n6574;
wire      [7:0] n6575;
wire            n6576;
wire      [7:0] n6577;
wire            n6578;
wire      [7:0] n6579;
wire      [7:0] n658;
wire            n6580;
wire      [7:0] n6581;
wire            n6582;
wire      [7:0] n6583;
wire            n6584;
wire      [7:0] n6585;
wire            n6586;
wire      [7:0] n6587;
wire            n6588;
wire      [7:0] n6589;
wire            n659;
wire            n6590;
wire      [7:0] n6591;
wire            n6592;
wire      [7:0] n6593;
wire            n6594;
wire      [7:0] n6595;
wire            n6596;
wire      [7:0] n6597;
wire            n6598;
wire      [7:0] n6599;
wire      [7:0] n66;
wire            n6600;
wire      [7:0] n6601;
wire            n6602;
wire      [7:0] n6603;
wire            n6604;
wire      [7:0] n6605;
wire            n6606;
wire      [7:0] n6607;
wire            n6608;
wire      [7:0] n6609;
wire      [7:0] n661;
wire            n6610;
wire      [7:0] n6611;
wire            n6612;
wire      [7:0] n6613;
wire            n6614;
wire      [7:0] n6615;
wire            n6616;
wire      [7:0] n6617;
wire            n6618;
wire      [7:0] n6619;
wire            n662;
wire            n6620;
wire      [7:0] n6621;
wire            n6622;
wire      [7:0] n6623;
wire            n6624;
wire      [7:0] n6625;
wire            n6626;
wire      [7:0] n6627;
wire            n6628;
wire      [7:0] n6629;
wire      [7:0] n663;
wire            n6630;
wire      [7:0] n6631;
wire            n6632;
wire      [7:0] n6633;
wire            n6634;
wire      [7:0] n6635;
wire            n6636;
wire      [7:0] n6637;
wire            n6638;
wire      [7:0] n6639;
wire            n664;
wire            n6640;
wire      [7:0] n6641;
wire            n6642;
wire      [7:0] n6643;
wire            n6644;
wire      [7:0] n6645;
wire            n6646;
wire      [7:0] n6647;
wire            n6648;
wire      [7:0] n6649;
wire      [7:0] n665;
wire            n6650;
wire      [7:0] n6651;
wire            n6652;
wire      [7:0] n6653;
wire            n6654;
wire      [7:0] n6655;
wire            n6656;
wire      [7:0] n6657;
wire            n6658;
wire      [7:0] n6659;
wire            n666;
wire            n6660;
wire      [7:0] n6661;
wire            n6662;
wire      [7:0] n6663;
wire            n6664;
wire      [7:0] n6665;
wire            n6666;
wire      [7:0] n6667;
wire            n6668;
wire      [7:0] n6669;
wire      [7:0] n667;
wire            n6670;
wire      [7:0] n6671;
wire            n6672;
wire      [7:0] n6673;
wire            n6674;
wire      [7:0] n6675;
wire            n6676;
wire      [7:0] n6677;
wire            n6678;
wire      [7:0] n6679;
wire            n668;
wire            n6680;
wire      [7:0] n6681;
wire            n6682;
wire      [7:0] n6683;
wire            n6684;
wire      [7:0] n6685;
wire            n6686;
wire      [7:0] n6687;
wire            n6688;
wire      [7:0] n6689;
wire            n6690;
wire      [7:0] n6691;
wire            n6692;
wire      [7:0] n6693;
wire            n6694;
wire      [7:0] n6695;
wire            n6696;
wire      [7:0] n6697;
wire            n6698;
wire      [7:0] n6699;
wire      [7:0] n670;
wire            n6700;
wire      [7:0] n6701;
wire            n6702;
wire      [7:0] n6703;
wire            n6704;
wire      [7:0] n6705;
wire            n6706;
wire      [7:0] n6707;
wire            n6708;
wire      [7:0] n6709;
wire            n671;
wire            n6710;
wire      [7:0] n6711;
wire            n6712;
wire      [7:0] n6713;
wire            n6714;
wire      [7:0] n6715;
wire            n6716;
wire      [7:0] n6717;
wire            n6718;
wire      [7:0] n6719;
wire            n6720;
wire      [7:0] n6721;
wire            n6722;
wire      [7:0] n6723;
wire            n6724;
wire      [7:0] n6725;
wire            n6726;
wire      [7:0] n6727;
wire            n6728;
wire      [7:0] n6729;
wire      [7:0] n673;
wire            n6730;
wire      [7:0] n6731;
wire            n6732;
wire      [7:0] n6733;
wire            n6734;
wire      [7:0] n6735;
wire            n6736;
wire      [7:0] n6737;
wire            n6738;
wire      [7:0] n6739;
wire            n674;
wire            n6740;
wire      [7:0] n6741;
wire            n6742;
wire      [7:0] n6743;
wire            n6744;
wire      [7:0] n6745;
wire            n6746;
wire      [7:0] n6747;
wire            n6748;
wire      [7:0] n6749;
wire      [7:0] n675;
wire            n6750;
wire      [7:0] n6751;
wire            n6752;
wire      [7:0] n6753;
wire            n6754;
wire      [7:0] n6755;
wire            n6756;
wire      [7:0] n6757;
wire            n6758;
wire      [7:0] n6759;
wire            n676;
wire            n6760;
wire      [7:0] n6761;
wire            n6762;
wire      [7:0] n6763;
wire            n6764;
wire      [7:0] n6765;
wire            n6766;
wire      [7:0] n6767;
wire            n6768;
wire      [7:0] n6769;
wire      [7:0] n677;
wire            n6770;
wire      [7:0] n6771;
wire            n6772;
wire      [7:0] n6773;
wire            n6774;
wire      [7:0] n6775;
wire            n6776;
wire      [7:0] n6777;
wire            n6778;
wire      [7:0] n6779;
wire            n678;
wire            n6780;
wire      [7:0] n6781;
wire            n6782;
wire      [7:0] n6783;
wire            n6784;
wire      [7:0] n6785;
wire            n6786;
wire      [7:0] n6787;
wire            n6788;
wire      [7:0] n6789;
wire      [7:0] n679;
wire            n6790;
wire      [7:0] n6791;
wire            n6792;
wire      [7:0] n6793;
wire            n6794;
wire      [7:0] n6795;
wire            n6796;
wire      [7:0] n6797;
wire            n6798;
wire      [7:0] n6799;
wire            n68;
wire            n680;
wire            n6800;
wire      [7:0] n6801;
wire            n6802;
wire      [7:0] n6803;
wire            n6804;
wire      [7:0] n6805;
wire            n6806;
wire      [7:0] n6807;
wire            n6808;
wire      [7:0] n6809;
wire      [7:0] n681;
wire            n6810;
wire      [7:0] n6811;
wire            n6812;
wire      [7:0] n6813;
wire            n6814;
wire      [7:0] n6815;
wire            n6816;
wire      [7:0] n6817;
wire            n6818;
wire      [7:0] n6819;
wire            n682;
wire            n6820;
wire      [7:0] n6821;
wire            n6822;
wire      [7:0] n6823;
wire            n6824;
wire      [7:0] n6825;
wire            n6826;
wire      [7:0] n6827;
wire            n6828;
wire      [7:0] n6829;
wire      [7:0] n683;
wire            n6830;
wire      [7:0] n6831;
wire            n6832;
wire      [7:0] n6833;
wire            n6834;
wire      [7:0] n6835;
wire            n6836;
wire      [7:0] n6837;
wire            n6838;
wire      [7:0] n6839;
wire            n684;
wire            n6840;
wire      [7:0] n6841;
wire            n6842;
wire      [7:0] n6843;
wire            n6844;
wire      [7:0] n6845;
wire            n6846;
wire      [7:0] n6847;
wire            n6848;
wire      [7:0] n6849;
wire      [7:0] n685;
wire            n6850;
wire      [7:0] n6851;
wire            n6852;
wire      [7:0] n6853;
wire            n6854;
wire      [7:0] n6855;
wire            n6856;
wire      [7:0] n6857;
wire            n6858;
wire      [7:0] n6859;
wire            n686;
wire            n6860;
wire      [7:0] n6861;
wire            n6862;
wire      [7:0] n6863;
wire            n6864;
wire      [7:0] n6865;
wire            n6866;
wire      [7:0] n6867;
wire            n6868;
wire      [7:0] n6869;
wire      [7:0] n687;
wire            n6870;
wire      [7:0] n6871;
wire            n6872;
wire      [7:0] n6873;
wire            n6874;
wire      [7:0] n6875;
wire            n6876;
wire      [7:0] n6877;
wire            n6878;
wire      [7:0] n6879;
wire            n688;
wire            n6880;
wire      [7:0] n6881;
wire            n6882;
wire      [7:0] n6883;
wire            n6884;
wire      [7:0] n6885;
wire            n6886;
wire      [7:0] n6887;
wire            n6888;
wire      [7:0] n6889;
wire      [7:0] n689;
wire            n6890;
wire      [7:0] n6891;
wire            n6892;
wire      [7:0] n6893;
wire            n6894;
wire      [7:0] n6895;
wire            n6896;
wire      [7:0] n6897;
wire            n6898;
wire      [7:0] n6899;
wire            n690;
wire            n6900;
wire      [7:0] n6901;
wire            n6902;
wire      [7:0] n6903;
wire            n6904;
wire      [7:0] n6905;
wire            n6906;
wire      [7:0] n6907;
wire            n6908;
wire      [7:0] n6909;
wire      [7:0] n691;
wire            n6910;
wire      [7:0] n6911;
wire            n6912;
wire      [7:0] n6913;
wire            n6914;
wire      [7:0] n6915;
wire            n6916;
wire      [7:0] n6917;
wire            n6918;
wire      [7:0] n6919;
wire            n692;
wire            n6920;
wire      [7:0] n6921;
wire            n6922;
wire      [7:0] n6923;
wire            n6924;
wire      [7:0] n6925;
wire            n6926;
wire      [7:0] n6927;
wire            n6928;
wire      [7:0] n6929;
wire      [7:0] n693;
wire            n6930;
wire      [7:0] n6931;
wire            n6932;
wire      [7:0] n6933;
wire            n6934;
wire      [7:0] n6935;
wire            n6936;
wire      [7:0] n6937;
wire            n6938;
wire      [7:0] n6939;
wire            n694;
wire            n6940;
wire      [7:0] n6941;
wire      [7:0] n6942;
wire      [7:0] n6943;
wire      [7:0] n6944;
wire      [7:0] n6945;
wire      [7:0] n6946;
wire      [7:0] n6947;
wire      [7:0] n6948;
wire      [7:0] n6949;
wire      [7:0] n695;
wire      [7:0] n6950;
wire      [7:0] n6951;
wire      [7:0] n6952;
wire      [7:0] n6953;
wire      [7:0] n6954;
wire      [7:0] n6955;
wire      [7:0] n6956;
wire      [7:0] n6957;
wire      [7:0] n6958;
wire      [7:0] n6959;
wire      [7:0] n6960;
wire      [7:0] n6961;
wire      [7:0] n6962;
wire      [7:0] n6963;
wire      [7:0] n6964;
wire      [7:0] n6965;
wire      [7:0] n6966;
wire      [7:0] n6967;
wire      [7:0] n6968;
wire      [7:0] n6969;
wire            n697;
wire      [7:0] n6970;
wire      [7:0] n6971;
wire      [7:0] n6972;
wire      [7:0] n6973;
wire      [7:0] n6974;
wire      [7:0] n6975;
wire      [7:0] n6976;
wire      [7:0] n6977;
wire      [7:0] n6978;
wire      [7:0] n6979;
wire      [7:0] n698;
wire      [7:0] n6980;
wire      [7:0] n6981;
wire      [7:0] n6982;
wire      [7:0] n6983;
wire      [7:0] n6984;
wire      [7:0] n6985;
wire      [7:0] n6986;
wire      [7:0] n6987;
wire      [7:0] n6988;
wire      [7:0] n6989;
wire            n699;
wire      [7:0] n6990;
wire      [7:0] n6991;
wire      [7:0] n6992;
wire      [7:0] n6993;
wire      [7:0] n6994;
wire      [7:0] n6995;
wire      [7:0] n6996;
wire      [7:0] n6997;
wire      [7:0] n6998;
wire      [7:0] n6999;
wire      [7:0] n70;
wire      [7:0] n700;
wire      [7:0] n7000;
wire      [7:0] n7001;
wire      [7:0] n7002;
wire      [7:0] n7003;
wire      [7:0] n7004;
wire      [7:0] n7005;
wire      [7:0] n7006;
wire      [7:0] n7007;
wire      [7:0] n7008;
wire      [7:0] n7009;
wire            n701;
wire      [7:0] n7010;
wire      [7:0] n7011;
wire      [7:0] n7012;
wire      [7:0] n7013;
wire      [7:0] n7014;
wire      [7:0] n7015;
wire      [7:0] n7016;
wire      [7:0] n7017;
wire      [7:0] n7018;
wire      [7:0] n7019;
wire      [7:0] n702;
wire      [7:0] n7020;
wire      [7:0] n7021;
wire      [7:0] n7022;
wire      [7:0] n7023;
wire      [7:0] n7024;
wire      [7:0] n7025;
wire      [7:0] n7026;
wire      [7:0] n7027;
wire      [7:0] n7028;
wire      [7:0] n7029;
wire            n703;
wire      [7:0] n7030;
wire      [7:0] n7031;
wire      [7:0] n7032;
wire      [7:0] n7033;
wire      [7:0] n7034;
wire      [7:0] n7035;
wire      [7:0] n7036;
wire      [7:0] n7037;
wire      [7:0] n7038;
wire      [7:0] n7039;
wire      [7:0] n704;
wire      [7:0] n7040;
wire      [7:0] n7041;
wire      [7:0] n7042;
wire      [7:0] n7043;
wire      [7:0] n7044;
wire      [7:0] n7045;
wire      [7:0] n7046;
wire      [7:0] n7047;
wire      [7:0] n7048;
wire      [7:0] n7049;
wire      [7:0] n7050;
wire      [7:0] n7051;
wire      [7:0] n7052;
wire      [7:0] n7053;
wire      [7:0] n7054;
wire      [7:0] n7055;
wire      [7:0] n7056;
wire      [7:0] n7057;
wire      [7:0] n7058;
wire      [7:0] n7059;
wire            n706;
wire      [7:0] n7060;
wire      [7:0] n7061;
wire      [7:0] n7062;
wire      [7:0] n7063;
wire      [7:0] n7064;
wire      [7:0] n7065;
wire      [7:0] n7066;
wire      [7:0] n7067;
wire      [7:0] n7068;
wire      [7:0] n7069;
wire      [7:0] n707;
wire      [7:0] n7070;
wire      [7:0] n7071;
wire      [7:0] n7072;
wire      [7:0] n7073;
wire      [7:0] n7074;
wire      [7:0] n7075;
wire      [7:0] n7076;
wire      [7:0] n7077;
wire      [7:0] n7078;
wire      [7:0] n7079;
wire            n708;
wire      [7:0] n7080;
wire      [7:0] n7081;
wire      [7:0] n7082;
wire      [7:0] n7083;
wire      [7:0] n7084;
wire      [7:0] n7085;
wire      [7:0] n7086;
wire      [7:0] n7087;
wire      [7:0] n7088;
wire      [7:0] n7089;
wire      [7:0] n709;
wire      [7:0] n7090;
wire      [7:0] n7091;
wire      [7:0] n7092;
wire      [7:0] n7093;
wire      [7:0] n7094;
wire      [7:0] n7095;
wire      [7:0] n7096;
wire      [7:0] n7097;
wire      [7:0] n7098;
wire      [7:0] n7099;
wire            n710;
wire      [7:0] n7100;
wire      [7:0] n7101;
wire      [7:0] n7102;
wire      [7:0] n7103;
wire      [7:0] n7104;
wire      [7:0] n7105;
wire      [7:0] n7106;
wire      [7:0] n7107;
wire      [7:0] n7108;
wire      [7:0] n7109;
wire      [7:0] n711;
wire      [7:0] n7110;
wire      [7:0] n7111;
wire      [7:0] n7112;
wire      [7:0] n7113;
wire      [7:0] n7114;
wire      [7:0] n7115;
wire      [7:0] n7116;
wire      [7:0] n7117;
wire      [7:0] n7118;
wire      [7:0] n7119;
wire            n712;
wire      [7:0] n7120;
wire      [7:0] n7121;
wire      [7:0] n7122;
wire      [7:0] n7123;
wire      [7:0] n7124;
wire      [7:0] n7125;
wire      [7:0] n7126;
wire      [7:0] n7127;
wire      [7:0] n7128;
wire      [7:0] n7129;
wire      [7:0] n713;
wire      [7:0] n7130;
wire      [7:0] n7131;
wire      [7:0] n7132;
wire      [7:0] n7133;
wire      [7:0] n7134;
wire      [7:0] n7135;
wire      [7:0] n7136;
wire      [7:0] n7137;
wire      [7:0] n7138;
wire      [7:0] n7139;
wire            n714;
wire      [7:0] n7140;
wire      [7:0] n7141;
wire      [7:0] n7142;
wire      [7:0] n7143;
wire      [7:0] n7144;
wire      [7:0] n7145;
wire      [7:0] n7146;
wire      [7:0] n7147;
wire      [7:0] n7148;
wire      [7:0] n7149;
wire      [7:0] n715;
wire      [7:0] n7150;
wire      [7:0] n7151;
wire      [7:0] n7152;
wire      [7:0] n7153;
wire      [7:0] n7154;
wire      [7:0] n7155;
wire      [7:0] n7156;
wire      [7:0] n7157;
wire      [7:0] n7158;
wire      [7:0] n7159;
wire            n716;
wire      [7:0] n7160;
wire      [7:0] n7161;
wire      [7:0] n7162;
wire      [7:0] n7163;
wire      [7:0] n7164;
wire      [7:0] n7165;
wire      [7:0] n7166;
wire      [7:0] n7167;
wire      [7:0] n7168;
wire      [7:0] n7169;
wire      [7:0] n717;
wire      [7:0] n7170;
wire      [7:0] n7171;
wire      [7:0] n7172;
wire      [7:0] n7173;
wire      [7:0] n7174;
wire      [7:0] n7175;
wire      [7:0] n7176;
wire      [7:0] n7177;
wire      [7:0] n7178;
wire      [7:0] n7179;
wire            n718;
wire      [7:0] n7180;
wire      [7:0] n7181;
wire      [7:0] n7182;
wire      [7:0] n7183;
wire      [7:0] n7184;
wire      [7:0] n7185;
wire      [7:0] n7186;
wire      [7:0] n7187;
wire      [7:0] n7188;
wire      [7:0] n7189;
wire      [7:0] n719;
wire      [7:0] n7190;
wire      [7:0] n7191;
wire      [7:0] n7192;
wire      [7:0] n7193;
wire      [7:0] n7194;
wire      [7:0] n7195;
wire      [7:0] n7196;
wire      [7:0] n7197;
wire            n7198;
wire      [7:0] n7199;
wire            n72;
wire            n720;
wire            n7200;
wire      [7:0] n7201;
wire            n7202;
wire      [7:0] n7203;
wire            n7204;
wire      [7:0] n7205;
wire            n7206;
wire      [7:0] n7207;
wire            n7208;
wire      [7:0] n7209;
wire      [7:0] n721;
wire            n7210;
wire      [7:0] n7211;
wire            n7212;
wire      [7:0] n7213;
wire            n7214;
wire      [7:0] n7215;
wire            n7216;
wire      [7:0] n7217;
wire            n7218;
wire      [7:0] n7219;
wire            n722;
wire            n7220;
wire      [7:0] n7221;
wire            n7222;
wire      [7:0] n7223;
wire            n7224;
wire      [7:0] n7225;
wire            n7226;
wire      [7:0] n7227;
wire            n7228;
wire      [7:0] n7229;
wire      [7:0] n723;
wire            n7230;
wire      [7:0] n7231;
wire            n7232;
wire      [7:0] n7233;
wire            n7234;
wire      [7:0] n7235;
wire            n7236;
wire      [7:0] n7237;
wire            n7238;
wire      [7:0] n7239;
wire            n724;
wire            n7240;
wire      [7:0] n7241;
wire            n7242;
wire      [7:0] n7243;
wire            n7244;
wire      [7:0] n7245;
wire            n7246;
wire      [7:0] n7247;
wire            n7248;
wire      [7:0] n7249;
wire      [7:0] n725;
wire            n7250;
wire      [7:0] n7251;
wire            n7252;
wire      [7:0] n7253;
wire            n7254;
wire      [7:0] n7255;
wire            n7256;
wire      [7:0] n7257;
wire            n7258;
wire      [7:0] n7259;
wire            n726;
wire            n7260;
wire      [7:0] n7261;
wire            n7262;
wire      [7:0] n7263;
wire            n7264;
wire      [7:0] n7265;
wire            n7266;
wire      [7:0] n7267;
wire            n7268;
wire      [7:0] n7269;
wire      [7:0] n727;
wire            n7270;
wire      [7:0] n7271;
wire            n7272;
wire      [7:0] n7273;
wire            n7274;
wire      [7:0] n7275;
wire            n7276;
wire      [7:0] n7277;
wire            n7278;
wire      [7:0] n7279;
wire            n728;
wire            n7280;
wire      [7:0] n7281;
wire            n7282;
wire      [7:0] n7283;
wire            n7284;
wire      [7:0] n7285;
wire            n7286;
wire      [7:0] n7287;
wire            n7288;
wire      [7:0] n7289;
wire      [7:0] n729;
wire            n7290;
wire      [7:0] n7291;
wire            n7292;
wire      [7:0] n7293;
wire            n7294;
wire      [7:0] n7295;
wire            n7296;
wire      [7:0] n7297;
wire            n7298;
wire      [7:0] n7299;
wire            n730;
wire            n7300;
wire      [7:0] n7301;
wire            n7302;
wire      [7:0] n7303;
wire            n7304;
wire      [7:0] n7305;
wire            n7306;
wire      [7:0] n7307;
wire            n7308;
wire      [7:0] n7309;
wire      [7:0] n731;
wire            n7310;
wire      [7:0] n7311;
wire            n7312;
wire      [7:0] n7313;
wire            n7314;
wire      [7:0] n7315;
wire            n7316;
wire      [7:0] n7317;
wire            n7318;
wire      [7:0] n7319;
wire            n732;
wire            n7320;
wire      [7:0] n7321;
wire            n7322;
wire      [7:0] n7323;
wire            n7324;
wire      [7:0] n7325;
wire            n7326;
wire      [7:0] n7327;
wire            n7328;
wire      [7:0] n7329;
wire      [7:0] n733;
wire            n7330;
wire      [7:0] n7331;
wire            n7332;
wire      [7:0] n7333;
wire            n7334;
wire      [7:0] n7335;
wire            n7336;
wire      [7:0] n7337;
wire            n7338;
wire      [7:0] n7339;
wire            n734;
wire            n7340;
wire      [7:0] n7341;
wire            n7342;
wire      [7:0] n7343;
wire            n7344;
wire      [7:0] n7345;
wire            n7346;
wire      [7:0] n7347;
wire            n7348;
wire      [7:0] n7349;
wire      [7:0] n735;
wire            n7350;
wire      [7:0] n7351;
wire            n7352;
wire      [7:0] n7353;
wire            n7354;
wire      [7:0] n7355;
wire            n7356;
wire      [7:0] n7357;
wire            n7358;
wire      [7:0] n7359;
wire            n736;
wire            n7360;
wire      [7:0] n7361;
wire            n7362;
wire      [7:0] n7363;
wire            n7364;
wire      [7:0] n7365;
wire            n7366;
wire      [7:0] n7367;
wire            n7368;
wire      [7:0] n7369;
wire      [7:0] n737;
wire            n7370;
wire      [7:0] n7371;
wire            n7372;
wire      [7:0] n7373;
wire            n7374;
wire      [7:0] n7375;
wire            n7376;
wire      [7:0] n7377;
wire            n7378;
wire      [7:0] n7379;
wire            n738;
wire            n7380;
wire      [7:0] n7381;
wire            n7382;
wire      [7:0] n7383;
wire            n7384;
wire      [7:0] n7385;
wire            n7386;
wire      [7:0] n7387;
wire            n7388;
wire      [7:0] n7389;
wire      [7:0] n739;
wire            n7390;
wire      [7:0] n7391;
wire            n7392;
wire      [7:0] n7393;
wire            n7394;
wire      [7:0] n7395;
wire            n7396;
wire      [7:0] n7397;
wire            n7398;
wire      [7:0] n7399;
wire      [7:0] n74;
wire            n740;
wire            n7400;
wire      [7:0] n7401;
wire            n7402;
wire      [7:0] n7403;
wire            n7404;
wire      [7:0] n7405;
wire            n7406;
wire      [7:0] n7407;
wire            n7408;
wire      [7:0] n7409;
wire      [7:0] n741;
wire            n7410;
wire      [7:0] n7411;
wire            n7412;
wire      [7:0] n7413;
wire            n7414;
wire      [7:0] n7415;
wire            n7416;
wire      [7:0] n7417;
wire            n7418;
wire      [7:0] n7419;
wire            n742;
wire            n7420;
wire      [7:0] n7421;
wire            n7422;
wire      [7:0] n7423;
wire            n7424;
wire      [7:0] n7425;
wire            n7426;
wire      [7:0] n7427;
wire            n7428;
wire      [7:0] n7429;
wire      [7:0] n743;
wire            n7430;
wire      [7:0] n7431;
wire            n7432;
wire      [7:0] n7433;
wire            n7434;
wire      [7:0] n7435;
wire            n7436;
wire      [7:0] n7437;
wire            n7438;
wire      [7:0] n7439;
wire            n744;
wire            n7440;
wire      [7:0] n7441;
wire            n7442;
wire      [7:0] n7443;
wire            n7444;
wire      [7:0] n7445;
wire            n7446;
wire      [7:0] n7447;
wire            n7448;
wire      [7:0] n7449;
wire      [7:0] n745;
wire            n7450;
wire      [7:0] n7451;
wire            n7452;
wire      [7:0] n7453;
wire            n7454;
wire      [7:0] n7455;
wire            n7456;
wire      [7:0] n7457;
wire            n7458;
wire      [7:0] n7459;
wire            n746;
wire            n7460;
wire      [7:0] n7461;
wire            n7462;
wire      [7:0] n7463;
wire            n7464;
wire      [7:0] n7465;
wire            n7466;
wire      [7:0] n7467;
wire            n7468;
wire      [7:0] n7469;
wire      [7:0] n747;
wire            n7470;
wire      [7:0] n7471;
wire            n7472;
wire      [7:0] n7473;
wire            n7474;
wire      [7:0] n7475;
wire            n7476;
wire      [7:0] n7477;
wire            n7478;
wire      [7:0] n7479;
wire            n748;
wire            n7480;
wire      [7:0] n7481;
wire            n7482;
wire      [7:0] n7483;
wire            n7484;
wire      [7:0] n7485;
wire            n7486;
wire      [7:0] n7487;
wire            n7488;
wire      [7:0] n7489;
wire      [7:0] n749;
wire            n7490;
wire      [7:0] n7491;
wire            n7492;
wire      [7:0] n7493;
wire            n7494;
wire      [7:0] n7495;
wire            n7496;
wire      [7:0] n7497;
wire            n7498;
wire      [7:0] n7499;
wire            n750;
wire            n7500;
wire      [7:0] n7501;
wire            n7502;
wire      [7:0] n7503;
wire            n7504;
wire      [7:0] n7505;
wire            n7506;
wire      [7:0] n7507;
wire            n7508;
wire      [7:0] n7509;
wire            n7510;
wire      [7:0] n7511;
wire            n7512;
wire      [7:0] n7513;
wire            n7514;
wire      [7:0] n7515;
wire            n7516;
wire      [7:0] n7517;
wire            n7518;
wire      [7:0] n7519;
wire      [7:0] n752;
wire            n7520;
wire      [7:0] n7521;
wire            n7522;
wire      [7:0] n7523;
wire            n7524;
wire      [7:0] n7525;
wire            n7526;
wire      [7:0] n7527;
wire            n7528;
wire      [7:0] n7529;
wire            n753;
wire            n7530;
wire      [7:0] n7531;
wire            n7532;
wire      [7:0] n7533;
wire            n7534;
wire      [7:0] n7535;
wire            n7536;
wire      [7:0] n7537;
wire            n7538;
wire      [7:0] n7539;
wire      [7:0] n754;
wire            n7540;
wire      [7:0] n7541;
wire            n7542;
wire      [7:0] n7543;
wire            n7544;
wire      [7:0] n7545;
wire            n7546;
wire      [7:0] n7547;
wire            n7548;
wire      [7:0] n7549;
wire            n755;
wire            n7550;
wire      [7:0] n7551;
wire            n7552;
wire      [7:0] n7553;
wire            n7554;
wire      [7:0] n7555;
wire            n7556;
wire      [7:0] n7557;
wire            n7558;
wire      [7:0] n7559;
wire      [7:0] n756;
wire            n7560;
wire      [7:0] n7561;
wire            n7562;
wire      [7:0] n7563;
wire            n7564;
wire      [7:0] n7565;
wire            n7566;
wire      [7:0] n7567;
wire            n7568;
wire      [7:0] n7569;
wire            n757;
wire            n7570;
wire      [7:0] n7571;
wire            n7572;
wire      [7:0] n7573;
wire            n7574;
wire      [7:0] n7575;
wire            n7576;
wire      [7:0] n7577;
wire            n7578;
wire      [7:0] n7579;
wire      [7:0] n758;
wire            n7580;
wire      [7:0] n7581;
wire            n7582;
wire      [7:0] n7583;
wire            n7584;
wire      [7:0] n7585;
wire            n7586;
wire      [7:0] n7587;
wire            n7588;
wire      [7:0] n7589;
wire            n759;
wire            n7590;
wire      [7:0] n7591;
wire            n7592;
wire      [7:0] n7593;
wire            n7594;
wire      [7:0] n7595;
wire            n7596;
wire      [7:0] n7597;
wire            n7598;
wire      [7:0] n7599;
wire            n76;
wire      [7:0] n760;
wire            n7600;
wire      [7:0] n7601;
wire            n7602;
wire      [7:0] n7603;
wire            n7604;
wire      [7:0] n7605;
wire            n7606;
wire      [7:0] n7607;
wire            n7608;
wire      [7:0] n7609;
wire            n761;
wire            n7610;
wire      [7:0] n7611;
wire            n7612;
wire      [7:0] n7613;
wire            n7614;
wire      [7:0] n7615;
wire            n7616;
wire      [7:0] n7617;
wire            n7618;
wire      [7:0] n7619;
wire      [7:0] n762;
wire            n7620;
wire      [7:0] n7621;
wire            n7622;
wire      [7:0] n7623;
wire            n7624;
wire      [7:0] n7625;
wire            n7626;
wire      [7:0] n7627;
wire            n7628;
wire      [7:0] n7629;
wire            n763;
wire            n7630;
wire      [7:0] n7631;
wire            n7632;
wire      [7:0] n7633;
wire            n7634;
wire      [7:0] n7635;
wire            n7636;
wire      [7:0] n7637;
wire            n7638;
wire      [7:0] n7639;
wire      [7:0] n764;
wire            n7640;
wire      [7:0] n7641;
wire            n7642;
wire      [7:0] n7643;
wire            n7644;
wire      [7:0] n7645;
wire            n7646;
wire      [7:0] n7647;
wire            n7648;
wire      [7:0] n7649;
wire            n765;
wire            n7650;
wire      [7:0] n7651;
wire            n7652;
wire      [7:0] n7653;
wire            n7654;
wire      [7:0] n7655;
wire            n7656;
wire      [7:0] n7657;
wire            n7658;
wire      [7:0] n7659;
wire      [7:0] n766;
wire            n7660;
wire      [7:0] n7661;
wire            n7662;
wire      [7:0] n7663;
wire            n7664;
wire      [7:0] n7665;
wire            n7666;
wire      [7:0] n7667;
wire            n7668;
wire      [7:0] n7669;
wire            n767;
wire            n7670;
wire      [7:0] n7671;
wire            n7672;
wire      [7:0] n7673;
wire            n7674;
wire      [7:0] n7675;
wire            n7676;
wire      [7:0] n7677;
wire            n7678;
wire      [7:0] n7679;
wire      [7:0] n768;
wire            n7680;
wire      [7:0] n7681;
wire            n7682;
wire      [7:0] n7683;
wire            n7684;
wire      [7:0] n7685;
wire            n7686;
wire      [7:0] n7687;
wire            n7688;
wire      [7:0] n7689;
wire            n769;
wire            n7690;
wire      [7:0] n7691;
wire            n7692;
wire      [7:0] n7693;
wire            n7694;
wire      [7:0] n7695;
wire            n7696;
wire      [7:0] n7697;
wire            n7698;
wire      [7:0] n7699;
wire      [7:0] n770;
wire            n7700;
wire      [7:0] n7701;
wire            n7702;
wire      [7:0] n7703;
wire            n7704;
wire      [7:0] n7705;
wire            n7706;
wire      [7:0] n7707;
wire            n7708;
wire      [7:0] n7709;
wire      [7:0] n771;
wire      [7:0] n7710;
wire      [7:0] n7711;
wire      [7:0] n7712;
wire      [7:0] n7713;
wire      [7:0] n7714;
wire      [7:0] n7715;
wire      [7:0] n7716;
wire      [7:0] n7717;
wire      [7:0] n7718;
wire      [7:0] n7719;
wire      [7:0] n772;
wire      [7:0] n7720;
wire      [7:0] n7721;
wire      [7:0] n7722;
wire      [7:0] n7723;
wire      [7:0] n7724;
wire      [7:0] n7725;
wire      [7:0] n7726;
wire      [7:0] n7727;
wire      [7:0] n7728;
wire      [7:0] n7729;
wire      [7:0] n773;
wire      [7:0] n7730;
wire      [7:0] n7731;
wire      [7:0] n7732;
wire      [7:0] n7733;
wire      [7:0] n7734;
wire      [7:0] n7735;
wire      [7:0] n7736;
wire      [7:0] n7737;
wire      [7:0] n7738;
wire      [7:0] n7739;
wire      [7:0] n774;
wire      [7:0] n7740;
wire      [7:0] n7741;
wire      [7:0] n7742;
wire      [7:0] n7743;
wire      [7:0] n7744;
wire      [7:0] n7745;
wire      [7:0] n7746;
wire      [7:0] n7747;
wire      [7:0] n7748;
wire      [7:0] n7749;
wire      [7:0] n775;
wire      [7:0] n7750;
wire      [7:0] n7751;
wire      [7:0] n7752;
wire      [7:0] n7753;
wire      [7:0] n7754;
wire      [7:0] n7755;
wire      [7:0] n7756;
wire      [7:0] n7757;
wire      [7:0] n7758;
wire      [7:0] n7759;
wire      [7:0] n776;
wire      [7:0] n7760;
wire      [7:0] n7761;
wire      [7:0] n7762;
wire      [7:0] n7763;
wire      [7:0] n7764;
wire      [7:0] n7765;
wire      [7:0] n7766;
wire      [7:0] n7767;
wire      [7:0] n7768;
wire      [7:0] n7769;
wire      [7:0] n777;
wire      [7:0] n7770;
wire      [7:0] n7771;
wire      [7:0] n7772;
wire      [7:0] n7773;
wire      [7:0] n7774;
wire      [7:0] n7775;
wire      [7:0] n7776;
wire      [7:0] n7777;
wire      [7:0] n7778;
wire      [7:0] n7779;
wire      [7:0] n778;
wire      [7:0] n7780;
wire      [7:0] n7781;
wire      [7:0] n7782;
wire      [7:0] n7783;
wire      [7:0] n7784;
wire      [7:0] n7785;
wire      [7:0] n7786;
wire      [7:0] n7787;
wire      [7:0] n7788;
wire      [7:0] n7789;
wire      [7:0] n779;
wire      [7:0] n7790;
wire      [7:0] n7791;
wire      [7:0] n7792;
wire      [7:0] n7793;
wire      [7:0] n7794;
wire      [7:0] n7795;
wire      [7:0] n7796;
wire      [7:0] n7797;
wire      [7:0] n7798;
wire      [7:0] n7799;
wire      [7:0] n78;
wire      [7:0] n780;
wire      [7:0] n7800;
wire      [7:0] n7801;
wire      [7:0] n7802;
wire      [7:0] n7803;
wire      [7:0] n7804;
wire      [7:0] n7805;
wire      [7:0] n7806;
wire      [7:0] n7807;
wire      [7:0] n7808;
wire      [7:0] n7809;
wire      [7:0] n781;
wire      [7:0] n7810;
wire      [7:0] n7811;
wire      [7:0] n7812;
wire      [7:0] n7813;
wire      [7:0] n7814;
wire      [7:0] n7815;
wire      [7:0] n7816;
wire      [7:0] n7817;
wire      [7:0] n7818;
wire      [7:0] n7819;
wire      [7:0] n782;
wire      [7:0] n7820;
wire      [7:0] n7821;
wire      [7:0] n7822;
wire      [7:0] n7823;
wire      [7:0] n7824;
wire      [7:0] n7825;
wire      [7:0] n7826;
wire      [7:0] n7827;
wire      [7:0] n7828;
wire      [7:0] n7829;
wire      [7:0] n783;
wire      [7:0] n7830;
wire      [7:0] n7831;
wire      [7:0] n7832;
wire      [7:0] n7833;
wire      [7:0] n7834;
wire      [7:0] n7835;
wire      [7:0] n7836;
wire      [7:0] n7837;
wire      [7:0] n7838;
wire      [7:0] n7839;
wire      [7:0] n784;
wire      [7:0] n7840;
wire      [7:0] n7841;
wire      [7:0] n7842;
wire      [7:0] n7843;
wire      [7:0] n7844;
wire      [7:0] n7845;
wire      [7:0] n7846;
wire      [7:0] n7847;
wire      [7:0] n7848;
wire      [7:0] n7849;
wire      [7:0] n785;
wire      [7:0] n7850;
wire      [7:0] n7851;
wire      [7:0] n7852;
wire      [7:0] n7853;
wire      [7:0] n7854;
wire      [7:0] n7855;
wire      [7:0] n7856;
wire      [7:0] n7857;
wire      [7:0] n7858;
wire      [7:0] n7859;
wire      [7:0] n786;
wire      [7:0] n7860;
wire      [7:0] n7861;
wire      [7:0] n7862;
wire      [7:0] n7863;
wire      [7:0] n7864;
wire      [7:0] n7865;
wire      [7:0] n7866;
wire      [7:0] n7867;
wire      [7:0] n7868;
wire      [7:0] n7869;
wire      [7:0] n787;
wire      [7:0] n7870;
wire      [7:0] n7871;
wire      [7:0] n7872;
wire      [7:0] n7873;
wire      [7:0] n7874;
wire      [7:0] n7875;
wire      [7:0] n7876;
wire      [7:0] n7877;
wire      [7:0] n7878;
wire      [7:0] n7879;
wire      [7:0] n788;
wire      [7:0] n7880;
wire      [7:0] n7881;
wire      [7:0] n7882;
wire      [7:0] n7883;
wire      [7:0] n7884;
wire      [7:0] n7885;
wire      [7:0] n7886;
wire      [7:0] n7887;
wire      [7:0] n7888;
wire      [7:0] n7889;
wire      [7:0] n789;
wire      [7:0] n7890;
wire      [7:0] n7891;
wire      [7:0] n7892;
wire      [7:0] n7893;
wire      [7:0] n7894;
wire      [7:0] n7895;
wire      [7:0] n7896;
wire      [7:0] n7897;
wire      [7:0] n7898;
wire      [7:0] n7899;
wire      [7:0] n790;
wire      [7:0] n7900;
wire      [7:0] n7901;
wire      [7:0] n7902;
wire      [7:0] n7903;
wire      [7:0] n7904;
wire      [7:0] n7905;
wire      [7:0] n7906;
wire      [7:0] n7907;
wire      [7:0] n7908;
wire      [7:0] n7909;
wire      [7:0] n791;
wire      [7:0] n7910;
wire      [7:0] n7911;
wire      [7:0] n7912;
wire      [7:0] n7913;
wire      [7:0] n7914;
wire      [7:0] n7915;
wire      [7:0] n7916;
wire      [7:0] n7917;
wire      [7:0] n7918;
wire      [7:0] n7919;
wire      [7:0] n792;
wire      [7:0] n7920;
wire      [7:0] n7921;
wire      [7:0] n7922;
wire      [7:0] n7923;
wire      [7:0] n7924;
wire      [7:0] n7925;
wire      [7:0] n7926;
wire      [7:0] n7927;
wire      [7:0] n7928;
wire      [7:0] n7929;
wire      [7:0] n793;
wire      [7:0] n7930;
wire      [7:0] n7931;
wire      [7:0] n7932;
wire      [7:0] n7933;
wire      [7:0] n7934;
wire      [7:0] n7935;
wire      [7:0] n7936;
wire      [7:0] n7937;
wire      [7:0] n7938;
wire      [7:0] n7939;
wire      [7:0] n794;
wire      [7:0] n7940;
wire      [7:0] n7941;
wire      [7:0] n7942;
wire      [7:0] n7943;
wire      [7:0] n7944;
wire      [7:0] n7945;
wire      [7:0] n7946;
wire      [7:0] n7947;
wire      [7:0] n7948;
wire      [7:0] n7949;
wire      [7:0] n795;
wire      [7:0] n7950;
wire      [7:0] n7951;
wire      [7:0] n7952;
wire      [7:0] n7953;
wire      [7:0] n7954;
wire      [7:0] n7955;
wire      [7:0] n7956;
wire      [7:0] n7957;
wire      [7:0] n7958;
wire      [7:0] n7959;
wire      [7:0] n796;
wire      [7:0] n7960;
wire      [7:0] n7961;
wire      [7:0] n7962;
wire      [7:0] n7963;
wire      [7:0] n7964;
wire      [7:0] n7965;
wire      [7:0] n7966;
wire            n7967;
wire      [7:0] n7968;
wire            n7969;
wire      [7:0] n797;
wire      [7:0] n7970;
wire            n7971;
wire      [7:0] n7972;
wire            n7973;
wire      [7:0] n7974;
wire            n7975;
wire      [7:0] n7976;
wire            n7977;
wire      [7:0] n7978;
wire            n7979;
wire      [7:0] n798;
wire      [7:0] n7980;
wire            n7981;
wire      [7:0] n7982;
wire            n7983;
wire      [7:0] n7984;
wire            n7985;
wire      [7:0] n7986;
wire            n7987;
wire      [7:0] n7988;
wire            n7989;
wire      [7:0] n799;
wire      [7:0] n7990;
wire            n7991;
wire      [7:0] n7992;
wire            n7993;
wire      [7:0] n7994;
wire            n7995;
wire      [7:0] n7996;
wire            n7997;
wire      [7:0] n7998;
wire            n7999;
wire            n8;
wire            n80;
wire      [7:0] n800;
wire      [7:0] n8000;
wire            n8001;
wire      [7:0] n8002;
wire            n8003;
wire      [7:0] n8004;
wire            n8005;
wire      [7:0] n8006;
wire            n8007;
wire      [7:0] n8008;
wire            n8009;
wire      [7:0] n801;
wire      [7:0] n8010;
wire            n8011;
wire      [7:0] n8012;
wire            n8013;
wire      [7:0] n8014;
wire            n8015;
wire      [7:0] n8016;
wire            n8017;
wire      [7:0] n8018;
wire            n8019;
wire      [7:0] n802;
wire      [7:0] n8020;
wire            n8021;
wire      [7:0] n8022;
wire            n8023;
wire      [7:0] n8024;
wire            n8025;
wire      [7:0] n8026;
wire            n8027;
wire      [7:0] n8028;
wire            n8029;
wire      [7:0] n803;
wire      [7:0] n8030;
wire            n8031;
wire      [7:0] n8032;
wire            n8033;
wire      [7:0] n8034;
wire            n8035;
wire      [7:0] n8036;
wire            n8037;
wire      [7:0] n8038;
wire            n8039;
wire      [7:0] n804;
wire      [7:0] n8040;
wire            n8041;
wire      [7:0] n8042;
wire            n8043;
wire      [7:0] n8044;
wire            n8045;
wire      [7:0] n8046;
wire            n8047;
wire      [7:0] n8048;
wire            n8049;
wire      [7:0] n805;
wire      [7:0] n8050;
wire            n8051;
wire      [7:0] n8052;
wire            n8053;
wire      [7:0] n8054;
wire            n8055;
wire      [7:0] n8056;
wire            n8057;
wire      [7:0] n8058;
wire            n8059;
wire      [7:0] n806;
wire      [7:0] n8060;
wire            n8061;
wire      [7:0] n8062;
wire            n8063;
wire      [7:0] n8064;
wire            n8065;
wire      [7:0] n8066;
wire            n8067;
wire      [7:0] n8068;
wire            n8069;
wire      [7:0] n807;
wire      [7:0] n8070;
wire            n8071;
wire      [7:0] n8072;
wire            n8073;
wire      [7:0] n8074;
wire            n8075;
wire      [7:0] n8076;
wire            n8077;
wire      [7:0] n8078;
wire            n8079;
wire      [7:0] n808;
wire      [7:0] n8080;
wire            n8081;
wire      [7:0] n8082;
wire            n8083;
wire      [7:0] n8084;
wire            n8085;
wire      [7:0] n8086;
wire            n8087;
wire      [7:0] n8088;
wire            n8089;
wire      [7:0] n809;
wire      [7:0] n8090;
wire            n8091;
wire      [7:0] n8092;
wire            n8093;
wire      [7:0] n8094;
wire            n8095;
wire      [7:0] n8096;
wire            n8097;
wire      [7:0] n8098;
wire            n8099;
wire      [7:0] n810;
wire      [7:0] n8100;
wire            n8101;
wire      [7:0] n8102;
wire            n8103;
wire      [7:0] n8104;
wire            n8105;
wire      [7:0] n8106;
wire            n8107;
wire      [7:0] n8108;
wire            n8109;
wire      [7:0] n811;
wire      [7:0] n8110;
wire            n8111;
wire      [7:0] n8112;
wire            n8113;
wire      [7:0] n8114;
wire            n8115;
wire      [7:0] n8116;
wire            n8117;
wire      [7:0] n8118;
wire            n8119;
wire      [7:0] n812;
wire      [7:0] n8120;
wire            n8121;
wire      [7:0] n8122;
wire            n8123;
wire      [7:0] n8124;
wire            n8125;
wire      [7:0] n8126;
wire            n8127;
wire      [7:0] n8128;
wire            n8129;
wire      [7:0] n813;
wire      [7:0] n8130;
wire            n8131;
wire      [7:0] n8132;
wire            n8133;
wire      [7:0] n8134;
wire            n8135;
wire      [7:0] n8136;
wire            n8137;
wire      [7:0] n8138;
wire            n8139;
wire      [7:0] n814;
wire      [7:0] n8140;
wire            n8141;
wire      [7:0] n8142;
wire            n8143;
wire      [7:0] n8144;
wire            n8145;
wire      [7:0] n8146;
wire            n8147;
wire      [7:0] n8148;
wire            n8149;
wire      [7:0] n815;
wire      [7:0] n8150;
wire            n8151;
wire      [7:0] n8152;
wire            n8153;
wire      [7:0] n8154;
wire            n8155;
wire      [7:0] n8156;
wire            n8157;
wire      [7:0] n8158;
wire            n8159;
wire      [7:0] n816;
wire      [7:0] n8160;
wire            n8161;
wire      [7:0] n8162;
wire            n8163;
wire      [7:0] n8164;
wire            n8165;
wire      [7:0] n8166;
wire            n8167;
wire      [7:0] n8168;
wire            n8169;
wire      [7:0] n817;
wire      [7:0] n8170;
wire            n8171;
wire      [7:0] n8172;
wire            n8173;
wire      [7:0] n8174;
wire            n8175;
wire      [7:0] n8176;
wire            n8177;
wire      [7:0] n8178;
wire            n8179;
wire      [7:0] n818;
wire      [7:0] n8180;
wire            n8181;
wire      [7:0] n8182;
wire            n8183;
wire      [7:0] n8184;
wire            n8185;
wire      [7:0] n8186;
wire            n8187;
wire      [7:0] n8188;
wire            n8189;
wire      [7:0] n819;
wire      [7:0] n8190;
wire            n8191;
wire      [7:0] n8192;
wire            n8193;
wire      [7:0] n8194;
wire            n8195;
wire      [7:0] n8196;
wire            n8197;
wire      [7:0] n8198;
wire            n8199;
wire      [7:0] n82;
wire      [7:0] n820;
wire      [7:0] n8200;
wire            n8201;
wire      [7:0] n8202;
wire            n8203;
wire      [7:0] n8204;
wire            n8205;
wire      [7:0] n8206;
wire            n8207;
wire      [7:0] n8208;
wire            n8209;
wire      [7:0] n821;
wire      [7:0] n8210;
wire            n8211;
wire      [7:0] n8212;
wire            n8213;
wire      [7:0] n8214;
wire            n8215;
wire      [7:0] n8216;
wire            n8217;
wire      [7:0] n8218;
wire            n8219;
wire      [7:0] n822;
wire      [7:0] n8220;
wire            n8221;
wire      [7:0] n8222;
wire            n8223;
wire      [7:0] n8224;
wire            n8225;
wire      [7:0] n8226;
wire            n8227;
wire      [7:0] n8228;
wire            n8229;
wire      [7:0] n823;
wire      [7:0] n8230;
wire            n8231;
wire      [7:0] n8232;
wire            n8233;
wire      [7:0] n8234;
wire            n8235;
wire      [7:0] n8236;
wire            n8237;
wire      [7:0] n8238;
wire            n8239;
wire      [7:0] n824;
wire      [7:0] n8240;
wire            n8241;
wire      [7:0] n8242;
wire            n8243;
wire      [7:0] n8244;
wire            n8245;
wire      [7:0] n8246;
wire            n8247;
wire      [7:0] n8248;
wire            n8249;
wire      [7:0] n825;
wire      [7:0] n8250;
wire            n8251;
wire      [7:0] n8252;
wire            n8253;
wire      [7:0] n8254;
wire            n8255;
wire      [7:0] n8256;
wire            n8257;
wire      [7:0] n8258;
wire            n8259;
wire      [7:0] n826;
wire      [7:0] n8260;
wire            n8261;
wire      [7:0] n8262;
wire            n8263;
wire      [7:0] n8264;
wire            n8265;
wire      [7:0] n8266;
wire            n8267;
wire      [7:0] n8268;
wire            n8269;
wire      [7:0] n827;
wire      [7:0] n8270;
wire            n8271;
wire      [7:0] n8272;
wire            n8273;
wire      [7:0] n8274;
wire            n8275;
wire      [7:0] n8276;
wire            n8277;
wire      [7:0] n8278;
wire            n8279;
wire      [7:0] n828;
wire      [7:0] n8280;
wire            n8281;
wire      [7:0] n8282;
wire            n8283;
wire      [7:0] n8284;
wire            n8285;
wire      [7:0] n8286;
wire            n8287;
wire      [7:0] n8288;
wire            n8289;
wire      [7:0] n829;
wire      [7:0] n8290;
wire            n8291;
wire      [7:0] n8292;
wire            n8293;
wire      [7:0] n8294;
wire            n8295;
wire      [7:0] n8296;
wire            n8297;
wire      [7:0] n8298;
wire            n8299;
wire      [7:0] n830;
wire      [7:0] n8300;
wire            n8301;
wire      [7:0] n8302;
wire            n8303;
wire      [7:0] n8304;
wire            n8305;
wire      [7:0] n8306;
wire            n8307;
wire      [7:0] n8308;
wire            n8309;
wire      [7:0] n831;
wire      [7:0] n8310;
wire            n8311;
wire      [7:0] n8312;
wire            n8313;
wire      [7:0] n8314;
wire            n8315;
wire      [7:0] n8316;
wire            n8317;
wire      [7:0] n8318;
wire            n8319;
wire      [7:0] n832;
wire      [7:0] n8320;
wire            n8321;
wire      [7:0] n8322;
wire            n8323;
wire      [7:0] n8324;
wire            n8325;
wire      [7:0] n8326;
wire            n8327;
wire      [7:0] n8328;
wire            n8329;
wire      [7:0] n833;
wire      [7:0] n8330;
wire            n8331;
wire      [7:0] n8332;
wire            n8333;
wire      [7:0] n8334;
wire            n8335;
wire      [7:0] n8336;
wire            n8337;
wire      [7:0] n8338;
wire            n8339;
wire      [7:0] n834;
wire      [7:0] n8340;
wire            n8341;
wire      [7:0] n8342;
wire            n8343;
wire      [7:0] n8344;
wire            n8345;
wire      [7:0] n8346;
wire            n8347;
wire      [7:0] n8348;
wire            n8349;
wire      [7:0] n835;
wire      [7:0] n8350;
wire            n8351;
wire      [7:0] n8352;
wire            n8353;
wire      [7:0] n8354;
wire            n8355;
wire      [7:0] n8356;
wire            n8357;
wire      [7:0] n8358;
wire            n8359;
wire      [7:0] n836;
wire      [7:0] n8360;
wire            n8361;
wire      [7:0] n8362;
wire            n8363;
wire      [7:0] n8364;
wire            n8365;
wire      [7:0] n8366;
wire            n8367;
wire      [7:0] n8368;
wire            n8369;
wire      [7:0] n837;
wire      [7:0] n8370;
wire            n8371;
wire      [7:0] n8372;
wire            n8373;
wire      [7:0] n8374;
wire            n8375;
wire      [7:0] n8376;
wire            n8377;
wire      [7:0] n8378;
wire            n8379;
wire      [7:0] n838;
wire      [7:0] n8380;
wire            n8381;
wire      [7:0] n8382;
wire            n8383;
wire      [7:0] n8384;
wire            n8385;
wire      [7:0] n8386;
wire            n8387;
wire      [7:0] n8388;
wire            n8389;
wire      [7:0] n839;
wire      [7:0] n8390;
wire            n8391;
wire      [7:0] n8392;
wire            n8393;
wire      [7:0] n8394;
wire            n8395;
wire      [7:0] n8396;
wire            n8397;
wire      [7:0] n8398;
wire            n8399;
wire            n84;
wire      [7:0] n840;
wire      [7:0] n8400;
wire            n8401;
wire      [7:0] n8402;
wire            n8403;
wire      [7:0] n8404;
wire            n8405;
wire      [7:0] n8406;
wire            n8407;
wire      [7:0] n8408;
wire            n8409;
wire      [7:0] n841;
wire      [7:0] n8410;
wire            n8411;
wire      [7:0] n8412;
wire            n8413;
wire      [7:0] n8414;
wire            n8415;
wire      [7:0] n8416;
wire            n8417;
wire      [7:0] n8418;
wire            n8419;
wire      [7:0] n842;
wire      [7:0] n8420;
wire            n8421;
wire      [7:0] n8422;
wire            n8423;
wire      [7:0] n8424;
wire            n8425;
wire      [7:0] n8426;
wire            n8427;
wire      [7:0] n8428;
wire            n8429;
wire      [7:0] n843;
wire      [7:0] n8430;
wire            n8431;
wire      [7:0] n8432;
wire            n8433;
wire      [7:0] n8434;
wire            n8435;
wire      [7:0] n8436;
wire            n8437;
wire      [7:0] n8438;
wire            n8439;
wire      [7:0] n844;
wire      [7:0] n8440;
wire            n8441;
wire      [7:0] n8442;
wire            n8443;
wire      [7:0] n8444;
wire            n8445;
wire      [7:0] n8446;
wire            n8447;
wire      [7:0] n8448;
wire            n8449;
wire      [7:0] n845;
wire      [7:0] n8450;
wire            n8451;
wire      [7:0] n8452;
wire            n8453;
wire      [7:0] n8454;
wire            n8455;
wire      [7:0] n8456;
wire            n8457;
wire      [7:0] n8458;
wire            n8459;
wire      [7:0] n846;
wire      [7:0] n8460;
wire            n8461;
wire      [7:0] n8462;
wire            n8463;
wire      [7:0] n8464;
wire            n8465;
wire      [7:0] n8466;
wire            n8467;
wire      [7:0] n8468;
wire            n8469;
wire      [7:0] n847;
wire      [7:0] n8470;
wire            n8471;
wire      [7:0] n8472;
wire            n8473;
wire      [7:0] n8474;
wire            n8475;
wire      [7:0] n8476;
wire            n8477;
wire      [7:0] n8478;
wire      [7:0] n8479;
wire      [7:0] n848;
wire      [7:0] n8480;
wire      [7:0] n8481;
wire      [7:0] n8482;
wire      [7:0] n8483;
wire      [7:0] n8484;
wire      [7:0] n8485;
wire      [7:0] n8486;
wire      [7:0] n8487;
wire      [7:0] n8488;
wire      [7:0] n8489;
wire      [7:0] n849;
wire      [7:0] n8490;
wire      [7:0] n8491;
wire      [7:0] n8492;
wire      [7:0] n8493;
wire      [7:0] n8494;
wire      [7:0] n8495;
wire      [7:0] n8496;
wire      [7:0] n8497;
wire      [7:0] n8498;
wire      [7:0] n8499;
wire      [7:0] n850;
wire      [7:0] n8500;
wire      [7:0] n8501;
wire      [7:0] n8502;
wire      [7:0] n8503;
wire      [7:0] n8504;
wire      [7:0] n8505;
wire      [7:0] n8506;
wire      [7:0] n8507;
wire      [7:0] n8508;
wire      [7:0] n8509;
wire      [7:0] n851;
wire      [7:0] n8510;
wire      [7:0] n8511;
wire      [7:0] n8512;
wire      [7:0] n8513;
wire      [7:0] n8514;
wire      [7:0] n8515;
wire      [7:0] n8516;
wire      [7:0] n8517;
wire      [7:0] n8518;
wire      [7:0] n8519;
wire      [7:0] n852;
wire      [7:0] n8520;
wire      [7:0] n8521;
wire      [7:0] n8522;
wire      [7:0] n8523;
wire      [7:0] n8524;
wire      [7:0] n8525;
wire      [7:0] n8526;
wire      [7:0] n8527;
wire      [7:0] n8528;
wire      [7:0] n8529;
wire      [7:0] n853;
wire      [7:0] n8530;
wire      [7:0] n8531;
wire      [7:0] n8532;
wire      [7:0] n8533;
wire      [7:0] n8534;
wire      [7:0] n8535;
wire      [7:0] n8536;
wire      [7:0] n8537;
wire      [7:0] n8538;
wire      [7:0] n8539;
wire      [7:0] n854;
wire      [7:0] n8540;
wire      [7:0] n8541;
wire      [7:0] n8542;
wire      [7:0] n8543;
wire      [7:0] n8544;
wire      [7:0] n8545;
wire      [7:0] n8546;
wire      [7:0] n8547;
wire      [7:0] n8548;
wire      [7:0] n8549;
wire      [7:0] n855;
wire      [7:0] n8550;
wire      [7:0] n8551;
wire      [7:0] n8552;
wire      [7:0] n8553;
wire      [7:0] n8554;
wire      [7:0] n8555;
wire      [7:0] n8556;
wire      [7:0] n8557;
wire      [7:0] n8558;
wire      [7:0] n8559;
wire      [7:0] n856;
wire      [7:0] n8560;
wire      [7:0] n8561;
wire      [7:0] n8562;
wire      [7:0] n8563;
wire      [7:0] n8564;
wire      [7:0] n8565;
wire      [7:0] n8566;
wire      [7:0] n8567;
wire      [7:0] n8568;
wire      [7:0] n8569;
wire      [7:0] n857;
wire      [7:0] n8570;
wire      [7:0] n8571;
wire      [7:0] n8572;
wire      [7:0] n8573;
wire      [7:0] n8574;
wire      [7:0] n8575;
wire      [7:0] n8576;
wire      [7:0] n8577;
wire      [7:0] n8578;
wire      [7:0] n8579;
wire      [7:0] n858;
wire      [7:0] n8580;
wire      [7:0] n8581;
wire      [7:0] n8582;
wire      [7:0] n8583;
wire      [7:0] n8584;
wire      [7:0] n8585;
wire      [7:0] n8586;
wire      [7:0] n8587;
wire      [7:0] n8588;
wire      [7:0] n8589;
wire      [7:0] n859;
wire      [7:0] n8590;
wire      [7:0] n8591;
wire      [7:0] n8592;
wire      [7:0] n8593;
wire      [7:0] n8594;
wire      [7:0] n8595;
wire      [7:0] n8596;
wire      [7:0] n8597;
wire      [7:0] n8598;
wire      [7:0] n8599;
wire      [7:0] n86;
wire      [7:0] n860;
wire      [7:0] n8600;
wire      [7:0] n8601;
wire      [7:0] n8602;
wire      [7:0] n8603;
wire      [7:0] n8604;
wire      [7:0] n8605;
wire      [7:0] n8606;
wire      [7:0] n8607;
wire      [7:0] n8608;
wire      [7:0] n8609;
wire      [7:0] n861;
wire      [7:0] n8610;
wire      [7:0] n8611;
wire      [7:0] n8612;
wire      [7:0] n8613;
wire      [7:0] n8614;
wire      [7:0] n8615;
wire      [7:0] n8616;
wire      [7:0] n8617;
wire      [7:0] n8618;
wire      [7:0] n8619;
wire      [7:0] n862;
wire      [7:0] n8620;
wire      [7:0] n8621;
wire      [7:0] n8622;
wire      [7:0] n8623;
wire      [7:0] n8624;
wire      [7:0] n8625;
wire      [7:0] n8626;
wire      [7:0] n8627;
wire      [7:0] n8628;
wire      [7:0] n8629;
wire      [7:0] n863;
wire      [7:0] n8630;
wire      [7:0] n8631;
wire      [7:0] n8632;
wire      [7:0] n8633;
wire      [7:0] n8634;
wire      [7:0] n8635;
wire      [7:0] n8636;
wire      [7:0] n8637;
wire      [7:0] n8638;
wire      [7:0] n8639;
wire      [7:0] n864;
wire      [7:0] n8640;
wire      [7:0] n8641;
wire      [7:0] n8642;
wire      [7:0] n8643;
wire      [7:0] n8644;
wire      [7:0] n8645;
wire      [7:0] n8646;
wire      [7:0] n8647;
wire      [7:0] n8648;
wire      [7:0] n8649;
wire      [7:0] n865;
wire      [7:0] n8650;
wire      [7:0] n8651;
wire      [7:0] n8652;
wire      [7:0] n8653;
wire      [7:0] n8654;
wire      [7:0] n8655;
wire      [7:0] n8656;
wire      [7:0] n8657;
wire      [7:0] n8658;
wire      [7:0] n8659;
wire      [7:0] n866;
wire      [7:0] n8660;
wire      [7:0] n8661;
wire      [7:0] n8662;
wire      [7:0] n8663;
wire      [7:0] n8664;
wire      [7:0] n8665;
wire      [7:0] n8666;
wire      [7:0] n8667;
wire      [7:0] n8668;
wire      [7:0] n8669;
wire      [7:0] n867;
wire      [7:0] n8670;
wire      [7:0] n8671;
wire      [7:0] n8672;
wire      [7:0] n8673;
wire      [7:0] n8674;
wire      [7:0] n8675;
wire      [7:0] n8676;
wire      [7:0] n8677;
wire      [7:0] n8678;
wire      [7:0] n8679;
wire      [7:0] n868;
wire      [7:0] n8680;
wire      [7:0] n8681;
wire      [7:0] n8682;
wire      [7:0] n8683;
wire      [7:0] n8684;
wire      [7:0] n8685;
wire      [7:0] n8686;
wire      [7:0] n8687;
wire      [7:0] n8688;
wire      [7:0] n8689;
wire      [7:0] n869;
wire      [7:0] n8690;
wire      [7:0] n8691;
wire      [7:0] n8692;
wire      [7:0] n8693;
wire      [7:0] n8694;
wire      [7:0] n8695;
wire      [7:0] n8696;
wire      [7:0] n8697;
wire      [7:0] n8698;
wire      [7:0] n8699;
wire      [7:0] n870;
wire      [7:0] n8700;
wire      [7:0] n8701;
wire      [7:0] n8702;
wire      [7:0] n8703;
wire      [7:0] n8704;
wire      [7:0] n8705;
wire      [7:0] n8706;
wire      [7:0] n8707;
wire      [7:0] n8708;
wire      [7:0] n8709;
wire      [7:0] n871;
wire      [7:0] n8710;
wire      [7:0] n8711;
wire      [7:0] n8712;
wire      [7:0] n8713;
wire      [7:0] n8714;
wire      [7:0] n8715;
wire      [7:0] n8716;
wire      [7:0] n8717;
wire      [7:0] n8718;
wire      [7:0] n8719;
wire      [7:0] n872;
wire      [7:0] n8720;
wire      [7:0] n8721;
wire      [7:0] n8722;
wire      [7:0] n8723;
wire      [7:0] n8724;
wire      [7:0] n8725;
wire      [7:0] n8726;
wire      [7:0] n8727;
wire      [7:0] n8728;
wire      [7:0] n8729;
wire      [7:0] n873;
wire      [7:0] n8730;
wire      [7:0] n8731;
wire      [7:0] n8732;
wire      [7:0] n8733;
wire      [7:0] n8734;
wire      [7:0] n8735;
wire            n8736;
wire      [7:0] n8737;
wire            n8738;
wire      [7:0] n8739;
wire      [7:0] n874;
wire            n8740;
wire      [7:0] n8741;
wire            n8742;
wire      [7:0] n8743;
wire            n8744;
wire      [7:0] n8745;
wire            n8746;
wire      [7:0] n8747;
wire            n8748;
wire      [7:0] n8749;
wire      [7:0] n875;
wire            n8750;
wire      [7:0] n8751;
wire            n8752;
wire      [7:0] n8753;
wire            n8754;
wire      [7:0] n8755;
wire            n8756;
wire      [7:0] n8757;
wire            n8758;
wire      [7:0] n8759;
wire      [7:0] n876;
wire            n8760;
wire      [7:0] n8761;
wire            n8762;
wire      [7:0] n8763;
wire            n8764;
wire      [7:0] n8765;
wire            n8766;
wire      [7:0] n8767;
wire            n8768;
wire      [7:0] n8769;
wire      [7:0] n877;
wire            n8770;
wire      [7:0] n8771;
wire            n8772;
wire      [7:0] n8773;
wire            n8774;
wire      [7:0] n8775;
wire            n8776;
wire      [7:0] n8777;
wire            n8778;
wire      [7:0] n8779;
wire      [7:0] n878;
wire            n8780;
wire      [7:0] n8781;
wire            n8782;
wire      [7:0] n8783;
wire            n8784;
wire      [7:0] n8785;
wire            n8786;
wire      [7:0] n8787;
wire            n8788;
wire      [7:0] n8789;
wire      [7:0] n879;
wire            n8790;
wire      [7:0] n8791;
wire            n8792;
wire      [7:0] n8793;
wire            n8794;
wire      [7:0] n8795;
wire            n8796;
wire      [7:0] n8797;
wire            n8798;
wire      [7:0] n8799;
wire            n88;
wire      [7:0] n880;
wire            n8800;
wire      [7:0] n8801;
wire            n8802;
wire      [7:0] n8803;
wire            n8804;
wire      [7:0] n8805;
wire            n8806;
wire      [7:0] n8807;
wire            n8808;
wire      [7:0] n8809;
wire      [7:0] n881;
wire            n8810;
wire      [7:0] n8811;
wire            n8812;
wire      [7:0] n8813;
wire            n8814;
wire      [7:0] n8815;
wire            n8816;
wire      [7:0] n8817;
wire            n8818;
wire      [7:0] n8819;
wire      [7:0] n882;
wire            n8820;
wire      [7:0] n8821;
wire            n8822;
wire      [7:0] n8823;
wire            n8824;
wire      [7:0] n8825;
wire            n8826;
wire      [7:0] n8827;
wire            n8828;
wire      [7:0] n8829;
wire      [7:0] n883;
wire            n8830;
wire      [7:0] n8831;
wire            n8832;
wire      [7:0] n8833;
wire            n8834;
wire      [7:0] n8835;
wire            n8836;
wire      [7:0] n8837;
wire            n8838;
wire      [7:0] n8839;
wire      [7:0] n884;
wire            n8840;
wire      [7:0] n8841;
wire            n8842;
wire      [7:0] n8843;
wire            n8844;
wire      [7:0] n8845;
wire            n8846;
wire      [7:0] n8847;
wire            n8848;
wire      [7:0] n8849;
wire      [7:0] n885;
wire            n8850;
wire      [7:0] n8851;
wire            n8852;
wire      [7:0] n8853;
wire            n8854;
wire      [7:0] n8855;
wire            n8856;
wire      [7:0] n8857;
wire            n8858;
wire      [7:0] n8859;
wire      [7:0] n886;
wire            n8860;
wire      [7:0] n8861;
wire            n8862;
wire      [7:0] n8863;
wire            n8864;
wire      [7:0] n8865;
wire            n8866;
wire      [7:0] n8867;
wire            n8868;
wire      [7:0] n8869;
wire      [7:0] n887;
wire            n8870;
wire      [7:0] n8871;
wire            n8872;
wire      [7:0] n8873;
wire            n8874;
wire      [7:0] n8875;
wire            n8876;
wire      [7:0] n8877;
wire            n8878;
wire      [7:0] n8879;
wire      [7:0] n888;
wire            n8880;
wire      [7:0] n8881;
wire            n8882;
wire      [7:0] n8883;
wire            n8884;
wire      [7:0] n8885;
wire            n8886;
wire      [7:0] n8887;
wire            n8888;
wire      [7:0] n8889;
wire      [7:0] n889;
wire            n8890;
wire      [7:0] n8891;
wire            n8892;
wire      [7:0] n8893;
wire            n8894;
wire      [7:0] n8895;
wire            n8896;
wire      [7:0] n8897;
wire            n8898;
wire      [7:0] n8899;
wire      [7:0] n890;
wire            n8900;
wire      [7:0] n8901;
wire            n8902;
wire      [7:0] n8903;
wire            n8904;
wire      [7:0] n8905;
wire            n8906;
wire      [7:0] n8907;
wire            n8908;
wire      [7:0] n8909;
wire      [7:0] n891;
wire            n8910;
wire      [7:0] n8911;
wire            n8912;
wire      [7:0] n8913;
wire            n8914;
wire      [7:0] n8915;
wire            n8916;
wire      [7:0] n8917;
wire            n8918;
wire      [7:0] n8919;
wire      [7:0] n892;
wire            n8920;
wire      [7:0] n8921;
wire            n8922;
wire      [7:0] n8923;
wire            n8924;
wire      [7:0] n8925;
wire            n8926;
wire      [7:0] n8927;
wire            n8928;
wire      [7:0] n8929;
wire      [7:0] n893;
wire            n8930;
wire      [7:0] n8931;
wire            n8932;
wire      [7:0] n8933;
wire            n8934;
wire      [7:0] n8935;
wire            n8936;
wire      [7:0] n8937;
wire            n8938;
wire      [7:0] n8939;
wire      [7:0] n894;
wire            n8940;
wire      [7:0] n8941;
wire            n8942;
wire      [7:0] n8943;
wire            n8944;
wire      [7:0] n8945;
wire            n8946;
wire      [7:0] n8947;
wire            n8948;
wire      [7:0] n8949;
wire      [7:0] n895;
wire            n8950;
wire      [7:0] n8951;
wire            n8952;
wire      [7:0] n8953;
wire            n8954;
wire      [7:0] n8955;
wire            n8956;
wire      [7:0] n8957;
wire            n8958;
wire      [7:0] n8959;
wire      [7:0] n896;
wire            n8960;
wire      [7:0] n8961;
wire            n8962;
wire      [7:0] n8963;
wire            n8964;
wire      [7:0] n8965;
wire            n8966;
wire      [7:0] n8967;
wire            n8968;
wire      [7:0] n8969;
wire      [7:0] n897;
wire            n8970;
wire      [7:0] n8971;
wire            n8972;
wire      [7:0] n8973;
wire            n8974;
wire      [7:0] n8975;
wire            n8976;
wire      [7:0] n8977;
wire            n8978;
wire      [7:0] n8979;
wire      [7:0] n898;
wire            n8980;
wire      [7:0] n8981;
wire            n8982;
wire      [7:0] n8983;
wire            n8984;
wire      [7:0] n8985;
wire            n8986;
wire      [7:0] n8987;
wire            n8988;
wire      [7:0] n8989;
wire      [7:0] n899;
wire            n8990;
wire      [7:0] n8991;
wire            n8992;
wire      [7:0] n8993;
wire            n8994;
wire      [7:0] n8995;
wire            n8996;
wire      [7:0] n8997;
wire            n8998;
wire      [7:0] n8999;
wire      [7:0] n90;
wire      [7:0] n900;
wire            n9000;
wire      [7:0] n9001;
wire            n9002;
wire      [7:0] n9003;
wire            n9004;
wire      [7:0] n9005;
wire            n9006;
wire      [7:0] n9007;
wire            n9008;
wire      [7:0] n9009;
wire      [7:0] n901;
wire            n9010;
wire      [7:0] n9011;
wire            n9012;
wire      [7:0] n9013;
wire            n9014;
wire      [7:0] n9015;
wire            n9016;
wire      [7:0] n9017;
wire            n9018;
wire      [7:0] n9019;
wire      [7:0] n902;
wire            n9020;
wire      [7:0] n9021;
wire            n9022;
wire      [7:0] n9023;
wire            n9024;
wire      [7:0] n9025;
wire            n9026;
wire      [7:0] n9027;
wire            n9028;
wire      [7:0] n9029;
wire      [7:0] n903;
wire            n9030;
wire      [7:0] n9031;
wire            n9032;
wire      [7:0] n9033;
wire            n9034;
wire      [7:0] n9035;
wire            n9036;
wire      [7:0] n9037;
wire            n9038;
wire      [7:0] n9039;
wire      [7:0] n904;
wire            n9040;
wire      [7:0] n9041;
wire            n9042;
wire      [7:0] n9043;
wire            n9044;
wire      [7:0] n9045;
wire            n9046;
wire      [7:0] n9047;
wire            n9048;
wire      [7:0] n9049;
wire      [7:0] n905;
wire            n9050;
wire      [7:0] n9051;
wire            n9052;
wire      [7:0] n9053;
wire            n9054;
wire      [7:0] n9055;
wire            n9056;
wire      [7:0] n9057;
wire            n9058;
wire      [7:0] n9059;
wire      [7:0] n906;
wire            n9060;
wire      [7:0] n9061;
wire            n9062;
wire      [7:0] n9063;
wire            n9064;
wire      [7:0] n9065;
wire            n9066;
wire      [7:0] n9067;
wire            n9068;
wire      [7:0] n9069;
wire      [7:0] n907;
wire            n9070;
wire      [7:0] n9071;
wire            n9072;
wire      [7:0] n9073;
wire            n9074;
wire      [7:0] n9075;
wire            n9076;
wire      [7:0] n9077;
wire            n9078;
wire      [7:0] n9079;
wire      [7:0] n908;
wire            n9080;
wire      [7:0] n9081;
wire            n9082;
wire      [7:0] n9083;
wire            n9084;
wire      [7:0] n9085;
wire            n9086;
wire      [7:0] n9087;
wire            n9088;
wire      [7:0] n9089;
wire      [7:0] n909;
wire            n9090;
wire      [7:0] n9091;
wire            n9092;
wire      [7:0] n9093;
wire            n9094;
wire      [7:0] n9095;
wire            n9096;
wire      [7:0] n9097;
wire            n9098;
wire      [7:0] n9099;
wire      [7:0] n910;
wire            n9100;
wire      [7:0] n9101;
wire            n9102;
wire      [7:0] n9103;
wire            n9104;
wire      [7:0] n9105;
wire            n9106;
wire      [7:0] n9107;
wire            n9108;
wire      [7:0] n9109;
wire      [7:0] n911;
wire            n9110;
wire      [7:0] n9111;
wire            n9112;
wire      [7:0] n9113;
wire            n9114;
wire      [7:0] n9115;
wire            n9116;
wire      [7:0] n9117;
wire            n9118;
wire      [7:0] n9119;
wire      [7:0] n912;
wire            n9120;
wire      [7:0] n9121;
wire            n9122;
wire      [7:0] n9123;
wire            n9124;
wire      [7:0] n9125;
wire            n9126;
wire      [7:0] n9127;
wire            n9128;
wire      [7:0] n9129;
wire      [7:0] n913;
wire            n9130;
wire      [7:0] n9131;
wire            n9132;
wire      [7:0] n9133;
wire            n9134;
wire      [7:0] n9135;
wire            n9136;
wire      [7:0] n9137;
wire            n9138;
wire      [7:0] n9139;
wire      [7:0] n914;
wire            n9140;
wire      [7:0] n9141;
wire            n9142;
wire      [7:0] n9143;
wire            n9144;
wire      [7:0] n9145;
wire            n9146;
wire      [7:0] n9147;
wire            n9148;
wire      [7:0] n9149;
wire      [7:0] n915;
wire            n9150;
wire      [7:0] n9151;
wire            n9152;
wire      [7:0] n9153;
wire            n9154;
wire      [7:0] n9155;
wire            n9156;
wire      [7:0] n9157;
wire            n9158;
wire      [7:0] n9159;
wire      [7:0] n916;
wire            n9160;
wire      [7:0] n9161;
wire            n9162;
wire      [7:0] n9163;
wire            n9164;
wire      [7:0] n9165;
wire            n9166;
wire      [7:0] n9167;
wire            n9168;
wire      [7:0] n9169;
wire      [7:0] n917;
wire            n9170;
wire      [7:0] n9171;
wire            n9172;
wire      [7:0] n9173;
wire            n9174;
wire      [7:0] n9175;
wire            n9176;
wire      [7:0] n9177;
wire            n9178;
wire      [7:0] n9179;
wire      [7:0] n918;
wire            n9180;
wire      [7:0] n9181;
wire            n9182;
wire      [7:0] n9183;
wire            n9184;
wire      [7:0] n9185;
wire            n9186;
wire      [7:0] n9187;
wire            n9188;
wire      [7:0] n9189;
wire      [7:0] n919;
wire            n9190;
wire      [7:0] n9191;
wire            n9192;
wire      [7:0] n9193;
wire            n9194;
wire      [7:0] n9195;
wire            n9196;
wire      [7:0] n9197;
wire            n9198;
wire      [7:0] n9199;
wire            n92;
wire      [7:0] n920;
wire            n9200;
wire      [7:0] n9201;
wire            n9202;
wire      [7:0] n9203;
wire            n9204;
wire      [7:0] n9205;
wire            n9206;
wire      [7:0] n9207;
wire            n9208;
wire      [7:0] n9209;
wire      [7:0] n921;
wire            n9210;
wire      [7:0] n9211;
wire            n9212;
wire      [7:0] n9213;
wire            n9214;
wire      [7:0] n9215;
wire            n9216;
wire      [7:0] n9217;
wire            n9218;
wire      [7:0] n9219;
wire      [7:0] n922;
wire            n9220;
wire      [7:0] n9221;
wire            n9222;
wire      [7:0] n9223;
wire            n9224;
wire      [7:0] n9225;
wire            n9226;
wire      [7:0] n9227;
wire            n9228;
wire      [7:0] n9229;
wire      [7:0] n923;
wire            n9230;
wire      [7:0] n9231;
wire            n9232;
wire      [7:0] n9233;
wire            n9234;
wire      [7:0] n9235;
wire            n9236;
wire      [7:0] n9237;
wire            n9238;
wire      [7:0] n9239;
wire      [7:0] n924;
wire            n9240;
wire      [7:0] n9241;
wire            n9242;
wire      [7:0] n9243;
wire            n9244;
wire      [7:0] n9245;
wire            n9246;
wire      [7:0] n9247;
wire      [7:0] n9248;
wire      [7:0] n9249;
wire      [7:0] n925;
wire      [7:0] n9250;
wire      [7:0] n9251;
wire      [7:0] n9252;
wire      [7:0] n9253;
wire      [7:0] n9254;
wire      [7:0] n9255;
wire      [7:0] n9256;
wire      [7:0] n9257;
wire      [7:0] n9258;
wire      [7:0] n9259;
wire      [7:0] n926;
wire      [7:0] n9260;
wire      [7:0] n9261;
wire      [7:0] n9262;
wire      [7:0] n9263;
wire      [7:0] n9264;
wire      [7:0] n9265;
wire      [7:0] n9266;
wire      [7:0] n9267;
wire      [7:0] n9268;
wire      [7:0] n9269;
wire      [7:0] n927;
wire      [7:0] n9270;
wire      [7:0] n9271;
wire      [7:0] n9272;
wire      [7:0] n9273;
wire      [7:0] n9274;
wire      [7:0] n9275;
wire      [7:0] n9276;
wire      [7:0] n9277;
wire      [7:0] n9278;
wire      [7:0] n9279;
wire      [7:0] n928;
wire      [7:0] n9280;
wire      [7:0] n9281;
wire      [7:0] n9282;
wire      [7:0] n9283;
wire      [7:0] n9284;
wire      [7:0] n9285;
wire      [7:0] n9286;
wire      [7:0] n9287;
wire      [7:0] n9288;
wire      [7:0] n9289;
wire      [7:0] n929;
wire      [7:0] n9290;
wire      [7:0] n9291;
wire      [7:0] n9292;
wire      [7:0] n9293;
wire      [7:0] n9294;
wire      [7:0] n9295;
wire      [7:0] n9296;
wire      [7:0] n9297;
wire      [7:0] n9298;
wire      [7:0] n9299;
wire      [7:0] n930;
wire      [7:0] n9300;
wire      [7:0] n9301;
wire      [7:0] n9302;
wire      [7:0] n9303;
wire      [7:0] n9304;
wire      [7:0] n9305;
wire      [7:0] n9306;
wire      [7:0] n9307;
wire      [7:0] n9308;
wire      [7:0] n9309;
wire      [7:0] n931;
wire      [7:0] n9310;
wire      [7:0] n9311;
wire      [7:0] n9312;
wire      [7:0] n9313;
wire      [7:0] n9314;
wire      [7:0] n9315;
wire      [7:0] n9316;
wire      [7:0] n9317;
wire      [7:0] n9318;
wire      [7:0] n9319;
wire      [7:0] n932;
wire      [7:0] n9320;
wire      [7:0] n9321;
wire      [7:0] n9322;
wire      [7:0] n9323;
wire      [7:0] n9324;
wire      [7:0] n9325;
wire      [7:0] n9326;
wire      [7:0] n9327;
wire      [7:0] n9328;
wire      [7:0] n9329;
wire      [7:0] n933;
wire      [7:0] n9330;
wire      [7:0] n9331;
wire      [7:0] n9332;
wire      [7:0] n9333;
wire      [7:0] n9334;
wire      [7:0] n9335;
wire      [7:0] n9336;
wire      [7:0] n9337;
wire      [7:0] n9338;
wire      [7:0] n9339;
wire      [7:0] n934;
wire      [7:0] n9340;
wire      [7:0] n9341;
wire      [7:0] n9342;
wire      [7:0] n9343;
wire      [7:0] n9344;
wire      [7:0] n9345;
wire      [7:0] n9346;
wire      [7:0] n9347;
wire      [7:0] n9348;
wire      [7:0] n9349;
wire      [7:0] n935;
wire      [7:0] n9350;
wire      [7:0] n9351;
wire      [7:0] n9352;
wire      [7:0] n9353;
wire      [7:0] n9354;
wire      [7:0] n9355;
wire      [7:0] n9356;
wire      [7:0] n9357;
wire      [7:0] n9358;
wire      [7:0] n9359;
wire      [7:0] n936;
wire      [7:0] n9360;
wire      [7:0] n9361;
wire      [7:0] n9362;
wire      [7:0] n9363;
wire      [7:0] n9364;
wire      [7:0] n9365;
wire      [7:0] n9366;
wire      [7:0] n9367;
wire      [7:0] n9368;
wire      [7:0] n9369;
wire      [7:0] n937;
wire      [7:0] n9370;
wire      [7:0] n9371;
wire      [7:0] n9372;
wire      [7:0] n9373;
wire      [7:0] n9374;
wire      [7:0] n9375;
wire      [7:0] n9376;
wire      [7:0] n9377;
wire      [7:0] n9378;
wire      [7:0] n9379;
wire      [7:0] n938;
wire      [7:0] n9380;
wire      [7:0] n9381;
wire      [7:0] n9382;
wire      [7:0] n9383;
wire      [7:0] n9384;
wire      [7:0] n9385;
wire      [7:0] n9386;
wire      [7:0] n9387;
wire      [7:0] n9388;
wire      [7:0] n9389;
wire      [7:0] n939;
wire      [7:0] n9390;
wire      [7:0] n9391;
wire      [7:0] n9392;
wire      [7:0] n9393;
wire      [7:0] n9394;
wire      [7:0] n9395;
wire      [7:0] n9396;
wire      [7:0] n9397;
wire      [7:0] n9398;
wire      [7:0] n9399;
wire      [7:0] n94;
wire      [7:0] n940;
wire      [7:0] n9400;
wire      [7:0] n9401;
wire      [7:0] n9402;
wire      [7:0] n9403;
wire      [7:0] n9404;
wire      [7:0] n9405;
wire      [7:0] n9406;
wire      [7:0] n9407;
wire      [7:0] n9408;
wire      [7:0] n9409;
wire      [7:0] n941;
wire      [7:0] n9410;
wire      [7:0] n9411;
wire      [7:0] n9412;
wire      [7:0] n9413;
wire      [7:0] n9414;
wire      [7:0] n9415;
wire      [7:0] n9416;
wire      [7:0] n9417;
wire      [7:0] n9418;
wire      [7:0] n9419;
wire      [7:0] n942;
wire      [7:0] n9420;
wire      [7:0] n9421;
wire      [7:0] n9422;
wire      [7:0] n9423;
wire      [7:0] n9424;
wire      [7:0] n9425;
wire      [7:0] n9426;
wire      [7:0] n9427;
wire      [7:0] n9428;
wire      [7:0] n9429;
wire      [7:0] n943;
wire      [7:0] n9430;
wire      [7:0] n9431;
wire      [7:0] n9432;
wire      [7:0] n9433;
wire      [7:0] n9434;
wire      [7:0] n9435;
wire      [7:0] n9436;
wire      [7:0] n9437;
wire      [7:0] n9438;
wire      [7:0] n9439;
wire      [7:0] n944;
wire      [7:0] n9440;
wire      [7:0] n9441;
wire      [7:0] n9442;
wire      [7:0] n9443;
wire      [7:0] n9444;
wire      [7:0] n9445;
wire      [7:0] n9446;
wire      [7:0] n9447;
wire      [7:0] n9448;
wire      [7:0] n9449;
wire      [7:0] n945;
wire      [7:0] n9450;
wire      [7:0] n9451;
wire      [7:0] n9452;
wire      [7:0] n9453;
wire      [7:0] n9454;
wire      [7:0] n9455;
wire      [7:0] n9456;
wire      [7:0] n9457;
wire      [7:0] n9458;
wire      [7:0] n9459;
wire      [7:0] n946;
wire      [7:0] n9460;
wire      [7:0] n9461;
wire      [7:0] n9462;
wire      [7:0] n9463;
wire      [7:0] n9464;
wire      [7:0] n9465;
wire      [7:0] n9466;
wire      [7:0] n9467;
wire      [7:0] n9468;
wire      [7:0] n9469;
wire      [7:0] n947;
wire      [7:0] n9470;
wire      [7:0] n9471;
wire      [7:0] n9472;
wire      [7:0] n9473;
wire      [7:0] n9474;
wire      [7:0] n9475;
wire      [7:0] n9476;
wire      [7:0] n9477;
wire      [7:0] n9478;
wire      [7:0] n9479;
wire      [7:0] n948;
wire      [7:0] n9480;
wire      [7:0] n9481;
wire      [7:0] n9482;
wire      [7:0] n9483;
wire      [7:0] n9484;
wire      [7:0] n9485;
wire      [7:0] n9486;
wire      [7:0] n9487;
wire      [7:0] n9488;
wire      [7:0] n9489;
wire      [7:0] n949;
wire      [7:0] n9490;
wire      [7:0] n9491;
wire      [7:0] n9492;
wire      [7:0] n9493;
wire      [7:0] n9494;
wire      [7:0] n9495;
wire      [7:0] n9496;
wire      [7:0] n9497;
wire      [7:0] n9498;
wire      [7:0] n9499;
wire      [7:0] n950;
wire      [7:0] n9500;
wire      [7:0] n9501;
wire      [7:0] n9502;
wire      [7:0] n9503;
wire      [7:0] n9504;
wire            n9505;
wire      [7:0] n9506;
wire            n9507;
wire      [7:0] n9508;
wire            n9509;
wire      [7:0] n951;
wire      [7:0] n9510;
wire            n9511;
wire      [7:0] n9512;
wire            n9513;
wire      [7:0] n9514;
wire            n9515;
wire      [7:0] n9516;
wire            n9517;
wire      [7:0] n9518;
wire            n9519;
wire      [7:0] n952;
wire      [7:0] n9520;
wire            n9521;
wire      [7:0] n9522;
wire            n9523;
wire      [7:0] n9524;
wire            n9525;
wire      [7:0] n9526;
wire            n9527;
wire      [7:0] n9528;
wire            n9529;
wire      [7:0] n953;
wire      [7:0] n9530;
wire            n9531;
wire      [7:0] n9532;
wire            n9533;
wire      [7:0] n9534;
wire            n9535;
wire      [7:0] n9536;
wire            n9537;
wire      [7:0] n9538;
wire            n9539;
wire      [7:0] n954;
wire      [7:0] n9540;
wire            n9541;
wire      [7:0] n9542;
wire            n9543;
wire      [7:0] n9544;
wire            n9545;
wire      [7:0] n9546;
wire            n9547;
wire      [7:0] n9548;
wire            n9549;
wire      [7:0] n955;
wire      [7:0] n9550;
wire            n9551;
wire      [7:0] n9552;
wire            n9553;
wire      [7:0] n9554;
wire            n9555;
wire      [7:0] n9556;
wire            n9557;
wire      [7:0] n9558;
wire            n9559;
wire      [7:0] n956;
wire      [7:0] n9560;
wire            n9561;
wire      [7:0] n9562;
wire            n9563;
wire      [7:0] n9564;
wire            n9565;
wire      [7:0] n9566;
wire            n9567;
wire      [7:0] n9568;
wire            n9569;
wire      [7:0] n957;
wire      [7:0] n9570;
wire            n9571;
wire      [7:0] n9572;
wire            n9573;
wire      [7:0] n9574;
wire            n9575;
wire      [7:0] n9576;
wire            n9577;
wire      [7:0] n9578;
wire            n9579;
wire      [7:0] n958;
wire      [7:0] n9580;
wire            n9581;
wire      [7:0] n9582;
wire            n9583;
wire      [7:0] n9584;
wire            n9585;
wire      [7:0] n9586;
wire            n9587;
wire      [7:0] n9588;
wire            n9589;
wire      [7:0] n959;
wire      [7:0] n9590;
wire            n9591;
wire      [7:0] n9592;
wire            n9593;
wire      [7:0] n9594;
wire            n9595;
wire      [7:0] n9596;
wire            n9597;
wire      [7:0] n9598;
wire            n9599;
wire            n96;
wire      [7:0] n960;
wire      [7:0] n9600;
wire            n9601;
wire      [7:0] n9602;
wire            n9603;
wire      [7:0] n9604;
wire            n9605;
wire      [7:0] n9606;
wire            n9607;
wire      [7:0] n9608;
wire            n9609;
wire      [7:0] n961;
wire      [7:0] n9610;
wire            n9611;
wire      [7:0] n9612;
wire            n9613;
wire      [7:0] n9614;
wire            n9615;
wire      [7:0] n9616;
wire            n9617;
wire      [7:0] n9618;
wire            n9619;
wire      [7:0] n962;
wire      [7:0] n9620;
wire            n9621;
wire      [7:0] n9622;
wire            n9623;
wire      [7:0] n9624;
wire            n9625;
wire      [7:0] n9626;
wire            n9627;
wire      [7:0] n9628;
wire            n9629;
wire      [7:0] n963;
wire      [7:0] n9630;
wire            n9631;
wire      [7:0] n9632;
wire            n9633;
wire      [7:0] n9634;
wire            n9635;
wire      [7:0] n9636;
wire            n9637;
wire      [7:0] n9638;
wire            n9639;
wire      [7:0] n964;
wire      [7:0] n9640;
wire            n9641;
wire      [7:0] n9642;
wire            n9643;
wire      [7:0] n9644;
wire            n9645;
wire      [7:0] n9646;
wire            n9647;
wire      [7:0] n9648;
wire            n9649;
wire      [7:0] n965;
wire      [7:0] n9650;
wire            n9651;
wire      [7:0] n9652;
wire            n9653;
wire      [7:0] n9654;
wire            n9655;
wire      [7:0] n9656;
wire            n9657;
wire      [7:0] n9658;
wire            n9659;
wire      [7:0] n966;
wire      [7:0] n9660;
wire            n9661;
wire      [7:0] n9662;
wire            n9663;
wire      [7:0] n9664;
wire            n9665;
wire      [7:0] n9666;
wire            n9667;
wire      [7:0] n9668;
wire            n9669;
wire      [7:0] n967;
wire      [7:0] n9670;
wire            n9671;
wire      [7:0] n9672;
wire            n9673;
wire      [7:0] n9674;
wire            n9675;
wire      [7:0] n9676;
wire            n9677;
wire      [7:0] n9678;
wire            n9679;
wire      [7:0] n968;
wire      [7:0] n9680;
wire            n9681;
wire      [7:0] n9682;
wire            n9683;
wire      [7:0] n9684;
wire            n9685;
wire      [7:0] n9686;
wire            n9687;
wire      [7:0] n9688;
wire            n9689;
wire      [7:0] n969;
wire      [7:0] n9690;
wire            n9691;
wire      [7:0] n9692;
wire            n9693;
wire      [7:0] n9694;
wire            n9695;
wire      [7:0] n9696;
wire            n9697;
wire      [7:0] n9698;
wire            n9699;
wire      [7:0] n970;
wire      [7:0] n9700;
wire            n9701;
wire      [7:0] n9702;
wire            n9703;
wire      [7:0] n9704;
wire            n9705;
wire      [7:0] n9706;
wire            n9707;
wire      [7:0] n9708;
wire            n9709;
wire      [7:0] n971;
wire      [7:0] n9710;
wire            n9711;
wire      [7:0] n9712;
wire            n9713;
wire      [7:0] n9714;
wire            n9715;
wire      [7:0] n9716;
wire            n9717;
wire      [7:0] n9718;
wire            n9719;
wire      [7:0] n972;
wire      [7:0] n9720;
wire            n9721;
wire      [7:0] n9722;
wire            n9723;
wire      [7:0] n9724;
wire            n9725;
wire      [7:0] n9726;
wire            n9727;
wire      [7:0] n9728;
wire            n9729;
wire      [7:0] n973;
wire      [7:0] n9730;
wire            n9731;
wire      [7:0] n9732;
wire            n9733;
wire      [7:0] n9734;
wire            n9735;
wire      [7:0] n9736;
wire            n9737;
wire      [7:0] n9738;
wire            n9739;
wire      [7:0] n974;
wire      [7:0] n9740;
wire            n9741;
wire      [7:0] n9742;
wire            n9743;
wire      [7:0] n9744;
wire            n9745;
wire      [7:0] n9746;
wire            n9747;
wire      [7:0] n9748;
wire            n9749;
wire      [7:0] n975;
wire      [7:0] n9750;
wire            n9751;
wire      [7:0] n9752;
wire            n9753;
wire      [7:0] n9754;
wire            n9755;
wire      [7:0] n9756;
wire            n9757;
wire      [7:0] n9758;
wire            n9759;
wire      [7:0] n976;
wire      [7:0] n9760;
wire            n9761;
wire      [7:0] n9762;
wire            n9763;
wire      [7:0] n9764;
wire            n9765;
wire      [7:0] n9766;
wire            n9767;
wire      [7:0] n9768;
wire            n9769;
wire      [7:0] n977;
wire      [7:0] n9770;
wire            n9771;
wire      [7:0] n9772;
wire            n9773;
wire      [7:0] n9774;
wire            n9775;
wire      [7:0] n9776;
wire            n9777;
wire      [7:0] n9778;
wire            n9779;
wire      [7:0] n978;
wire      [7:0] n9780;
wire            n9781;
wire      [7:0] n9782;
wire            n9783;
wire      [7:0] n9784;
wire            n9785;
wire      [7:0] n9786;
wire            n9787;
wire      [7:0] n9788;
wire            n9789;
wire      [7:0] n979;
wire      [7:0] n9790;
wire            n9791;
wire      [7:0] n9792;
wire            n9793;
wire      [7:0] n9794;
wire            n9795;
wire      [7:0] n9796;
wire            n9797;
wire      [7:0] n9798;
wire            n9799;
wire      [7:0] n98;
wire      [7:0] n980;
wire      [7:0] n9800;
wire            n9801;
wire      [7:0] n9802;
wire            n9803;
wire      [7:0] n9804;
wire            n9805;
wire      [7:0] n9806;
wire            n9807;
wire      [7:0] n9808;
wire            n9809;
wire      [7:0] n981;
wire      [7:0] n9810;
wire            n9811;
wire      [7:0] n9812;
wire            n9813;
wire      [7:0] n9814;
wire            n9815;
wire      [7:0] n9816;
wire            n9817;
wire      [7:0] n9818;
wire            n9819;
wire      [7:0] n982;
wire      [7:0] n9820;
wire            n9821;
wire      [7:0] n9822;
wire            n9823;
wire      [7:0] n9824;
wire            n9825;
wire      [7:0] n9826;
wire            n9827;
wire      [7:0] n9828;
wire            n9829;
wire      [7:0] n983;
wire      [7:0] n9830;
wire            n9831;
wire      [7:0] n9832;
wire            n9833;
wire      [7:0] n9834;
wire            n9835;
wire      [7:0] n9836;
wire            n9837;
wire      [7:0] n9838;
wire            n9839;
wire      [7:0] n984;
wire      [7:0] n9840;
wire            n9841;
wire      [7:0] n9842;
wire            n9843;
wire      [7:0] n9844;
wire            n9845;
wire      [7:0] n9846;
wire            n9847;
wire      [7:0] n9848;
wire            n9849;
wire      [7:0] n985;
wire      [7:0] n9850;
wire            n9851;
wire      [7:0] n9852;
wire            n9853;
wire      [7:0] n9854;
wire            n9855;
wire      [7:0] n9856;
wire            n9857;
wire      [7:0] n9858;
wire            n9859;
wire      [7:0] n986;
wire      [7:0] n9860;
wire            n9861;
wire      [7:0] n9862;
wire            n9863;
wire      [7:0] n9864;
wire            n9865;
wire      [7:0] n9866;
wire            n9867;
wire      [7:0] n9868;
wire            n9869;
wire      [7:0] n987;
wire      [7:0] n9870;
wire            n9871;
wire      [7:0] n9872;
wire            n9873;
wire      [7:0] n9874;
wire            n9875;
wire      [7:0] n9876;
wire            n9877;
wire      [7:0] n9878;
wire            n9879;
wire      [7:0] n988;
wire      [7:0] n9880;
wire            n9881;
wire      [7:0] n9882;
wire            n9883;
wire      [7:0] n9884;
wire            n9885;
wire      [7:0] n9886;
wire            n9887;
wire      [7:0] n9888;
wire            n9889;
wire      [7:0] n989;
wire      [7:0] n9890;
wire            n9891;
wire      [7:0] n9892;
wire            n9893;
wire      [7:0] n9894;
wire            n9895;
wire      [7:0] n9896;
wire            n9897;
wire      [7:0] n9898;
wire            n9899;
wire      [7:0] n990;
wire      [7:0] n9900;
wire            n9901;
wire      [7:0] n9902;
wire            n9903;
wire      [7:0] n9904;
wire            n9905;
wire      [7:0] n9906;
wire            n9907;
wire      [7:0] n9908;
wire            n9909;
wire      [7:0] n991;
wire      [7:0] n9910;
wire            n9911;
wire      [7:0] n9912;
wire            n9913;
wire      [7:0] n9914;
wire            n9915;
wire      [7:0] n9916;
wire            n9917;
wire      [7:0] n9918;
wire            n9919;
wire      [7:0] n992;
wire      [7:0] n9920;
wire            n9921;
wire      [7:0] n9922;
wire            n9923;
wire      [7:0] n9924;
wire            n9925;
wire      [7:0] n9926;
wire            n9927;
wire      [7:0] n9928;
wire            n9929;
wire      [7:0] n993;
wire      [7:0] n9930;
wire            n9931;
wire      [7:0] n9932;
wire            n9933;
wire      [7:0] n9934;
wire            n9935;
wire      [7:0] n9936;
wire            n9937;
wire      [7:0] n9938;
wire            n9939;
wire      [7:0] n994;
wire      [7:0] n9940;
wire            n9941;
wire      [7:0] n9942;
wire            n9943;
wire      [7:0] n9944;
wire            n9945;
wire      [7:0] n9946;
wire            n9947;
wire      [7:0] n9948;
wire            n9949;
wire      [7:0] n995;
wire      [7:0] n9950;
wire            n9951;
wire      [7:0] n9952;
wire            n9953;
wire      [7:0] n9954;
wire            n9955;
wire      [7:0] n9956;
wire            n9957;
wire      [7:0] n9958;
wire            n9959;
wire      [7:0] n996;
wire      [7:0] n9960;
wire            n9961;
wire      [7:0] n9962;
wire            n9963;
wire      [7:0] n9964;
wire            n9965;
wire      [7:0] n9966;
wire            n9967;
wire      [7:0] n9968;
wire            n9969;
wire      [7:0] n997;
wire      [7:0] n9970;
wire            n9971;
wire      [7:0] n9972;
wire            n9973;
wire      [7:0] n9974;
wire            n9975;
wire      [7:0] n9976;
wire            n9977;
wire      [7:0] n9978;
wire            n9979;
wire      [7:0] n998;
wire      [7:0] n9980;
wire            n9981;
wire      [7:0] n9982;
wire            n9983;
wire      [7:0] n9984;
wire            n9985;
wire      [7:0] n9986;
wire            n9987;
wire      [7:0] n9988;
wire            n9989;
wire      [7:0] n999;
wire      [7:0] n9990;
wire            n9991;
wire      [7:0] n9992;
wire            n9993;
wire      [7:0] n9994;
wire            n9995;
wire      [7:0] n9996;
wire            n9997;
wire      [7:0] n9998;
wire            n9999;
wire            rst;
(* keep *) wire    [127:0] state_in_randinit;
(* keep *) wire    [127:0] state_out_randinit;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign bv_128_0_n1 = 128'h0 ;
assign n2 = state_in[127:120] ;
assign bv_8_255_n3 = 8'hff ;
assign n4 =  ( n2 ) == ( bv_8_255_n3 )  ;
assign bv_8_44_n5 = 8'h2c ;
assign n6 = state_in[127:120] ;
assign bv_8_254_n7 = 8'hfe ;
assign n8 =  ( n6 ) == ( bv_8_254_n7 )  ;
assign bv_8_109_n9 = 8'h6d ;
assign n10 = state_in[127:120] ;
assign bv_8_253_n11 = 8'hfd ;
assign n12 =  ( n10 ) == ( bv_8_253_n11 )  ;
assign bv_8_168_n13 = 8'ha8 ;
assign n14 = state_in[127:120] ;
assign bv_8_252_n15 = 8'hfc ;
assign n16 =  ( n14 ) == ( bv_8_252_n15 )  ;
assign bv_8_123_n17 = 8'h7b ;
assign n18 = state_in[127:120] ;
assign bv_8_251_n19 = 8'hfb ;
assign n20 =  ( n18 ) == ( bv_8_251_n19 )  ;
assign bv_8_30_n21 = 8'h1e ;
assign n22 = state_in[127:120] ;
assign bv_8_250_n23 = 8'hfa ;
assign n24 =  ( n22 ) == ( bv_8_250_n23 )  ;
assign bv_8_90_n25 = 8'h5a ;
assign n26 = state_in[127:120] ;
assign bv_8_249_n27 = 8'hf9 ;
assign n28 =  ( n26 ) == ( bv_8_249_n27 )  ;
assign bv_8_41_n29 = 8'h29 ;
assign n30 = state_in[127:120] ;
assign bv_8_248_n31 = 8'hf8 ;
assign n32 =  ( n30 ) == ( bv_8_248_n31 )  ;
assign bv_8_130_n33 = 8'h82 ;
assign n34 = state_in[127:120] ;
assign bv_8_247_n35 = 8'hf7 ;
assign n36 =  ( n34 ) == ( bv_8_247_n35 )  ;
assign bv_8_208_n37 = 8'hd0 ;
assign n38 = state_in[127:120] ;
assign bv_8_246_n39 = 8'hf6 ;
assign n40 =  ( n38 ) == ( bv_8_246_n39 )  ;
assign bv_8_132_n41 = 8'h84 ;
assign n42 = state_in[127:120] ;
assign bv_8_245_n43 = 8'hf5 ;
assign n44 =  ( n42 ) == ( bv_8_245_n43 )  ;
assign bv_8_215_n45 = 8'hd7 ;
assign n46 = state_in[127:120] ;
assign bv_8_244_n47 = 8'hf4 ;
assign n48 =  ( n46 ) == ( bv_8_244_n47 )  ;
assign bv_8_101_n49 = 8'h65 ;
assign n50 = state_in[127:120] ;
assign bv_8_243_n51 = 8'hf3 ;
assign n52 =  ( n50 ) == ( bv_8_243_n51 )  ;
assign bv_8_26_n53 = 8'h1a ;
assign n54 = state_in[127:120] ;
assign bv_8_242_n55 = 8'hf2 ;
assign n56 =  ( n54 ) == ( bv_8_242_n55 )  ;
assign bv_8_9_n57 = 8'h9 ;
assign n58 = state_in[127:120] ;
assign bv_8_241_n59 = 8'hf1 ;
assign n60 =  ( n58 ) == ( bv_8_241_n59 )  ;
assign bv_8_89_n61 = 8'h59 ;
assign n62 = state_in[127:120] ;
assign bv_8_240_n63 = 8'hf0 ;
assign n64 =  ( n62 ) == ( bv_8_240_n63 )  ;
assign bv_8_3_n65 = 8'h3 ;
assign n66 = state_in[127:120] ;
assign bv_8_239_n67 = 8'hef ;
assign n68 =  ( n66 ) == ( bv_8_239_n67 )  ;
assign bv_8_165_n69 = 8'ha5 ;
assign n70 = state_in[127:120] ;
assign bv_8_238_n71 = 8'hee ;
assign n72 =  ( n70 ) == ( bv_8_238_n71 )  ;
assign bv_8_80_n73 = 8'h50 ;
assign n74 = state_in[127:120] ;
assign bv_8_237_n75 = 8'hed ;
assign n76 =  ( n74 ) == ( bv_8_237_n75 )  ;
assign bv_8_170_n77 = 8'haa ;
assign n78 = state_in[127:120] ;
assign bv_8_236_n79 = 8'hec ;
assign n80 =  ( n78 ) == ( bv_8_236_n79 )  ;
assign bv_8_135_n81 = 8'h87 ;
assign n82 = state_in[127:120] ;
assign bv_8_235_n83 = 8'heb ;
assign n84 =  ( n82 ) == ( bv_8_235_n83 )  ;
assign bv_8_201_n85 = 8'hc9 ;
assign n86 = state_in[127:120] ;
assign bv_8_234_n87 = 8'hea ;
assign n88 =  ( n86 ) == ( bv_8_234_n87 )  ;
assign bv_8_21_n89 = 8'h15 ;
assign n90 = state_in[127:120] ;
assign bv_8_233_n91 = 8'he9 ;
assign n92 =  ( n90 ) == ( bv_8_233_n91 )  ;
assign bv_8_60_n93 = 8'h3c ;
assign n94 = state_in[127:120] ;
assign bv_8_232_n95 = 8'he8 ;
assign n96 =  ( n94 ) == ( bv_8_232_n95 )  ;
assign bv_8_45_n97 = 8'h2d ;
assign n98 = state_in[127:120] ;
assign bv_8_231_n99 = 8'he7 ;
assign n100 =  ( n98 ) == ( bv_8_231_n99 )  ;
assign bv_8_51_n101 = 8'h33 ;
assign n102 = state_in[127:120] ;
assign bv_8_230_n103 = 8'he6 ;
assign n104 =  ( n102 ) == ( bv_8_230_n103 )  ;
assign bv_8_7_n105 = 8'h7 ;
assign n106 = state_in[127:120] ;
assign bv_8_229_n107 = 8'he5 ;
assign n108 =  ( n106 ) == ( bv_8_229_n107 )  ;
assign bv_8_169_n109 = 8'ha9 ;
assign n110 = state_in[127:120] ;
assign bv_8_228_n111 = 8'he4 ;
assign n112 =  ( n110 ) == ( bv_8_228_n111 )  ;
assign bv_8_210_n113 = 8'hd2 ;
assign n114 = state_in[127:120] ;
assign bv_8_227_n115 = 8'he3 ;
assign n116 =  ( n114 ) == ( bv_8_227_n115 )  ;
assign bv_8_34_n117 = 8'h22 ;
assign n118 = state_in[127:120] ;
assign bv_8_226_n119 = 8'he2 ;
assign n120 =  ( n118 ) == ( bv_8_226_n119 )  ;
assign bv_8_43_n121 = 8'h2b ;
assign n122 = state_in[127:120] ;
assign bv_8_225_n123 = 8'he1 ;
assign n124 =  ( n122 ) == ( bv_8_225_n123 )  ;
assign n125 = state_in[127:120] ;
assign bv_8_224_n126 = 8'he0 ;
assign n127 =  ( n125 ) == ( bv_8_224_n126 )  ;
assign bv_8_217_n128 = 8'hd9 ;
assign n129 = state_in[127:120] ;
assign bv_8_223_n130 = 8'hdf ;
assign n131 =  ( n129 ) == ( bv_8_223_n130 )  ;
assign bv_8_39_n132 = 8'h27 ;
assign n133 = state_in[127:120] ;
assign bv_8_222_n134 = 8'hde ;
assign n135 =  ( n133 ) == ( bv_8_222_n134 )  ;
assign bv_8_58_n136 = 8'h3a ;
assign n137 = state_in[127:120] ;
assign bv_8_221_n138 = 8'hdd ;
assign n139 =  ( n137 ) == ( bv_8_221_n138 )  ;
assign bv_8_153_n140 = 8'h99 ;
assign n141 = state_in[127:120] ;
assign bv_8_220_n142 = 8'hdc ;
assign n143 =  ( n141 ) == ( bv_8_220_n142 )  ;
assign bv_8_23_n144 = 8'h17 ;
assign n145 = state_in[127:120] ;
assign bv_8_219_n146 = 8'hdb ;
assign n147 =  ( n145 ) == ( bv_8_219_n146 )  ;
assign bv_8_105_n148 = 8'h69 ;
assign n149 = state_in[127:120] ;
assign bv_8_218_n150 = 8'hda ;
assign n151 =  ( n149 ) == ( bv_8_218_n150 )  ;
assign bv_8_174_n152 = 8'hae ;
assign n153 = state_in[127:120] ;
assign n154 =  ( n153 ) == ( bv_8_217_n128 )  ;
assign bv_8_106_n155 = 8'h6a ;
assign n156 = state_in[127:120] ;
assign bv_8_216_n157 = 8'hd8 ;
assign n158 =  ( n156 ) == ( bv_8_216_n157 )  ;
assign bv_8_194_n159 = 8'hc2 ;
assign n160 = state_in[127:120] ;
assign n161 =  ( n160 ) == ( bv_8_215_n45 )  ;
assign bv_8_28_n162 = 8'h1c ;
assign n163 = state_in[127:120] ;
assign bv_8_214_n164 = 8'hd6 ;
assign n165 =  ( n163 ) == ( bv_8_214_n164 )  ;
assign n166 = state_in[127:120] ;
assign bv_8_213_n167 = 8'hd5 ;
assign n168 =  ( n166 ) == ( bv_8_213_n167 )  ;
assign bv_8_6_n169 = 8'h6 ;
assign n170 = state_in[127:120] ;
assign bv_8_212_n171 = 8'hd4 ;
assign n172 =  ( n170 ) == ( bv_8_212_n171 )  ;
assign bv_8_144_n173 = 8'h90 ;
assign n174 = state_in[127:120] ;
assign bv_8_211_n175 = 8'hd3 ;
assign n176 =  ( n174 ) == ( bv_8_211_n175 )  ;
assign bv_8_204_n177 = 8'hcc ;
assign n178 = state_in[127:120] ;
assign n179 =  ( n178 ) == ( bv_8_210_n113 )  ;
assign bv_8_113_n180 = 8'h71 ;
assign n181 = state_in[127:120] ;
assign bv_8_209_n182 = 8'hd1 ;
assign n183 =  ( n181 ) == ( bv_8_209_n182 )  ;
assign bv_8_124_n184 = 8'h7c ;
assign n185 = state_in[127:120] ;
assign n186 =  ( n185 ) == ( bv_8_208_n37 )  ;
assign n187 = state_in[127:120] ;
assign bv_8_207_n188 = 8'hcf ;
assign n189 =  ( n187 ) == ( bv_8_207_n188 )  ;
assign bv_8_15_n190 = 8'hf ;
assign n191 = state_in[127:120] ;
assign bv_8_206_n192 = 8'hce ;
assign n193 =  ( n191 ) == ( bv_8_206_n192 )  ;
assign bv_8_13_n194 = 8'hd ;
assign n195 = state_in[127:120] ;
assign bv_8_205_n196 = 8'hcd ;
assign n197 =  ( n195 ) == ( bv_8_205_n196 )  ;
assign bv_8_97_n198 = 8'h61 ;
assign n199 = state_in[127:120] ;
assign n200 =  ( n199 ) == ( bv_8_204_n177 )  ;
assign bv_8_150_n201 = 8'h96 ;
assign n202 = state_in[127:120] ;
assign bv_8_203_n203 = 8'hcb ;
assign n204 =  ( n202 ) == ( bv_8_203_n203 )  ;
assign bv_8_62_n205 = 8'h3e ;
assign n206 = state_in[127:120] ;
assign bv_8_202_n207 = 8'hca ;
assign n208 =  ( n206 ) == ( bv_8_202_n207 )  ;
assign n209 = state_in[127:120] ;
assign n210 =  ( n209 ) == ( bv_8_201_n85 )  ;
assign bv_8_161_n211 = 8'ha1 ;
assign n212 = state_in[127:120] ;
assign bv_8_200_n213 = 8'hc8 ;
assign n214 =  ( n212 ) == ( bv_8_200_n213 )  ;
assign n215 = state_in[127:120] ;
assign bv_8_199_n216 = 8'hc7 ;
assign n217 =  ( n215 ) == ( bv_8_199_n216 )  ;
assign bv_8_151_n218 = 8'h97 ;
assign n219 = state_in[127:120] ;
assign bv_8_198_n220 = 8'hc6 ;
assign n221 =  ( n219 ) == ( bv_8_198_n220 )  ;
assign bv_8_115_n222 = 8'h73 ;
assign n223 = state_in[127:120] ;
assign bv_8_197_n224 = 8'hc5 ;
assign n225 =  ( n223 ) == ( bv_8_197_n224 )  ;
assign bv_8_87_n226 = 8'h57 ;
assign n227 = state_in[127:120] ;
assign bv_8_196_n228 = 8'hc4 ;
assign n229 =  ( n227 ) == ( bv_8_196_n228 )  ;
assign bv_8_56_n230 = 8'h38 ;
assign n231 = state_in[127:120] ;
assign bv_8_195_n232 = 8'hc3 ;
assign n233 =  ( n231 ) == ( bv_8_195_n232 )  ;
assign bv_8_92_n234 = 8'h5c ;
assign n235 = state_in[127:120] ;
assign n236 =  ( n235 ) == ( bv_8_194_n159 )  ;
assign bv_8_74_n237 = 8'h4a ;
assign n238 = state_in[127:120] ;
assign bv_8_193_n239 = 8'hc1 ;
assign n240 =  ( n238 ) == ( bv_8_193_n239 )  ;
assign n241 = state_in[127:120] ;
assign bv_8_192_n242 = 8'hc0 ;
assign n243 =  ( n241 ) == ( bv_8_192_n242 )  ;
assign bv_8_111_n244 = 8'h6f ;
assign n245 = state_in[127:120] ;
assign bv_8_191_n246 = 8'hbf ;
assign n247 =  ( n245 ) == ( bv_8_191_n246 )  ;
assign bv_8_16_n248 = 8'h10 ;
assign n249 = state_in[127:120] ;
assign bv_8_190_n250 = 8'hbe ;
assign n251 =  ( n249 ) == ( bv_8_190_n250 )  ;
assign bv_8_71_n252 = 8'h47 ;
assign n253 = state_in[127:120] ;
assign bv_8_189_n254 = 8'hbd ;
assign n255 =  ( n253 ) == ( bv_8_189_n254 )  ;
assign n256 = state_in[127:120] ;
assign bv_8_188_n257 = 8'hbc ;
assign n258 =  ( n256 ) == ( bv_8_188_n257 )  ;
assign n259 = state_in[127:120] ;
assign bv_8_187_n260 = 8'hbb ;
assign n261 =  ( n259 ) == ( bv_8_187_n260 )  ;
assign n262 = state_in[127:120] ;
assign bv_8_186_n263 = 8'hba ;
assign n264 =  ( n262 ) == ( bv_8_186_n263 )  ;
assign n265 = state_in[127:120] ;
assign bv_8_185_n266 = 8'hb9 ;
assign n267 =  ( n265 ) == ( bv_8_185_n266 )  ;
assign bv_8_172_n268 = 8'hac ;
assign n269 = state_in[127:120] ;
assign bv_8_184_n270 = 8'hb8 ;
assign n271 =  ( n269 ) == ( bv_8_184_n270 )  ;
assign n272 = state_in[127:120] ;
assign bv_8_183_n273 = 8'hb7 ;
assign n274 =  ( n272 ) == ( bv_8_183_n273 )  ;
assign bv_8_73_n275 = 8'h49 ;
assign n276 = state_in[127:120] ;
assign bv_8_182_n277 = 8'hb6 ;
assign n278 =  ( n276 ) == ( bv_8_182_n277 )  ;
assign bv_8_156_n279 = 8'h9c ;
assign n280 = state_in[127:120] ;
assign bv_8_181_n281 = 8'hb5 ;
assign n282 =  ( n280 ) == ( bv_8_181_n281 )  ;
assign bv_8_177_n283 = 8'hb1 ;
assign n284 = state_in[127:120] ;
assign bv_8_180_n285 = 8'hb4 ;
assign n286 =  ( n284 ) == ( bv_8_180_n285 )  ;
assign bv_8_1_n287 = 8'h1 ;
assign n288 = state_in[127:120] ;
assign bv_8_179_n289 = 8'hb3 ;
assign n290 =  ( n288 ) == ( bv_8_179_n289 )  ;
assign n291 = state_in[127:120] ;
assign bv_8_178_n292 = 8'hb2 ;
assign n293 =  ( n291 ) == ( bv_8_178_n292 )  ;
assign bv_8_110_n294 = 8'h6e ;
assign n295 = state_in[127:120] ;
assign n296 =  ( n295 ) == ( bv_8_177_n283 )  ;
assign bv_8_139_n297 = 8'h8b ;
assign n298 = state_in[127:120] ;
assign bv_8_176_n299 = 8'hb0 ;
assign n300 =  ( n298 ) == ( bv_8_176_n299 )  ;
assign n301 = state_in[127:120] ;
assign bv_8_175_n302 = 8'haf ;
assign n303 =  ( n301 ) == ( bv_8_175_n302 )  ;
assign n304 = state_in[127:120] ;
assign n305 =  ( n304 ) == ( bv_8_174_n152 )  ;
assign n306 = state_in[127:120] ;
assign bv_8_173_n307 = 8'had ;
assign n308 =  ( n306 ) == ( bv_8_173_n307 )  ;
assign bv_8_49_n309 = 8'h31 ;
assign n310 = state_in[127:120] ;
assign n311 =  ( n310 ) == ( bv_8_172_n268 )  ;
assign bv_8_57_n312 = 8'h39 ;
assign n313 = state_in[127:120] ;
assign bv_8_171_n314 = 8'hab ;
assign n315 =  ( n313 ) == ( bv_8_171_n314 )  ;
assign n316 = state_in[127:120] ;
assign n317 =  ( n316 ) == ( bv_8_170_n77 )  ;
assign bv_8_67_n318 = 8'h43 ;
assign n319 = state_in[127:120] ;
assign n320 =  ( n319 ) == ( bv_8_169_n109 )  ;
assign n321 = state_in[127:120] ;
assign n322 =  ( n321 ) == ( bv_8_168_n13 )  ;
assign bv_8_159_n323 = 8'h9f ;
assign n324 = state_in[127:120] ;
assign bv_8_167_n325 = 8'ha7 ;
assign n326 =  ( n324 ) == ( bv_8_167_n325 )  ;
assign n327 = state_in[127:120] ;
assign bv_8_166_n328 = 8'ha6 ;
assign n329 =  ( n327 ) == ( bv_8_166_n328 )  ;
assign bv_8_72_n330 = 8'h48 ;
assign n331 = state_in[127:120] ;
assign n332 =  ( n331 ) == ( bv_8_165_n69 )  ;
assign bv_8_12_n333 = 8'hc ;
assign n334 = state_in[127:120] ;
assign bv_8_164_n335 = 8'ha4 ;
assign n336 =  ( n334 ) == ( bv_8_164_n335 )  ;
assign bv_8_146_n337 = 8'h92 ;
assign n338 = state_in[127:120] ;
assign bv_8_163_n339 = 8'ha3 ;
assign n340 =  ( n338 ) == ( bv_8_163_n339 )  ;
assign bv_8_20_n341 = 8'h14 ;
assign n342 = state_in[127:120] ;
assign bv_8_162_n343 = 8'ha2 ;
assign n344 =  ( n342 ) == ( bv_8_162_n343 )  ;
assign bv_8_116_n345 = 8'h74 ;
assign n346 = state_in[127:120] ;
assign n347 =  ( n346 ) == ( bv_8_161_n211 )  ;
assign bv_8_100_n348 = 8'h64 ;
assign n349 = state_in[127:120] ;
assign bv_8_160_n350 = 8'ha0 ;
assign n351 =  ( n349 ) == ( bv_8_160_n350 )  ;
assign n352 = state_in[127:120] ;
assign n353 =  ( n352 ) == ( bv_8_159_n323 )  ;
assign n354 = state_in[127:120] ;
assign bv_8_158_n355 = 8'h9e ;
assign n356 =  ( n354 ) == ( bv_8_158_n355 )  ;
assign bv_8_22_n357 = 8'h16 ;
assign n358 = state_in[127:120] ;
assign bv_8_157_n359 = 8'h9d ;
assign n360 =  ( n358 ) == ( bv_8_157_n359 )  ;
assign n361 = state_in[127:120] ;
assign n362 =  ( n361 ) == ( bv_8_156_n279 )  ;
assign n363 = state_in[127:120] ;
assign bv_8_155_n364 = 8'h9b ;
assign n365 =  ( n363 ) == ( bv_8_155_n364 )  ;
assign bv_8_40_n366 = 8'h28 ;
assign n367 = state_in[127:120] ;
assign bv_8_154_n368 = 8'h9a ;
assign n369 =  ( n367 ) == ( bv_8_154_n368 )  ;
assign bv_8_107_n370 = 8'h6b ;
assign n371 = state_in[127:120] ;
assign n372 =  ( n371 ) == ( bv_8_153_n140 )  ;
assign n373 = state_in[127:120] ;
assign bv_8_152_n374 = 8'h98 ;
assign n375 =  ( n373 ) == ( bv_8_152_n374 )  ;
assign bv_8_140_n376 = 8'h8c ;
assign n377 = state_in[127:120] ;
assign n378 =  ( n377 ) == ( bv_8_151_n218 )  ;
assign bv_8_11_n379 = 8'hb ;
assign n380 = state_in[127:120] ;
assign n381 =  ( n380 ) == ( bv_8_150_n201 )  ;
assign bv_8_59_n382 = 8'h3b ;
assign n383 = state_in[127:120] ;
assign bv_8_149_n384 = 8'h95 ;
assign n385 =  ( n383 ) == ( bv_8_149_n384 )  ;
assign bv_8_84_n386 = 8'h54 ;
assign n387 = state_in[127:120] ;
assign bv_8_148_n388 = 8'h94 ;
assign n389 =  ( n387 ) == ( bv_8_148_n388 )  ;
assign bv_8_68_n390 = 8'h44 ;
assign n391 = state_in[127:120] ;
assign bv_8_147_n392 = 8'h93 ;
assign n393 =  ( n391 ) == ( bv_8_147_n392 )  ;
assign n394 = state_in[127:120] ;
assign n395 =  ( n394 ) == ( bv_8_146_n337 )  ;
assign n396 = state_in[127:120] ;
assign bv_8_145_n397 = 8'h91 ;
assign n398 =  ( n396 ) == ( bv_8_145_n397 )  ;
assign bv_8_25_n399 = 8'h19 ;
assign n400 = state_in[127:120] ;
assign n401 =  ( n400 ) == ( bv_8_144_n173 )  ;
assign n402 = state_in[127:120] ;
assign bv_8_143_n403 = 8'h8f ;
assign n404 =  ( n402 ) == ( bv_8_143_n403 )  ;
assign n405 = state_in[127:120] ;
assign bv_8_142_n406 = 8'h8e ;
assign n407 =  ( n405 ) == ( bv_8_142_n406 )  ;
assign bv_8_50_n408 = 8'h32 ;
assign n409 = state_in[127:120] ;
assign bv_8_141_n410 = 8'h8d ;
assign n411 =  ( n409 ) == ( bv_8_141_n410 )  ;
assign n412 = state_in[127:120] ;
assign n413 =  ( n412 ) == ( bv_8_140_n376 )  ;
assign n414 = state_in[127:120] ;
assign n415 =  ( n414 ) == ( bv_8_139_n297 )  ;
assign bv_8_122_n416 = 8'h7a ;
assign n417 = state_in[127:120] ;
assign bv_8_138_n418 = 8'h8a ;
assign n419 =  ( n417 ) == ( bv_8_138_n418 )  ;
assign n420 = state_in[127:120] ;
assign bv_8_137_n421 = 8'h89 ;
assign n422 =  ( n420 ) == ( bv_8_137_n421 )  ;
assign bv_8_85_n423 = 8'h55 ;
assign n424 = state_in[127:120] ;
assign bv_8_136_n425 = 8'h88 ;
assign n426 =  ( n424 ) == ( bv_8_136_n425 )  ;
assign n427 = state_in[127:120] ;
assign n428 =  ( n427 ) == ( bv_8_135_n81 )  ;
assign bv_8_46_n429 = 8'h2e ;
assign n430 = state_in[127:120] ;
assign bv_8_134_n431 = 8'h86 ;
assign n432 =  ( n430 ) == ( bv_8_134_n431 )  ;
assign n433 = state_in[127:120] ;
assign bv_8_133_n434 = 8'h85 ;
assign n435 =  ( n433 ) == ( bv_8_133_n434 )  ;
assign bv_8_53_n436 = 8'h35 ;
assign n437 = state_in[127:120] ;
assign n438 =  ( n437 ) == ( bv_8_132_n41 )  ;
assign n439 = state_in[127:120] ;
assign bv_8_131_n440 = 8'h83 ;
assign n441 =  ( n439 ) == ( bv_8_131_n440 )  ;
assign n442 = state_in[127:120] ;
assign n443 =  ( n442 ) == ( bv_8_130_n33 )  ;
assign bv_8_38_n444 = 8'h26 ;
assign n445 = state_in[127:120] ;
assign bv_8_129_n446 = 8'h81 ;
assign n447 =  ( n445 ) == ( bv_8_129_n446 )  ;
assign bv_8_24_n448 = 8'h18 ;
assign n449 = state_in[127:120] ;
assign bv_8_128_n450 = 8'h80 ;
assign n451 =  ( n449 ) == ( bv_8_128_n450 )  ;
assign n452 = state_in[127:120] ;
assign bv_8_127_n453 = 8'h7f ;
assign n454 =  ( n452 ) == ( bv_8_127_n453 )  ;
assign n455 = state_in[127:120] ;
assign bv_8_126_n456 = 8'h7e ;
assign n457 =  ( n455 ) == ( bv_8_126_n456 )  ;
assign n458 = state_in[127:120] ;
assign bv_8_125_n459 = 8'h7d ;
assign n460 =  ( n458 ) == ( bv_8_125_n459 )  ;
assign n461 = state_in[127:120] ;
assign n462 =  ( n461 ) == ( bv_8_124_n184 )  ;
assign bv_8_32_n463 = 8'h20 ;
assign n464 = state_in[127:120] ;
assign n465 =  ( n464 ) == ( bv_8_123_n17 )  ;
assign bv_8_66_n466 = 8'h42 ;
assign n467 = state_in[127:120] ;
assign n468 =  ( n467 ) == ( bv_8_122_n416 )  ;
assign n469 = state_in[127:120] ;
assign bv_8_121_n470 = 8'h79 ;
assign n471 =  ( n469 ) == ( bv_8_121_n470 )  ;
assign bv_8_119_n472 = 8'h77 ;
assign n473 = state_in[127:120] ;
assign bv_8_120_n474 = 8'h78 ;
assign n475 =  ( n473 ) == ( bv_8_120_n474 )  ;
assign bv_8_99_n476 = 8'h63 ;
assign n477 = state_in[127:120] ;
assign n478 =  ( n477 ) == ( bv_8_119_n472 )  ;
assign n479 = state_in[127:120] ;
assign bv_8_118_n480 = 8'h76 ;
assign n481 =  ( n479 ) == ( bv_8_118_n480 )  ;
assign bv_8_112_n482 = 8'h70 ;
assign n483 = state_in[127:120] ;
assign bv_8_117_n484 = 8'h75 ;
assign n485 =  ( n483 ) == ( bv_8_117_n484 )  ;
assign bv_8_33_n486 = 8'h21 ;
assign n487 = state_in[127:120] ;
assign n488 =  ( n487 ) == ( bv_8_116_n345 )  ;
assign bv_8_63_n489 = 8'h3f ;
assign n490 = state_in[127:120] ;
assign n491 =  ( n490 ) == ( bv_8_115_n222 )  ;
assign bv_8_5_n492 = 8'h5 ;
assign n493 = state_in[127:120] ;
assign bv_8_114_n494 = 8'h72 ;
assign n495 =  ( n493 ) == ( bv_8_114_n494 )  ;
assign n496 = state_in[127:120] ;
assign n497 =  ( n496 ) == ( bv_8_113_n180 )  ;
assign bv_8_93_n498 = 8'h5d ;
assign n499 = state_in[127:120] ;
assign n500 =  ( n499 ) == ( bv_8_112_n482 )  ;
assign n501 = state_in[127:120] ;
assign n502 =  ( n501 ) == ( bv_8_111_n244 )  ;
assign bv_8_75_n503 = 8'h4b ;
assign n504 = state_in[127:120] ;
assign n505 =  ( n504 ) == ( bv_8_110_n294 )  ;
assign bv_8_37_n506 = 8'h25 ;
assign n507 = state_in[127:120] ;
assign n508 =  ( n507 ) == ( bv_8_109_n9 )  ;
assign n509 = state_in[127:120] ;
assign bv_8_108_n510 = 8'h6c ;
assign n511 =  ( n509 ) == ( bv_8_108_n510 )  ;
assign n512 = state_in[127:120] ;
assign n513 =  ( n512 ) == ( bv_8_107_n370 )  ;
assign n514 = state_in[127:120] ;
assign n515 =  ( n514 ) == ( bv_8_106_n155 )  ;
assign bv_8_4_n516 = 8'h4 ;
assign n517 = state_in[127:120] ;
assign n518 =  ( n517 ) == ( bv_8_105_n148 )  ;
assign n519 = state_in[127:120] ;
assign bv_8_104_n520 = 8'h68 ;
assign n521 =  ( n519 ) == ( bv_8_104_n520 )  ;
assign n522 = state_in[127:120] ;
assign bv_8_103_n523 = 8'h67 ;
assign n524 =  ( n522 ) == ( bv_8_103_n523 )  ;
assign bv_8_17_n525 = 8'h11 ;
assign n526 = state_in[127:120] ;
assign bv_8_102_n527 = 8'h66 ;
assign n528 =  ( n526 ) == ( bv_8_102_n527 )  ;
assign n529 = state_in[127:120] ;
assign n530 =  ( n529 ) == ( bv_8_101_n49 )  ;
assign n531 = state_in[127:120] ;
assign n532 =  ( n531 ) == ( bv_8_100_n348 )  ;
assign n533 = state_in[127:120] ;
assign n534 =  ( n533 ) == ( bv_8_99_n476 )  ;
assign n535 = state_in[127:120] ;
assign bv_8_98_n536 = 8'h62 ;
assign n537 =  ( n535 ) == ( bv_8_98_n536 )  ;
assign bv_8_79_n538 = 8'h4f ;
assign n539 = state_in[127:120] ;
assign n540 =  ( n539 ) == ( bv_8_97_n198 )  ;
assign n541 = state_in[127:120] ;
assign bv_8_96_n542 = 8'h60 ;
assign n543 =  ( n541 ) == ( bv_8_96_n542 )  ;
assign n544 = state_in[127:120] ;
assign bv_8_95_n545 = 8'h5f ;
assign n546 =  ( n544 ) == ( bv_8_95_n545 )  ;
assign n547 = state_in[127:120] ;
assign bv_8_94_n548 = 8'h5e ;
assign n549 =  ( n547 ) == ( bv_8_94_n548 )  ;
assign n550 = state_in[127:120] ;
assign n551 =  ( n550 ) == ( bv_8_93_n498 )  ;
assign n552 = state_in[127:120] ;
assign n553 =  ( n552 ) == ( bv_8_92_n234 )  ;
assign n554 = state_in[127:120] ;
assign bv_8_91_n555 = 8'h5b ;
assign n556 =  ( n554 ) == ( bv_8_91_n555 )  ;
assign n557 = state_in[127:120] ;
assign n558 =  ( n557 ) == ( bv_8_90_n25 )  ;
assign n559 = state_in[127:120] ;
assign n560 =  ( n559 ) == ( bv_8_89_n61 )  ;
assign n561 = state_in[127:120] ;
assign bv_8_88_n562 = 8'h58 ;
assign n563 =  ( n561 ) == ( bv_8_88_n562 )  ;
assign n564 = state_in[127:120] ;
assign n565 =  ( n564 ) == ( bv_8_87_n226 )  ;
assign n566 = state_in[127:120] ;
assign bv_8_86_n567 = 8'h56 ;
assign n568 =  ( n566 ) == ( bv_8_86_n567 )  ;
assign n569 = state_in[127:120] ;
assign n570 =  ( n569 ) == ( bv_8_85_n423 )  ;
assign n571 = state_in[127:120] ;
assign n572 =  ( n571 ) == ( bv_8_84_n386 )  ;
assign bv_8_64_n573 = 8'h40 ;
assign n574 = state_in[127:120] ;
assign bv_8_83_n575 = 8'h53 ;
assign n576 =  ( n574 ) == ( bv_8_83_n575 )  ;
assign n577 = state_in[127:120] ;
assign bv_8_82_n578 = 8'h52 ;
assign n579 =  ( n577 ) == ( bv_8_82_n578 )  ;
assign bv_8_0_n580 = 8'h0 ;
assign n581 = state_in[127:120] ;
assign bv_8_81_n582 = 8'h51 ;
assign n583 =  ( n581 ) == ( bv_8_81_n582 )  ;
assign n584 = state_in[127:120] ;
assign n585 =  ( n584 ) == ( bv_8_80_n73 )  ;
assign n586 = state_in[127:120] ;
assign n587 =  ( n586 ) == ( bv_8_79_n538 )  ;
assign bv_8_19_n588 = 8'h13 ;
assign n589 = state_in[127:120] ;
assign bv_8_78_n590 = 8'h4e ;
assign n591 =  ( n589 ) == ( bv_8_78_n590 )  ;
assign n592 = state_in[127:120] ;
assign bv_8_77_n593 = 8'h4d ;
assign n594 =  ( n592 ) == ( bv_8_77_n593 )  ;
assign n595 = state_in[127:120] ;
assign bv_8_76_n596 = 8'h4c ;
assign n597 =  ( n595 ) == ( bv_8_76_n596 )  ;
assign n598 = state_in[127:120] ;
assign n599 =  ( n598 ) == ( bv_8_75_n503 )  ;
assign n600 = state_in[127:120] ;
assign n601 =  ( n600 ) == ( bv_8_74_n237 )  ;
assign n602 = state_in[127:120] ;
assign n603 =  ( n602 ) == ( bv_8_73_n275 )  ;
assign n604 = state_in[127:120] ;
assign n605 =  ( n604 ) == ( bv_8_72_n330 )  ;
assign n606 = state_in[127:120] ;
assign n607 =  ( n606 ) == ( bv_8_71_n252 )  ;
assign n608 = state_in[127:120] ;
assign bv_8_70_n609 = 8'h46 ;
assign n610 =  ( n608 ) == ( bv_8_70_n609 )  ;
assign n611 = state_in[127:120] ;
assign bv_8_69_n612 = 8'h45 ;
assign n613 =  ( n611 ) == ( bv_8_69_n612 )  ;
assign n614 = state_in[127:120] ;
assign n615 =  ( n614 ) == ( bv_8_68_n390 )  ;
assign bv_8_54_n616 = 8'h36 ;
assign n617 = state_in[127:120] ;
assign n618 =  ( n617 ) == ( bv_8_67_n318 )  ;
assign bv_8_52_n619 = 8'h34 ;
assign n620 = state_in[127:120] ;
assign n621 =  ( n620 ) == ( bv_8_66_n466 )  ;
assign n622 = state_in[127:120] ;
assign bv_8_65_n623 = 8'h41 ;
assign n624 =  ( n622 ) == ( bv_8_65_n623 )  ;
assign bv_8_29_n625 = 8'h1d ;
assign n626 = state_in[127:120] ;
assign n627 =  ( n626 ) == ( bv_8_64_n573 )  ;
assign bv_8_18_n628 = 8'h12 ;
assign n629 = state_in[127:120] ;
assign n630 =  ( n629 ) == ( bv_8_63_n489 )  ;
assign n631 = state_in[127:120] ;
assign n632 =  ( n631 ) == ( bv_8_62_n205 )  ;
assign n633 = state_in[127:120] ;
assign bv_8_61_n634 = 8'h3d ;
assign n635 =  ( n633 ) == ( bv_8_61_n634 )  ;
assign n636 = state_in[127:120] ;
assign n637 =  ( n636 ) == ( bv_8_60_n93 )  ;
assign n638 = state_in[127:120] ;
assign n639 =  ( n638 ) == ( bv_8_59_n382 )  ;
assign n640 = state_in[127:120] ;
assign n641 =  ( n640 ) == ( bv_8_58_n136 )  ;
assign bv_8_27_n642 = 8'h1b ;
assign n643 = state_in[127:120] ;
assign n644 =  ( n643 ) == ( bv_8_57_n312 )  ;
assign bv_8_36_n645 = 8'h24 ;
assign n646 = state_in[127:120] ;
assign n647 =  ( n646 ) == ( bv_8_56_n230 )  ;
assign bv_8_14_n648 = 8'he ;
assign n649 = state_in[127:120] ;
assign bv_8_55_n650 = 8'h37 ;
assign n651 =  ( n649 ) == ( bv_8_55_n650 )  ;
assign bv_8_47_n652 = 8'h2f ;
assign n653 = state_in[127:120] ;
assign n654 =  ( n653 ) == ( bv_8_54_n616 )  ;
assign bv_8_10_n655 = 8'ha ;
assign n656 = state_in[127:120] ;
assign n657 =  ( n656 ) == ( bv_8_53_n436 )  ;
assign n658 = state_in[127:120] ;
assign n659 =  ( n658 ) == ( bv_8_52_n619 )  ;
assign bv_8_48_n660 = 8'h30 ;
assign n661 = state_in[127:120] ;
assign n662 =  ( n661 ) == ( bv_8_51_n101 )  ;
assign n663 = state_in[127:120] ;
assign n664 =  ( n663 ) == ( bv_8_50_n408 )  ;
assign n665 = state_in[127:120] ;
assign n666 =  ( n665 ) == ( bv_8_49_n309 )  ;
assign n667 = state_in[127:120] ;
assign n668 =  ( n667 ) == ( bv_8_48_n660 )  ;
assign bv_8_8_n669 = 8'h8 ;
assign n670 = state_in[127:120] ;
assign n671 =  ( n670 ) == ( bv_8_47_n652 )  ;
assign bv_8_42_n672 = 8'h2a ;
assign n673 = state_in[127:120] ;
assign n674 =  ( n673 ) == ( bv_8_46_n429 )  ;
assign n675 = state_in[127:120] ;
assign n676 =  ( n675 ) == ( bv_8_45_n97 )  ;
assign n677 = state_in[127:120] ;
assign n678 =  ( n677 ) == ( bv_8_44_n5 )  ;
assign n679 = state_in[127:120] ;
assign n680 =  ( n679 ) == ( bv_8_43_n121 )  ;
assign n681 = state_in[127:120] ;
assign n682 =  ( n681 ) == ( bv_8_42_n672 )  ;
assign n683 = state_in[127:120] ;
assign n684 =  ( n683 ) == ( bv_8_41_n29 )  ;
assign n685 = state_in[127:120] ;
assign n686 =  ( n685 ) == ( bv_8_40_n366 )  ;
assign n687 = state_in[127:120] ;
assign n688 =  ( n687 ) == ( bv_8_39_n132 )  ;
assign n689 = state_in[127:120] ;
assign n690 =  ( n689 ) == ( bv_8_38_n444 )  ;
assign n691 = state_in[127:120] ;
assign n692 =  ( n691 ) == ( bv_8_37_n506 )  ;
assign n693 = state_in[127:120] ;
assign n694 =  ( n693 ) == ( bv_8_36_n645 )  ;
assign n695 = state_in[127:120] ;
assign bv_8_35_n696 = 8'h23 ;
assign n697 =  ( n695 ) == ( bv_8_35_n696 )  ;
assign n698 = state_in[127:120] ;
assign n699 =  ( n698 ) == ( bv_8_34_n117 )  ;
assign n700 = state_in[127:120] ;
assign n701 =  ( n700 ) == ( bv_8_33_n486 )  ;
assign n702 = state_in[127:120] ;
assign n703 =  ( n702 ) == ( bv_8_32_n463 )  ;
assign n704 = state_in[127:120] ;
assign bv_8_31_n705 = 8'h1f ;
assign n706 =  ( n704 ) == ( bv_8_31_n705 )  ;
assign n707 = state_in[127:120] ;
assign n708 =  ( n707 ) == ( bv_8_30_n21 )  ;
assign n709 = state_in[127:120] ;
assign n710 =  ( n709 ) == ( bv_8_29_n625 )  ;
assign n711 = state_in[127:120] ;
assign n712 =  ( n711 ) == ( bv_8_28_n162 )  ;
assign n713 = state_in[127:120] ;
assign n714 =  ( n713 ) == ( bv_8_27_n642 )  ;
assign n715 = state_in[127:120] ;
assign n716 =  ( n715 ) == ( bv_8_26_n53 )  ;
assign n717 = state_in[127:120] ;
assign n718 =  ( n717 ) == ( bv_8_25_n399 )  ;
assign n719 = state_in[127:120] ;
assign n720 =  ( n719 ) == ( bv_8_24_n448 )  ;
assign n721 = state_in[127:120] ;
assign n722 =  ( n721 ) == ( bv_8_23_n144 )  ;
assign n723 = state_in[127:120] ;
assign n724 =  ( n723 ) == ( bv_8_22_n357 )  ;
assign n725 = state_in[127:120] ;
assign n726 =  ( n725 ) == ( bv_8_21_n89 )  ;
assign n727 = state_in[127:120] ;
assign n728 =  ( n727 ) == ( bv_8_20_n341 )  ;
assign n729 = state_in[127:120] ;
assign n730 =  ( n729 ) == ( bv_8_19_n588 )  ;
assign n731 = state_in[127:120] ;
assign n732 =  ( n731 ) == ( bv_8_18_n628 )  ;
assign n733 = state_in[127:120] ;
assign n734 =  ( n733 ) == ( bv_8_17_n525 )  ;
assign n735 = state_in[127:120] ;
assign n736 =  ( n735 ) == ( bv_8_16_n248 )  ;
assign n737 = state_in[127:120] ;
assign n738 =  ( n737 ) == ( bv_8_15_n190 )  ;
assign n739 = state_in[127:120] ;
assign n740 =  ( n739 ) == ( bv_8_14_n648 )  ;
assign n741 = state_in[127:120] ;
assign n742 =  ( n741 ) == ( bv_8_13_n194 )  ;
assign n743 = state_in[127:120] ;
assign n744 =  ( n743 ) == ( bv_8_12_n333 )  ;
assign n745 = state_in[127:120] ;
assign n746 =  ( n745 ) == ( bv_8_11_n379 )  ;
assign n747 = state_in[127:120] ;
assign n748 =  ( n747 ) == ( bv_8_10_n655 )  ;
assign n749 = state_in[127:120] ;
assign n750 =  ( n749 ) == ( bv_8_9_n57 )  ;
assign bv_8_2_n751 = 8'h2 ;
assign n752 = state_in[127:120] ;
assign n753 =  ( n752 ) == ( bv_8_8_n669 )  ;
assign n754 = state_in[127:120] ;
assign n755 =  ( n754 ) == ( bv_8_7_n105 )  ;
assign n756 = state_in[127:120] ;
assign n757 =  ( n756 ) == ( bv_8_6_n169 )  ;
assign n758 = state_in[127:120] ;
assign n759 =  ( n758 ) == ( bv_8_5_n492 )  ;
assign n760 = state_in[127:120] ;
assign n761 =  ( n760 ) == ( bv_8_4_n516 )  ;
assign n762 = state_in[127:120] ;
assign n763 =  ( n762 ) == ( bv_8_3_n65 )  ;
assign n764 = state_in[127:120] ;
assign n765 =  ( n764 ) == ( bv_8_2_n751 )  ;
assign n766 = state_in[127:120] ;
assign n767 =  ( n766 ) == ( bv_8_1_n287 )  ;
assign n768 = state_in[127:120] ;
assign n769 =  ( n768 ) == ( bv_8_0_n580 )  ;
assign n770 =  ( n769 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n771 =  ( n767 ) ? ( bv_8_248_n31 ) : ( n770 ) ;
assign n772 =  ( n765 ) ? ( bv_8_238_n71 ) : ( n771 ) ;
assign n773 =  ( n763 ) ? ( bv_8_246_n39 ) : ( n772 ) ;
assign n774 =  ( n761 ) ? ( bv_8_255_n3 ) : ( n773 ) ;
assign n775 =  ( n759 ) ? ( bv_8_214_n164 ) : ( n774 ) ;
assign n776 =  ( n757 ) ? ( bv_8_222_n134 ) : ( n775 ) ;
assign n777 =  ( n755 ) ? ( bv_8_145_n397 ) : ( n776 ) ;
assign n778 =  ( n753 ) ? ( bv_8_96_n542 ) : ( n777 ) ;
assign n779 =  ( n750 ) ? ( bv_8_2_n751 ) : ( n778 ) ;
assign n780 =  ( n748 ) ? ( bv_8_206_n192 ) : ( n779 ) ;
assign n781 =  ( n746 ) ? ( bv_8_86_n567 ) : ( n780 ) ;
assign n782 =  ( n744 ) ? ( bv_8_231_n99 ) : ( n781 ) ;
assign n783 =  ( n742 ) ? ( bv_8_181_n281 ) : ( n782 ) ;
assign n784 =  ( n740 ) ? ( bv_8_77_n593 ) : ( n783 ) ;
assign n785 =  ( n738 ) ? ( bv_8_236_n79 ) : ( n784 ) ;
assign n786 =  ( n736 ) ? ( bv_8_143_n403 ) : ( n785 ) ;
assign n787 =  ( n734 ) ? ( bv_8_31_n705 ) : ( n786 ) ;
assign n788 =  ( n732 ) ? ( bv_8_137_n421 ) : ( n787 ) ;
assign n789 =  ( n730 ) ? ( bv_8_250_n23 ) : ( n788 ) ;
assign n790 =  ( n728 ) ? ( bv_8_239_n67 ) : ( n789 ) ;
assign n791 =  ( n726 ) ? ( bv_8_178_n292 ) : ( n790 ) ;
assign n792 =  ( n724 ) ? ( bv_8_142_n406 ) : ( n791 ) ;
assign n793 =  ( n722 ) ? ( bv_8_251_n19 ) : ( n792 ) ;
assign n794 =  ( n720 ) ? ( bv_8_65_n623 ) : ( n793 ) ;
assign n795 =  ( n718 ) ? ( bv_8_179_n289 ) : ( n794 ) ;
assign n796 =  ( n716 ) ? ( bv_8_95_n545 ) : ( n795 ) ;
assign n797 =  ( n714 ) ? ( bv_8_69_n612 ) : ( n796 ) ;
assign n798 =  ( n712 ) ? ( bv_8_35_n696 ) : ( n797 ) ;
assign n799 =  ( n710 ) ? ( bv_8_83_n575 ) : ( n798 ) ;
assign n800 =  ( n708 ) ? ( bv_8_228_n111 ) : ( n799 ) ;
assign n801 =  ( n706 ) ? ( bv_8_155_n364 ) : ( n800 ) ;
assign n802 =  ( n703 ) ? ( bv_8_117_n484 ) : ( n801 ) ;
assign n803 =  ( n701 ) ? ( bv_8_225_n123 ) : ( n802 ) ;
assign n804 =  ( n699 ) ? ( bv_8_61_n634 ) : ( n803 ) ;
assign n805 =  ( n697 ) ? ( bv_8_76_n596 ) : ( n804 ) ;
assign n806 =  ( n694 ) ? ( bv_8_108_n510 ) : ( n805 ) ;
assign n807 =  ( n692 ) ? ( bv_8_126_n456 ) : ( n806 ) ;
assign n808 =  ( n690 ) ? ( bv_8_245_n43 ) : ( n807 ) ;
assign n809 =  ( n688 ) ? ( bv_8_131_n440 ) : ( n808 ) ;
assign n810 =  ( n686 ) ? ( bv_8_104_n520 ) : ( n809 ) ;
assign n811 =  ( n684 ) ? ( bv_8_81_n582 ) : ( n810 ) ;
assign n812 =  ( n682 ) ? ( bv_8_209_n182 ) : ( n811 ) ;
assign n813 =  ( n680 ) ? ( bv_8_249_n27 ) : ( n812 ) ;
assign n814 =  ( n678 ) ? ( bv_8_226_n119 ) : ( n813 ) ;
assign n815 =  ( n676 ) ? ( bv_8_171_n314 ) : ( n814 ) ;
assign n816 =  ( n674 ) ? ( bv_8_98_n536 ) : ( n815 ) ;
assign n817 =  ( n671 ) ? ( bv_8_42_n672 ) : ( n816 ) ;
assign n818 =  ( n668 ) ? ( bv_8_8_n669 ) : ( n817 ) ;
assign n819 =  ( n666 ) ? ( bv_8_149_n384 ) : ( n818 ) ;
assign n820 =  ( n664 ) ? ( bv_8_70_n609 ) : ( n819 ) ;
assign n821 =  ( n662 ) ? ( bv_8_157_n359 ) : ( n820 ) ;
assign n822 =  ( n659 ) ? ( bv_8_48_n660 ) : ( n821 ) ;
assign n823 =  ( n657 ) ? ( bv_8_55_n650 ) : ( n822 ) ;
assign n824 =  ( n654 ) ? ( bv_8_10_n655 ) : ( n823 ) ;
assign n825 =  ( n651 ) ? ( bv_8_47_n652 ) : ( n824 ) ;
assign n826 =  ( n647 ) ? ( bv_8_14_n648 ) : ( n825 ) ;
assign n827 =  ( n644 ) ? ( bv_8_36_n645 ) : ( n826 ) ;
assign n828 =  ( n641 ) ? ( bv_8_27_n642 ) : ( n827 ) ;
assign n829 =  ( n639 ) ? ( bv_8_223_n130 ) : ( n828 ) ;
assign n830 =  ( n637 ) ? ( bv_8_205_n196 ) : ( n829 ) ;
assign n831 =  ( n635 ) ? ( bv_8_78_n590 ) : ( n830 ) ;
assign n832 =  ( n632 ) ? ( bv_8_127_n453 ) : ( n831 ) ;
assign n833 =  ( n630 ) ? ( bv_8_234_n87 ) : ( n832 ) ;
assign n834 =  ( n627 ) ? ( bv_8_18_n628 ) : ( n833 ) ;
assign n835 =  ( n624 ) ? ( bv_8_29_n625 ) : ( n834 ) ;
assign n836 =  ( n621 ) ? ( bv_8_88_n562 ) : ( n835 ) ;
assign n837 =  ( n618 ) ? ( bv_8_52_n619 ) : ( n836 ) ;
assign n838 =  ( n615 ) ? ( bv_8_54_n616 ) : ( n837 ) ;
assign n839 =  ( n613 ) ? ( bv_8_220_n142 ) : ( n838 ) ;
assign n840 =  ( n610 ) ? ( bv_8_180_n285 ) : ( n839 ) ;
assign n841 =  ( n607 ) ? ( bv_8_91_n555 ) : ( n840 ) ;
assign n842 =  ( n605 ) ? ( bv_8_164_n335 ) : ( n841 ) ;
assign n843 =  ( n603 ) ? ( bv_8_118_n480 ) : ( n842 ) ;
assign n844 =  ( n601 ) ? ( bv_8_183_n273 ) : ( n843 ) ;
assign n845 =  ( n599 ) ? ( bv_8_125_n459 ) : ( n844 ) ;
assign n846 =  ( n597 ) ? ( bv_8_82_n578 ) : ( n845 ) ;
assign n847 =  ( n594 ) ? ( bv_8_221_n138 ) : ( n846 ) ;
assign n848 =  ( n591 ) ? ( bv_8_94_n548 ) : ( n847 ) ;
assign n849 =  ( n587 ) ? ( bv_8_19_n588 ) : ( n848 ) ;
assign n850 =  ( n585 ) ? ( bv_8_166_n328 ) : ( n849 ) ;
assign n851 =  ( n583 ) ? ( bv_8_185_n266 ) : ( n850 ) ;
assign n852 =  ( n579 ) ? ( bv_8_0_n580 ) : ( n851 ) ;
assign n853 =  ( n576 ) ? ( bv_8_193_n239 ) : ( n852 ) ;
assign n854 =  ( n572 ) ? ( bv_8_64_n573 ) : ( n853 ) ;
assign n855 =  ( n570 ) ? ( bv_8_227_n115 ) : ( n854 ) ;
assign n856 =  ( n568 ) ? ( bv_8_121_n470 ) : ( n855 ) ;
assign n857 =  ( n565 ) ? ( bv_8_182_n277 ) : ( n856 ) ;
assign n858 =  ( n563 ) ? ( bv_8_212_n171 ) : ( n857 ) ;
assign n859 =  ( n560 ) ? ( bv_8_141_n410 ) : ( n858 ) ;
assign n860 =  ( n558 ) ? ( bv_8_103_n523 ) : ( n859 ) ;
assign n861 =  ( n556 ) ? ( bv_8_114_n494 ) : ( n860 ) ;
assign n862 =  ( n553 ) ? ( bv_8_148_n388 ) : ( n861 ) ;
assign n863 =  ( n551 ) ? ( bv_8_152_n374 ) : ( n862 ) ;
assign n864 =  ( n549 ) ? ( bv_8_176_n299 ) : ( n863 ) ;
assign n865 =  ( n546 ) ? ( bv_8_133_n434 ) : ( n864 ) ;
assign n866 =  ( n543 ) ? ( bv_8_187_n260 ) : ( n865 ) ;
assign n867 =  ( n540 ) ? ( bv_8_197_n224 ) : ( n866 ) ;
assign n868 =  ( n537 ) ? ( bv_8_79_n538 ) : ( n867 ) ;
assign n869 =  ( n534 ) ? ( bv_8_237_n75 ) : ( n868 ) ;
assign n870 =  ( n532 ) ? ( bv_8_134_n431 ) : ( n869 ) ;
assign n871 =  ( n530 ) ? ( bv_8_154_n368 ) : ( n870 ) ;
assign n872 =  ( n528 ) ? ( bv_8_102_n527 ) : ( n871 ) ;
assign n873 =  ( n524 ) ? ( bv_8_17_n525 ) : ( n872 ) ;
assign n874 =  ( n521 ) ? ( bv_8_138_n418 ) : ( n873 ) ;
assign n875 =  ( n518 ) ? ( bv_8_233_n91 ) : ( n874 ) ;
assign n876 =  ( n515 ) ? ( bv_8_4_n516 ) : ( n875 ) ;
assign n877 =  ( n513 ) ? ( bv_8_254_n7 ) : ( n876 ) ;
assign n878 =  ( n511 ) ? ( bv_8_160_n350 ) : ( n877 ) ;
assign n879 =  ( n508 ) ? ( bv_8_120_n474 ) : ( n878 ) ;
assign n880 =  ( n505 ) ? ( bv_8_37_n506 ) : ( n879 ) ;
assign n881 =  ( n502 ) ? ( bv_8_75_n503 ) : ( n880 ) ;
assign n882 =  ( n500 ) ? ( bv_8_162_n343 ) : ( n881 ) ;
assign n883 =  ( n497 ) ? ( bv_8_93_n498 ) : ( n882 ) ;
assign n884 =  ( n495 ) ? ( bv_8_128_n450 ) : ( n883 ) ;
assign n885 =  ( n491 ) ? ( bv_8_5_n492 ) : ( n884 ) ;
assign n886 =  ( n488 ) ? ( bv_8_63_n489 ) : ( n885 ) ;
assign n887 =  ( n485 ) ? ( bv_8_33_n486 ) : ( n886 ) ;
assign n888 =  ( n481 ) ? ( bv_8_112_n482 ) : ( n887 ) ;
assign n889 =  ( n478 ) ? ( bv_8_241_n59 ) : ( n888 ) ;
assign n890 =  ( n475 ) ? ( bv_8_99_n476 ) : ( n889 ) ;
assign n891 =  ( n471 ) ? ( bv_8_119_n472 ) : ( n890 ) ;
assign n892 =  ( n468 ) ? ( bv_8_175_n302 ) : ( n891 ) ;
assign n893 =  ( n465 ) ? ( bv_8_66_n466 ) : ( n892 ) ;
assign n894 =  ( n462 ) ? ( bv_8_32_n463 ) : ( n893 ) ;
assign n895 =  ( n460 ) ? ( bv_8_229_n107 ) : ( n894 ) ;
assign n896 =  ( n457 ) ? ( bv_8_253_n11 ) : ( n895 ) ;
assign n897 =  ( n454 ) ? ( bv_8_191_n246 ) : ( n896 ) ;
assign n898 =  ( n451 ) ? ( bv_8_129_n446 ) : ( n897 ) ;
assign n899 =  ( n447 ) ? ( bv_8_24_n448 ) : ( n898 ) ;
assign n900 =  ( n443 ) ? ( bv_8_38_n444 ) : ( n899 ) ;
assign n901 =  ( n441 ) ? ( bv_8_195_n232 ) : ( n900 ) ;
assign n902 =  ( n438 ) ? ( bv_8_190_n250 ) : ( n901 ) ;
assign n903 =  ( n435 ) ? ( bv_8_53_n436 ) : ( n902 ) ;
assign n904 =  ( n432 ) ? ( bv_8_136_n425 ) : ( n903 ) ;
assign n905 =  ( n428 ) ? ( bv_8_46_n429 ) : ( n904 ) ;
assign n906 =  ( n426 ) ? ( bv_8_147_n392 ) : ( n905 ) ;
assign n907 =  ( n422 ) ? ( bv_8_85_n423 ) : ( n906 ) ;
assign n908 =  ( n419 ) ? ( bv_8_252_n15 ) : ( n907 ) ;
assign n909 =  ( n415 ) ? ( bv_8_122_n416 ) : ( n908 ) ;
assign n910 =  ( n413 ) ? ( bv_8_200_n213 ) : ( n909 ) ;
assign n911 =  ( n411 ) ? ( bv_8_186_n263 ) : ( n910 ) ;
assign n912 =  ( n407 ) ? ( bv_8_50_n408 ) : ( n911 ) ;
assign n913 =  ( n404 ) ? ( bv_8_230_n103 ) : ( n912 ) ;
assign n914 =  ( n401 ) ? ( bv_8_192_n242 ) : ( n913 ) ;
assign n915 =  ( n398 ) ? ( bv_8_25_n399 ) : ( n914 ) ;
assign n916 =  ( n395 ) ? ( bv_8_158_n355 ) : ( n915 ) ;
assign n917 =  ( n393 ) ? ( bv_8_163_n339 ) : ( n916 ) ;
assign n918 =  ( n389 ) ? ( bv_8_68_n390 ) : ( n917 ) ;
assign n919 =  ( n385 ) ? ( bv_8_84_n386 ) : ( n918 ) ;
assign n920 =  ( n381 ) ? ( bv_8_59_n382 ) : ( n919 ) ;
assign n921 =  ( n378 ) ? ( bv_8_11_n379 ) : ( n920 ) ;
assign n922 =  ( n375 ) ? ( bv_8_140_n376 ) : ( n921 ) ;
assign n923 =  ( n372 ) ? ( bv_8_199_n216 ) : ( n922 ) ;
assign n924 =  ( n369 ) ? ( bv_8_107_n370 ) : ( n923 ) ;
assign n925 =  ( n365 ) ? ( bv_8_40_n366 ) : ( n924 ) ;
assign n926 =  ( n362 ) ? ( bv_8_167_n325 ) : ( n925 ) ;
assign n927 =  ( n360 ) ? ( bv_8_188_n257 ) : ( n926 ) ;
assign n928 =  ( n356 ) ? ( bv_8_22_n357 ) : ( n927 ) ;
assign n929 =  ( n353 ) ? ( bv_8_173_n307 ) : ( n928 ) ;
assign n930 =  ( n351 ) ? ( bv_8_219_n146 ) : ( n929 ) ;
assign n931 =  ( n347 ) ? ( bv_8_100_n348 ) : ( n930 ) ;
assign n932 =  ( n344 ) ? ( bv_8_116_n345 ) : ( n931 ) ;
assign n933 =  ( n340 ) ? ( bv_8_20_n341 ) : ( n932 ) ;
assign n934 =  ( n336 ) ? ( bv_8_146_n337 ) : ( n933 ) ;
assign n935 =  ( n332 ) ? ( bv_8_12_n333 ) : ( n934 ) ;
assign n936 =  ( n329 ) ? ( bv_8_72_n330 ) : ( n935 ) ;
assign n937 =  ( n326 ) ? ( bv_8_184_n270 ) : ( n936 ) ;
assign n938 =  ( n322 ) ? ( bv_8_159_n323 ) : ( n937 ) ;
assign n939 =  ( n320 ) ? ( bv_8_189_n254 ) : ( n938 ) ;
assign n940 =  ( n317 ) ? ( bv_8_67_n318 ) : ( n939 ) ;
assign n941 =  ( n315 ) ? ( bv_8_196_n228 ) : ( n940 ) ;
assign n942 =  ( n311 ) ? ( bv_8_57_n312 ) : ( n941 ) ;
assign n943 =  ( n308 ) ? ( bv_8_49_n309 ) : ( n942 ) ;
assign n944 =  ( n305 ) ? ( bv_8_211_n175 ) : ( n943 ) ;
assign n945 =  ( n303 ) ? ( bv_8_242_n55 ) : ( n944 ) ;
assign n946 =  ( n300 ) ? ( bv_8_213_n167 ) : ( n945 ) ;
assign n947 =  ( n296 ) ? ( bv_8_139_n297 ) : ( n946 ) ;
assign n948 =  ( n293 ) ? ( bv_8_110_n294 ) : ( n947 ) ;
assign n949 =  ( n290 ) ? ( bv_8_218_n150 ) : ( n948 ) ;
assign n950 =  ( n286 ) ? ( bv_8_1_n287 ) : ( n949 ) ;
assign n951 =  ( n282 ) ? ( bv_8_177_n283 ) : ( n950 ) ;
assign n952 =  ( n278 ) ? ( bv_8_156_n279 ) : ( n951 ) ;
assign n953 =  ( n274 ) ? ( bv_8_73_n275 ) : ( n952 ) ;
assign n954 =  ( n271 ) ? ( bv_8_216_n157 ) : ( n953 ) ;
assign n955 =  ( n267 ) ? ( bv_8_172_n268 ) : ( n954 ) ;
assign n956 =  ( n264 ) ? ( bv_8_243_n51 ) : ( n955 ) ;
assign n957 =  ( n261 ) ? ( bv_8_207_n188 ) : ( n956 ) ;
assign n958 =  ( n258 ) ? ( bv_8_202_n207 ) : ( n957 ) ;
assign n959 =  ( n255 ) ? ( bv_8_244_n47 ) : ( n958 ) ;
assign n960 =  ( n251 ) ? ( bv_8_71_n252 ) : ( n959 ) ;
assign n961 =  ( n247 ) ? ( bv_8_16_n248 ) : ( n960 ) ;
assign n962 =  ( n243 ) ? ( bv_8_111_n244 ) : ( n961 ) ;
assign n963 =  ( n240 ) ? ( bv_8_240_n63 ) : ( n962 ) ;
assign n964 =  ( n236 ) ? ( bv_8_74_n237 ) : ( n963 ) ;
assign n965 =  ( n233 ) ? ( bv_8_92_n234 ) : ( n964 ) ;
assign n966 =  ( n229 ) ? ( bv_8_56_n230 ) : ( n965 ) ;
assign n967 =  ( n225 ) ? ( bv_8_87_n226 ) : ( n966 ) ;
assign n968 =  ( n221 ) ? ( bv_8_115_n222 ) : ( n967 ) ;
assign n969 =  ( n217 ) ? ( bv_8_151_n218 ) : ( n968 ) ;
assign n970 =  ( n214 ) ? ( bv_8_203_n203 ) : ( n969 ) ;
assign n971 =  ( n210 ) ? ( bv_8_161_n211 ) : ( n970 ) ;
assign n972 =  ( n208 ) ? ( bv_8_232_n95 ) : ( n971 ) ;
assign n973 =  ( n204 ) ? ( bv_8_62_n205 ) : ( n972 ) ;
assign n974 =  ( n200 ) ? ( bv_8_150_n201 ) : ( n973 ) ;
assign n975 =  ( n197 ) ? ( bv_8_97_n198 ) : ( n974 ) ;
assign n976 =  ( n193 ) ? ( bv_8_13_n194 ) : ( n975 ) ;
assign n977 =  ( n189 ) ? ( bv_8_15_n190 ) : ( n976 ) ;
assign n978 =  ( n186 ) ? ( bv_8_224_n126 ) : ( n977 ) ;
assign n979 =  ( n183 ) ? ( bv_8_124_n184 ) : ( n978 ) ;
assign n980 =  ( n179 ) ? ( bv_8_113_n180 ) : ( n979 ) ;
assign n981 =  ( n176 ) ? ( bv_8_204_n177 ) : ( n980 ) ;
assign n982 =  ( n172 ) ? ( bv_8_144_n173 ) : ( n981 ) ;
assign n983 =  ( n168 ) ? ( bv_8_6_n169 ) : ( n982 ) ;
assign n984 =  ( n165 ) ? ( bv_8_247_n35 ) : ( n983 ) ;
assign n985 =  ( n161 ) ? ( bv_8_28_n162 ) : ( n984 ) ;
assign n986 =  ( n158 ) ? ( bv_8_194_n159 ) : ( n985 ) ;
assign n987 =  ( n154 ) ? ( bv_8_106_n155 ) : ( n986 ) ;
assign n988 =  ( n151 ) ? ( bv_8_174_n152 ) : ( n987 ) ;
assign n989 =  ( n147 ) ? ( bv_8_105_n148 ) : ( n988 ) ;
assign n990 =  ( n143 ) ? ( bv_8_23_n144 ) : ( n989 ) ;
assign n991 =  ( n139 ) ? ( bv_8_153_n140 ) : ( n990 ) ;
assign n992 =  ( n135 ) ? ( bv_8_58_n136 ) : ( n991 ) ;
assign n993 =  ( n131 ) ? ( bv_8_39_n132 ) : ( n992 ) ;
assign n994 =  ( n127 ) ? ( bv_8_217_n128 ) : ( n993 ) ;
assign n995 =  ( n124 ) ? ( bv_8_235_n83 ) : ( n994 ) ;
assign n996 =  ( n120 ) ? ( bv_8_43_n121 ) : ( n995 ) ;
assign n997 =  ( n116 ) ? ( bv_8_34_n117 ) : ( n996 ) ;
assign n998 =  ( n112 ) ? ( bv_8_210_n113 ) : ( n997 ) ;
assign n999 =  ( n108 ) ? ( bv_8_169_n109 ) : ( n998 ) ;
assign n1000 =  ( n104 ) ? ( bv_8_7_n105 ) : ( n999 ) ;
assign n1001 =  ( n100 ) ? ( bv_8_51_n101 ) : ( n1000 ) ;
assign n1002 =  ( n96 ) ? ( bv_8_45_n97 ) : ( n1001 ) ;
assign n1003 =  ( n92 ) ? ( bv_8_60_n93 ) : ( n1002 ) ;
assign n1004 =  ( n88 ) ? ( bv_8_21_n89 ) : ( n1003 ) ;
assign n1005 =  ( n84 ) ? ( bv_8_201_n85 ) : ( n1004 ) ;
assign n1006 =  ( n80 ) ? ( bv_8_135_n81 ) : ( n1005 ) ;
assign n1007 =  ( n76 ) ? ( bv_8_170_n77 ) : ( n1006 ) ;
assign n1008 =  ( n72 ) ? ( bv_8_80_n73 ) : ( n1007 ) ;
assign n1009 =  ( n68 ) ? ( bv_8_165_n69 ) : ( n1008 ) ;
assign n1010 =  ( n64 ) ? ( bv_8_3_n65 ) : ( n1009 ) ;
assign n1011 =  ( n60 ) ? ( bv_8_89_n61 ) : ( n1010 ) ;
assign n1012 =  ( n56 ) ? ( bv_8_9_n57 ) : ( n1011 ) ;
assign n1013 =  ( n52 ) ? ( bv_8_26_n53 ) : ( n1012 ) ;
assign n1014 =  ( n48 ) ? ( bv_8_101_n49 ) : ( n1013 ) ;
assign n1015 =  ( n44 ) ? ( bv_8_215_n45 ) : ( n1014 ) ;
assign n1016 =  ( n40 ) ? ( bv_8_132_n41 ) : ( n1015 ) ;
assign n1017 =  ( n36 ) ? ( bv_8_208_n37 ) : ( n1016 ) ;
assign n1018 =  ( n32 ) ? ( bv_8_130_n33 ) : ( n1017 ) ;
assign n1019 =  ( n28 ) ? ( bv_8_41_n29 ) : ( n1018 ) ;
assign n1020 =  ( n24 ) ? ( bv_8_90_n25 ) : ( n1019 ) ;
assign n1021 =  ( n20 ) ? ( bv_8_30_n21 ) : ( n1020 ) ;
assign n1022 =  ( n16 ) ? ( bv_8_123_n17 ) : ( n1021 ) ;
assign n1023 =  ( n12 ) ? ( bv_8_168_n13 ) : ( n1022 ) ;
assign n1024 =  ( n8 ) ? ( bv_8_109_n9 ) : ( n1023 ) ;
assign n1025 =  ( n4 ) ? ( bv_8_44_n5 ) : ( n1024 ) ;
assign n1026 = state_in[87:80] ;
assign n1027 =  ( n1026 ) == ( bv_8_255_n3 )  ;
assign n1028 = state_in[87:80] ;
assign n1029 =  ( n1028 ) == ( bv_8_254_n7 )  ;
assign n1030 = state_in[87:80] ;
assign n1031 =  ( n1030 ) == ( bv_8_253_n11 )  ;
assign n1032 = state_in[87:80] ;
assign n1033 =  ( n1032 ) == ( bv_8_252_n15 )  ;
assign n1034 = state_in[87:80] ;
assign n1035 =  ( n1034 ) == ( bv_8_251_n19 )  ;
assign n1036 = state_in[87:80] ;
assign n1037 =  ( n1036 ) == ( bv_8_250_n23 )  ;
assign n1038 = state_in[87:80] ;
assign n1039 =  ( n1038 ) == ( bv_8_249_n27 )  ;
assign n1040 = state_in[87:80] ;
assign n1041 =  ( n1040 ) == ( bv_8_248_n31 )  ;
assign n1042 = state_in[87:80] ;
assign n1043 =  ( n1042 ) == ( bv_8_247_n35 )  ;
assign n1044 = state_in[87:80] ;
assign n1045 =  ( n1044 ) == ( bv_8_246_n39 )  ;
assign n1046 = state_in[87:80] ;
assign n1047 =  ( n1046 ) == ( bv_8_245_n43 )  ;
assign n1048 = state_in[87:80] ;
assign n1049 =  ( n1048 ) == ( bv_8_244_n47 )  ;
assign n1050 = state_in[87:80] ;
assign n1051 =  ( n1050 ) == ( bv_8_243_n51 )  ;
assign n1052 = state_in[87:80] ;
assign n1053 =  ( n1052 ) == ( bv_8_242_n55 )  ;
assign n1054 = state_in[87:80] ;
assign n1055 =  ( n1054 ) == ( bv_8_241_n59 )  ;
assign n1056 = state_in[87:80] ;
assign n1057 =  ( n1056 ) == ( bv_8_240_n63 )  ;
assign n1058 = state_in[87:80] ;
assign n1059 =  ( n1058 ) == ( bv_8_239_n67 )  ;
assign n1060 = state_in[87:80] ;
assign n1061 =  ( n1060 ) == ( bv_8_238_n71 )  ;
assign n1062 = state_in[87:80] ;
assign n1063 =  ( n1062 ) == ( bv_8_237_n75 )  ;
assign n1064 = state_in[87:80] ;
assign n1065 =  ( n1064 ) == ( bv_8_236_n79 )  ;
assign n1066 = state_in[87:80] ;
assign n1067 =  ( n1066 ) == ( bv_8_235_n83 )  ;
assign n1068 = state_in[87:80] ;
assign n1069 =  ( n1068 ) == ( bv_8_234_n87 )  ;
assign n1070 = state_in[87:80] ;
assign n1071 =  ( n1070 ) == ( bv_8_233_n91 )  ;
assign n1072 = state_in[87:80] ;
assign n1073 =  ( n1072 ) == ( bv_8_232_n95 )  ;
assign n1074 = state_in[87:80] ;
assign n1075 =  ( n1074 ) == ( bv_8_231_n99 )  ;
assign n1076 = state_in[87:80] ;
assign n1077 =  ( n1076 ) == ( bv_8_230_n103 )  ;
assign n1078 = state_in[87:80] ;
assign n1079 =  ( n1078 ) == ( bv_8_229_n107 )  ;
assign n1080 = state_in[87:80] ;
assign n1081 =  ( n1080 ) == ( bv_8_228_n111 )  ;
assign n1082 = state_in[87:80] ;
assign n1083 =  ( n1082 ) == ( bv_8_227_n115 )  ;
assign n1084 = state_in[87:80] ;
assign n1085 =  ( n1084 ) == ( bv_8_226_n119 )  ;
assign n1086 = state_in[87:80] ;
assign n1087 =  ( n1086 ) == ( bv_8_225_n123 )  ;
assign n1088 = state_in[87:80] ;
assign n1089 =  ( n1088 ) == ( bv_8_224_n126 )  ;
assign n1090 = state_in[87:80] ;
assign n1091 =  ( n1090 ) == ( bv_8_223_n130 )  ;
assign n1092 = state_in[87:80] ;
assign n1093 =  ( n1092 ) == ( bv_8_222_n134 )  ;
assign n1094 = state_in[87:80] ;
assign n1095 =  ( n1094 ) == ( bv_8_221_n138 )  ;
assign n1096 = state_in[87:80] ;
assign n1097 =  ( n1096 ) == ( bv_8_220_n142 )  ;
assign n1098 = state_in[87:80] ;
assign n1099 =  ( n1098 ) == ( bv_8_219_n146 )  ;
assign n1100 = state_in[87:80] ;
assign n1101 =  ( n1100 ) == ( bv_8_218_n150 )  ;
assign n1102 = state_in[87:80] ;
assign n1103 =  ( n1102 ) == ( bv_8_217_n128 )  ;
assign n1104 = state_in[87:80] ;
assign n1105 =  ( n1104 ) == ( bv_8_216_n157 )  ;
assign n1106 = state_in[87:80] ;
assign n1107 =  ( n1106 ) == ( bv_8_215_n45 )  ;
assign n1108 = state_in[87:80] ;
assign n1109 =  ( n1108 ) == ( bv_8_214_n164 )  ;
assign n1110 = state_in[87:80] ;
assign n1111 =  ( n1110 ) == ( bv_8_213_n167 )  ;
assign n1112 = state_in[87:80] ;
assign n1113 =  ( n1112 ) == ( bv_8_212_n171 )  ;
assign n1114 = state_in[87:80] ;
assign n1115 =  ( n1114 ) == ( bv_8_211_n175 )  ;
assign n1116 = state_in[87:80] ;
assign n1117 =  ( n1116 ) == ( bv_8_210_n113 )  ;
assign n1118 = state_in[87:80] ;
assign n1119 =  ( n1118 ) == ( bv_8_209_n182 )  ;
assign n1120 = state_in[87:80] ;
assign n1121 =  ( n1120 ) == ( bv_8_208_n37 )  ;
assign n1122 = state_in[87:80] ;
assign n1123 =  ( n1122 ) == ( bv_8_207_n188 )  ;
assign n1124 = state_in[87:80] ;
assign n1125 =  ( n1124 ) == ( bv_8_206_n192 )  ;
assign n1126 = state_in[87:80] ;
assign n1127 =  ( n1126 ) == ( bv_8_205_n196 )  ;
assign n1128 = state_in[87:80] ;
assign n1129 =  ( n1128 ) == ( bv_8_204_n177 )  ;
assign n1130 = state_in[87:80] ;
assign n1131 =  ( n1130 ) == ( bv_8_203_n203 )  ;
assign n1132 = state_in[87:80] ;
assign n1133 =  ( n1132 ) == ( bv_8_202_n207 )  ;
assign n1134 = state_in[87:80] ;
assign n1135 =  ( n1134 ) == ( bv_8_201_n85 )  ;
assign n1136 = state_in[87:80] ;
assign n1137 =  ( n1136 ) == ( bv_8_200_n213 )  ;
assign n1138 = state_in[87:80] ;
assign n1139 =  ( n1138 ) == ( bv_8_199_n216 )  ;
assign n1140 = state_in[87:80] ;
assign n1141 =  ( n1140 ) == ( bv_8_198_n220 )  ;
assign n1142 = state_in[87:80] ;
assign n1143 =  ( n1142 ) == ( bv_8_197_n224 )  ;
assign n1144 = state_in[87:80] ;
assign n1145 =  ( n1144 ) == ( bv_8_196_n228 )  ;
assign n1146 = state_in[87:80] ;
assign n1147 =  ( n1146 ) == ( bv_8_195_n232 )  ;
assign n1148 = state_in[87:80] ;
assign n1149 =  ( n1148 ) == ( bv_8_194_n159 )  ;
assign n1150 = state_in[87:80] ;
assign n1151 =  ( n1150 ) == ( bv_8_193_n239 )  ;
assign n1152 = state_in[87:80] ;
assign n1153 =  ( n1152 ) == ( bv_8_192_n242 )  ;
assign n1154 = state_in[87:80] ;
assign n1155 =  ( n1154 ) == ( bv_8_191_n246 )  ;
assign n1156 = state_in[87:80] ;
assign n1157 =  ( n1156 ) == ( bv_8_190_n250 )  ;
assign n1158 = state_in[87:80] ;
assign n1159 =  ( n1158 ) == ( bv_8_189_n254 )  ;
assign n1160 = state_in[87:80] ;
assign n1161 =  ( n1160 ) == ( bv_8_188_n257 )  ;
assign n1162 = state_in[87:80] ;
assign n1163 =  ( n1162 ) == ( bv_8_187_n260 )  ;
assign n1164 = state_in[87:80] ;
assign n1165 =  ( n1164 ) == ( bv_8_186_n263 )  ;
assign n1166 = state_in[87:80] ;
assign n1167 =  ( n1166 ) == ( bv_8_185_n266 )  ;
assign n1168 = state_in[87:80] ;
assign n1169 =  ( n1168 ) == ( bv_8_184_n270 )  ;
assign n1170 = state_in[87:80] ;
assign n1171 =  ( n1170 ) == ( bv_8_183_n273 )  ;
assign n1172 = state_in[87:80] ;
assign n1173 =  ( n1172 ) == ( bv_8_182_n277 )  ;
assign n1174 = state_in[87:80] ;
assign n1175 =  ( n1174 ) == ( bv_8_181_n281 )  ;
assign n1176 = state_in[87:80] ;
assign n1177 =  ( n1176 ) == ( bv_8_180_n285 )  ;
assign n1178 = state_in[87:80] ;
assign n1179 =  ( n1178 ) == ( bv_8_179_n289 )  ;
assign n1180 = state_in[87:80] ;
assign n1181 =  ( n1180 ) == ( bv_8_178_n292 )  ;
assign n1182 = state_in[87:80] ;
assign n1183 =  ( n1182 ) == ( bv_8_177_n283 )  ;
assign n1184 = state_in[87:80] ;
assign n1185 =  ( n1184 ) == ( bv_8_176_n299 )  ;
assign n1186 = state_in[87:80] ;
assign n1187 =  ( n1186 ) == ( bv_8_175_n302 )  ;
assign n1188 = state_in[87:80] ;
assign n1189 =  ( n1188 ) == ( bv_8_174_n152 )  ;
assign n1190 = state_in[87:80] ;
assign n1191 =  ( n1190 ) == ( bv_8_173_n307 )  ;
assign n1192 = state_in[87:80] ;
assign n1193 =  ( n1192 ) == ( bv_8_172_n268 )  ;
assign n1194 = state_in[87:80] ;
assign n1195 =  ( n1194 ) == ( bv_8_171_n314 )  ;
assign n1196 = state_in[87:80] ;
assign n1197 =  ( n1196 ) == ( bv_8_170_n77 )  ;
assign n1198 = state_in[87:80] ;
assign n1199 =  ( n1198 ) == ( bv_8_169_n109 )  ;
assign n1200 = state_in[87:80] ;
assign n1201 =  ( n1200 ) == ( bv_8_168_n13 )  ;
assign n1202 = state_in[87:80] ;
assign n1203 =  ( n1202 ) == ( bv_8_167_n325 )  ;
assign n1204 = state_in[87:80] ;
assign n1205 =  ( n1204 ) == ( bv_8_166_n328 )  ;
assign n1206 = state_in[87:80] ;
assign n1207 =  ( n1206 ) == ( bv_8_165_n69 )  ;
assign n1208 = state_in[87:80] ;
assign n1209 =  ( n1208 ) == ( bv_8_164_n335 )  ;
assign n1210 = state_in[87:80] ;
assign n1211 =  ( n1210 ) == ( bv_8_163_n339 )  ;
assign n1212 = state_in[87:80] ;
assign n1213 =  ( n1212 ) == ( bv_8_162_n343 )  ;
assign n1214 = state_in[87:80] ;
assign n1215 =  ( n1214 ) == ( bv_8_161_n211 )  ;
assign n1216 = state_in[87:80] ;
assign n1217 =  ( n1216 ) == ( bv_8_160_n350 )  ;
assign n1218 = state_in[87:80] ;
assign n1219 =  ( n1218 ) == ( bv_8_159_n323 )  ;
assign n1220 = state_in[87:80] ;
assign n1221 =  ( n1220 ) == ( bv_8_158_n355 )  ;
assign n1222 = state_in[87:80] ;
assign n1223 =  ( n1222 ) == ( bv_8_157_n359 )  ;
assign n1224 = state_in[87:80] ;
assign n1225 =  ( n1224 ) == ( bv_8_156_n279 )  ;
assign n1226 = state_in[87:80] ;
assign n1227 =  ( n1226 ) == ( bv_8_155_n364 )  ;
assign n1228 = state_in[87:80] ;
assign n1229 =  ( n1228 ) == ( bv_8_154_n368 )  ;
assign n1230 = state_in[87:80] ;
assign n1231 =  ( n1230 ) == ( bv_8_153_n140 )  ;
assign n1232 = state_in[87:80] ;
assign n1233 =  ( n1232 ) == ( bv_8_152_n374 )  ;
assign n1234 = state_in[87:80] ;
assign n1235 =  ( n1234 ) == ( bv_8_151_n218 )  ;
assign n1236 = state_in[87:80] ;
assign n1237 =  ( n1236 ) == ( bv_8_150_n201 )  ;
assign n1238 = state_in[87:80] ;
assign n1239 =  ( n1238 ) == ( bv_8_149_n384 )  ;
assign n1240 = state_in[87:80] ;
assign n1241 =  ( n1240 ) == ( bv_8_148_n388 )  ;
assign n1242 = state_in[87:80] ;
assign n1243 =  ( n1242 ) == ( bv_8_147_n392 )  ;
assign n1244 = state_in[87:80] ;
assign n1245 =  ( n1244 ) == ( bv_8_146_n337 )  ;
assign n1246 = state_in[87:80] ;
assign n1247 =  ( n1246 ) == ( bv_8_145_n397 )  ;
assign n1248 = state_in[87:80] ;
assign n1249 =  ( n1248 ) == ( bv_8_144_n173 )  ;
assign n1250 = state_in[87:80] ;
assign n1251 =  ( n1250 ) == ( bv_8_143_n403 )  ;
assign n1252 = state_in[87:80] ;
assign n1253 =  ( n1252 ) == ( bv_8_142_n406 )  ;
assign n1254 = state_in[87:80] ;
assign n1255 =  ( n1254 ) == ( bv_8_141_n410 )  ;
assign n1256 = state_in[87:80] ;
assign n1257 =  ( n1256 ) == ( bv_8_140_n376 )  ;
assign n1258 = state_in[87:80] ;
assign n1259 =  ( n1258 ) == ( bv_8_139_n297 )  ;
assign n1260 = state_in[87:80] ;
assign n1261 =  ( n1260 ) == ( bv_8_138_n418 )  ;
assign n1262 = state_in[87:80] ;
assign n1263 =  ( n1262 ) == ( bv_8_137_n421 )  ;
assign n1264 = state_in[87:80] ;
assign n1265 =  ( n1264 ) == ( bv_8_136_n425 )  ;
assign n1266 = state_in[87:80] ;
assign n1267 =  ( n1266 ) == ( bv_8_135_n81 )  ;
assign n1268 = state_in[87:80] ;
assign n1269 =  ( n1268 ) == ( bv_8_134_n431 )  ;
assign n1270 = state_in[87:80] ;
assign n1271 =  ( n1270 ) == ( bv_8_133_n434 )  ;
assign n1272 = state_in[87:80] ;
assign n1273 =  ( n1272 ) == ( bv_8_132_n41 )  ;
assign n1274 = state_in[87:80] ;
assign n1275 =  ( n1274 ) == ( bv_8_131_n440 )  ;
assign n1276 = state_in[87:80] ;
assign n1277 =  ( n1276 ) == ( bv_8_130_n33 )  ;
assign n1278 = state_in[87:80] ;
assign n1279 =  ( n1278 ) == ( bv_8_129_n446 )  ;
assign n1280 = state_in[87:80] ;
assign n1281 =  ( n1280 ) == ( bv_8_128_n450 )  ;
assign n1282 = state_in[87:80] ;
assign n1283 =  ( n1282 ) == ( bv_8_127_n453 )  ;
assign n1284 = state_in[87:80] ;
assign n1285 =  ( n1284 ) == ( bv_8_126_n456 )  ;
assign n1286 = state_in[87:80] ;
assign n1287 =  ( n1286 ) == ( bv_8_125_n459 )  ;
assign n1288 = state_in[87:80] ;
assign n1289 =  ( n1288 ) == ( bv_8_124_n184 )  ;
assign n1290 = state_in[87:80] ;
assign n1291 =  ( n1290 ) == ( bv_8_123_n17 )  ;
assign n1292 = state_in[87:80] ;
assign n1293 =  ( n1292 ) == ( bv_8_122_n416 )  ;
assign n1294 = state_in[87:80] ;
assign n1295 =  ( n1294 ) == ( bv_8_121_n470 )  ;
assign n1296 = state_in[87:80] ;
assign n1297 =  ( n1296 ) == ( bv_8_120_n474 )  ;
assign n1298 = state_in[87:80] ;
assign n1299 =  ( n1298 ) == ( bv_8_119_n472 )  ;
assign n1300 = state_in[87:80] ;
assign n1301 =  ( n1300 ) == ( bv_8_118_n480 )  ;
assign n1302 = state_in[87:80] ;
assign n1303 =  ( n1302 ) == ( bv_8_117_n484 )  ;
assign n1304 = state_in[87:80] ;
assign n1305 =  ( n1304 ) == ( bv_8_116_n345 )  ;
assign n1306 = state_in[87:80] ;
assign n1307 =  ( n1306 ) == ( bv_8_115_n222 )  ;
assign n1308 = state_in[87:80] ;
assign n1309 =  ( n1308 ) == ( bv_8_114_n494 )  ;
assign n1310 = state_in[87:80] ;
assign n1311 =  ( n1310 ) == ( bv_8_113_n180 )  ;
assign n1312 = state_in[87:80] ;
assign n1313 =  ( n1312 ) == ( bv_8_112_n482 )  ;
assign n1314 = state_in[87:80] ;
assign n1315 =  ( n1314 ) == ( bv_8_111_n244 )  ;
assign n1316 = state_in[87:80] ;
assign n1317 =  ( n1316 ) == ( bv_8_110_n294 )  ;
assign n1318 = state_in[87:80] ;
assign n1319 =  ( n1318 ) == ( bv_8_109_n9 )  ;
assign n1320 = state_in[87:80] ;
assign n1321 =  ( n1320 ) == ( bv_8_108_n510 )  ;
assign n1322 = state_in[87:80] ;
assign n1323 =  ( n1322 ) == ( bv_8_107_n370 )  ;
assign n1324 = state_in[87:80] ;
assign n1325 =  ( n1324 ) == ( bv_8_106_n155 )  ;
assign n1326 = state_in[87:80] ;
assign n1327 =  ( n1326 ) == ( bv_8_105_n148 )  ;
assign n1328 = state_in[87:80] ;
assign n1329 =  ( n1328 ) == ( bv_8_104_n520 )  ;
assign n1330 = state_in[87:80] ;
assign n1331 =  ( n1330 ) == ( bv_8_103_n523 )  ;
assign n1332 = state_in[87:80] ;
assign n1333 =  ( n1332 ) == ( bv_8_102_n527 )  ;
assign n1334 = state_in[87:80] ;
assign n1335 =  ( n1334 ) == ( bv_8_101_n49 )  ;
assign n1336 = state_in[87:80] ;
assign n1337 =  ( n1336 ) == ( bv_8_100_n348 )  ;
assign n1338 = state_in[87:80] ;
assign n1339 =  ( n1338 ) == ( bv_8_99_n476 )  ;
assign n1340 = state_in[87:80] ;
assign n1341 =  ( n1340 ) == ( bv_8_98_n536 )  ;
assign n1342 = state_in[87:80] ;
assign n1343 =  ( n1342 ) == ( bv_8_97_n198 )  ;
assign n1344 = state_in[87:80] ;
assign n1345 =  ( n1344 ) == ( bv_8_96_n542 )  ;
assign n1346 = state_in[87:80] ;
assign n1347 =  ( n1346 ) == ( bv_8_95_n545 )  ;
assign n1348 = state_in[87:80] ;
assign n1349 =  ( n1348 ) == ( bv_8_94_n548 )  ;
assign n1350 = state_in[87:80] ;
assign n1351 =  ( n1350 ) == ( bv_8_93_n498 )  ;
assign n1352 = state_in[87:80] ;
assign n1353 =  ( n1352 ) == ( bv_8_92_n234 )  ;
assign n1354 = state_in[87:80] ;
assign n1355 =  ( n1354 ) == ( bv_8_91_n555 )  ;
assign n1356 = state_in[87:80] ;
assign n1357 =  ( n1356 ) == ( bv_8_90_n25 )  ;
assign n1358 = state_in[87:80] ;
assign n1359 =  ( n1358 ) == ( bv_8_89_n61 )  ;
assign n1360 = state_in[87:80] ;
assign n1361 =  ( n1360 ) == ( bv_8_88_n562 )  ;
assign n1362 = state_in[87:80] ;
assign n1363 =  ( n1362 ) == ( bv_8_87_n226 )  ;
assign n1364 = state_in[87:80] ;
assign n1365 =  ( n1364 ) == ( bv_8_86_n567 )  ;
assign n1366 = state_in[87:80] ;
assign n1367 =  ( n1366 ) == ( bv_8_85_n423 )  ;
assign n1368 = state_in[87:80] ;
assign n1369 =  ( n1368 ) == ( bv_8_84_n386 )  ;
assign n1370 = state_in[87:80] ;
assign n1371 =  ( n1370 ) == ( bv_8_83_n575 )  ;
assign n1372 = state_in[87:80] ;
assign n1373 =  ( n1372 ) == ( bv_8_82_n578 )  ;
assign n1374 = state_in[87:80] ;
assign n1375 =  ( n1374 ) == ( bv_8_81_n582 )  ;
assign n1376 = state_in[87:80] ;
assign n1377 =  ( n1376 ) == ( bv_8_80_n73 )  ;
assign n1378 = state_in[87:80] ;
assign n1379 =  ( n1378 ) == ( bv_8_79_n538 )  ;
assign n1380 = state_in[87:80] ;
assign n1381 =  ( n1380 ) == ( bv_8_78_n590 )  ;
assign n1382 = state_in[87:80] ;
assign n1383 =  ( n1382 ) == ( bv_8_77_n593 )  ;
assign n1384 = state_in[87:80] ;
assign n1385 =  ( n1384 ) == ( bv_8_76_n596 )  ;
assign n1386 = state_in[87:80] ;
assign n1387 =  ( n1386 ) == ( bv_8_75_n503 )  ;
assign n1388 = state_in[87:80] ;
assign n1389 =  ( n1388 ) == ( bv_8_74_n237 )  ;
assign n1390 = state_in[87:80] ;
assign n1391 =  ( n1390 ) == ( bv_8_73_n275 )  ;
assign n1392 = state_in[87:80] ;
assign n1393 =  ( n1392 ) == ( bv_8_72_n330 )  ;
assign n1394 = state_in[87:80] ;
assign n1395 =  ( n1394 ) == ( bv_8_71_n252 )  ;
assign n1396 = state_in[87:80] ;
assign n1397 =  ( n1396 ) == ( bv_8_70_n609 )  ;
assign n1398 = state_in[87:80] ;
assign n1399 =  ( n1398 ) == ( bv_8_69_n612 )  ;
assign n1400 = state_in[87:80] ;
assign n1401 =  ( n1400 ) == ( bv_8_68_n390 )  ;
assign n1402 = state_in[87:80] ;
assign n1403 =  ( n1402 ) == ( bv_8_67_n318 )  ;
assign n1404 = state_in[87:80] ;
assign n1405 =  ( n1404 ) == ( bv_8_66_n466 )  ;
assign n1406 = state_in[87:80] ;
assign n1407 =  ( n1406 ) == ( bv_8_65_n623 )  ;
assign n1408 = state_in[87:80] ;
assign n1409 =  ( n1408 ) == ( bv_8_64_n573 )  ;
assign n1410 = state_in[87:80] ;
assign n1411 =  ( n1410 ) == ( bv_8_63_n489 )  ;
assign n1412 = state_in[87:80] ;
assign n1413 =  ( n1412 ) == ( bv_8_62_n205 )  ;
assign n1414 = state_in[87:80] ;
assign n1415 =  ( n1414 ) == ( bv_8_61_n634 )  ;
assign n1416 = state_in[87:80] ;
assign n1417 =  ( n1416 ) == ( bv_8_60_n93 )  ;
assign n1418 = state_in[87:80] ;
assign n1419 =  ( n1418 ) == ( bv_8_59_n382 )  ;
assign n1420 = state_in[87:80] ;
assign n1421 =  ( n1420 ) == ( bv_8_58_n136 )  ;
assign n1422 = state_in[87:80] ;
assign n1423 =  ( n1422 ) == ( bv_8_57_n312 )  ;
assign n1424 = state_in[87:80] ;
assign n1425 =  ( n1424 ) == ( bv_8_56_n230 )  ;
assign n1426 = state_in[87:80] ;
assign n1427 =  ( n1426 ) == ( bv_8_55_n650 )  ;
assign n1428 = state_in[87:80] ;
assign n1429 =  ( n1428 ) == ( bv_8_54_n616 )  ;
assign n1430 = state_in[87:80] ;
assign n1431 =  ( n1430 ) == ( bv_8_53_n436 )  ;
assign n1432 = state_in[87:80] ;
assign n1433 =  ( n1432 ) == ( bv_8_52_n619 )  ;
assign n1434 = state_in[87:80] ;
assign n1435 =  ( n1434 ) == ( bv_8_51_n101 )  ;
assign n1436 = state_in[87:80] ;
assign n1437 =  ( n1436 ) == ( bv_8_50_n408 )  ;
assign n1438 = state_in[87:80] ;
assign n1439 =  ( n1438 ) == ( bv_8_49_n309 )  ;
assign n1440 = state_in[87:80] ;
assign n1441 =  ( n1440 ) == ( bv_8_48_n660 )  ;
assign n1442 = state_in[87:80] ;
assign n1443 =  ( n1442 ) == ( bv_8_47_n652 )  ;
assign n1444 = state_in[87:80] ;
assign n1445 =  ( n1444 ) == ( bv_8_46_n429 )  ;
assign n1446 = state_in[87:80] ;
assign n1447 =  ( n1446 ) == ( bv_8_45_n97 )  ;
assign n1448 = state_in[87:80] ;
assign n1449 =  ( n1448 ) == ( bv_8_44_n5 )  ;
assign n1450 = state_in[87:80] ;
assign n1451 =  ( n1450 ) == ( bv_8_43_n121 )  ;
assign n1452 = state_in[87:80] ;
assign n1453 =  ( n1452 ) == ( bv_8_42_n672 )  ;
assign n1454 = state_in[87:80] ;
assign n1455 =  ( n1454 ) == ( bv_8_41_n29 )  ;
assign n1456 = state_in[87:80] ;
assign n1457 =  ( n1456 ) == ( bv_8_40_n366 )  ;
assign n1458 = state_in[87:80] ;
assign n1459 =  ( n1458 ) == ( bv_8_39_n132 )  ;
assign n1460 = state_in[87:80] ;
assign n1461 =  ( n1460 ) == ( bv_8_38_n444 )  ;
assign n1462 = state_in[87:80] ;
assign n1463 =  ( n1462 ) == ( bv_8_37_n506 )  ;
assign n1464 = state_in[87:80] ;
assign n1465 =  ( n1464 ) == ( bv_8_36_n645 )  ;
assign n1466 = state_in[87:80] ;
assign n1467 =  ( n1466 ) == ( bv_8_35_n696 )  ;
assign n1468 = state_in[87:80] ;
assign n1469 =  ( n1468 ) == ( bv_8_34_n117 )  ;
assign n1470 = state_in[87:80] ;
assign n1471 =  ( n1470 ) == ( bv_8_33_n486 )  ;
assign n1472 = state_in[87:80] ;
assign n1473 =  ( n1472 ) == ( bv_8_32_n463 )  ;
assign n1474 = state_in[87:80] ;
assign n1475 =  ( n1474 ) == ( bv_8_31_n705 )  ;
assign n1476 = state_in[87:80] ;
assign n1477 =  ( n1476 ) == ( bv_8_30_n21 )  ;
assign n1478 = state_in[87:80] ;
assign n1479 =  ( n1478 ) == ( bv_8_29_n625 )  ;
assign n1480 = state_in[87:80] ;
assign n1481 =  ( n1480 ) == ( bv_8_28_n162 )  ;
assign n1482 = state_in[87:80] ;
assign n1483 =  ( n1482 ) == ( bv_8_27_n642 )  ;
assign n1484 = state_in[87:80] ;
assign n1485 =  ( n1484 ) == ( bv_8_26_n53 )  ;
assign n1486 = state_in[87:80] ;
assign n1487 =  ( n1486 ) == ( bv_8_25_n399 )  ;
assign n1488 = state_in[87:80] ;
assign n1489 =  ( n1488 ) == ( bv_8_24_n448 )  ;
assign n1490 = state_in[87:80] ;
assign n1491 =  ( n1490 ) == ( bv_8_23_n144 )  ;
assign n1492 = state_in[87:80] ;
assign n1493 =  ( n1492 ) == ( bv_8_22_n357 )  ;
assign n1494 = state_in[87:80] ;
assign n1495 =  ( n1494 ) == ( bv_8_21_n89 )  ;
assign n1496 = state_in[87:80] ;
assign n1497 =  ( n1496 ) == ( bv_8_20_n341 )  ;
assign n1498 = state_in[87:80] ;
assign n1499 =  ( n1498 ) == ( bv_8_19_n588 )  ;
assign n1500 = state_in[87:80] ;
assign n1501 =  ( n1500 ) == ( bv_8_18_n628 )  ;
assign n1502 = state_in[87:80] ;
assign n1503 =  ( n1502 ) == ( bv_8_17_n525 )  ;
assign n1504 = state_in[87:80] ;
assign n1505 =  ( n1504 ) == ( bv_8_16_n248 )  ;
assign n1506 = state_in[87:80] ;
assign n1507 =  ( n1506 ) == ( bv_8_15_n190 )  ;
assign n1508 = state_in[87:80] ;
assign n1509 =  ( n1508 ) == ( bv_8_14_n648 )  ;
assign n1510 = state_in[87:80] ;
assign n1511 =  ( n1510 ) == ( bv_8_13_n194 )  ;
assign n1512 = state_in[87:80] ;
assign n1513 =  ( n1512 ) == ( bv_8_12_n333 )  ;
assign n1514 = state_in[87:80] ;
assign n1515 =  ( n1514 ) == ( bv_8_11_n379 )  ;
assign n1516 = state_in[87:80] ;
assign n1517 =  ( n1516 ) == ( bv_8_10_n655 )  ;
assign n1518 = state_in[87:80] ;
assign n1519 =  ( n1518 ) == ( bv_8_9_n57 )  ;
assign n1520 = state_in[87:80] ;
assign n1521 =  ( n1520 ) == ( bv_8_8_n669 )  ;
assign n1522 = state_in[87:80] ;
assign n1523 =  ( n1522 ) == ( bv_8_7_n105 )  ;
assign n1524 = state_in[87:80] ;
assign n1525 =  ( n1524 ) == ( bv_8_6_n169 )  ;
assign n1526 = state_in[87:80] ;
assign n1527 =  ( n1526 ) == ( bv_8_5_n492 )  ;
assign n1528 = state_in[87:80] ;
assign n1529 =  ( n1528 ) == ( bv_8_4_n516 )  ;
assign n1530 = state_in[87:80] ;
assign n1531 =  ( n1530 ) == ( bv_8_3_n65 )  ;
assign n1532 = state_in[87:80] ;
assign n1533 =  ( n1532 ) == ( bv_8_2_n751 )  ;
assign n1534 = state_in[87:80] ;
assign n1535 =  ( n1534 ) == ( bv_8_1_n287 )  ;
assign n1536 = state_in[87:80] ;
assign n1537 =  ( n1536 ) == ( bv_8_0_n580 )  ;
assign n1538 =  ( n1537 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n1539 =  ( n1535 ) ? ( bv_8_124_n184 ) : ( n1538 ) ;
assign n1540 =  ( n1533 ) ? ( bv_8_119_n472 ) : ( n1539 ) ;
assign n1541 =  ( n1531 ) ? ( bv_8_123_n17 ) : ( n1540 ) ;
assign n1542 =  ( n1529 ) ? ( bv_8_242_n55 ) : ( n1541 ) ;
assign n1543 =  ( n1527 ) ? ( bv_8_107_n370 ) : ( n1542 ) ;
assign n1544 =  ( n1525 ) ? ( bv_8_111_n244 ) : ( n1543 ) ;
assign n1545 =  ( n1523 ) ? ( bv_8_197_n224 ) : ( n1544 ) ;
assign n1546 =  ( n1521 ) ? ( bv_8_48_n660 ) : ( n1545 ) ;
assign n1547 =  ( n1519 ) ? ( bv_8_1_n287 ) : ( n1546 ) ;
assign n1548 =  ( n1517 ) ? ( bv_8_103_n523 ) : ( n1547 ) ;
assign n1549 =  ( n1515 ) ? ( bv_8_43_n121 ) : ( n1548 ) ;
assign n1550 =  ( n1513 ) ? ( bv_8_254_n7 ) : ( n1549 ) ;
assign n1551 =  ( n1511 ) ? ( bv_8_215_n45 ) : ( n1550 ) ;
assign n1552 =  ( n1509 ) ? ( bv_8_171_n314 ) : ( n1551 ) ;
assign n1553 =  ( n1507 ) ? ( bv_8_118_n480 ) : ( n1552 ) ;
assign n1554 =  ( n1505 ) ? ( bv_8_202_n207 ) : ( n1553 ) ;
assign n1555 =  ( n1503 ) ? ( bv_8_130_n33 ) : ( n1554 ) ;
assign n1556 =  ( n1501 ) ? ( bv_8_201_n85 ) : ( n1555 ) ;
assign n1557 =  ( n1499 ) ? ( bv_8_125_n459 ) : ( n1556 ) ;
assign n1558 =  ( n1497 ) ? ( bv_8_250_n23 ) : ( n1557 ) ;
assign n1559 =  ( n1495 ) ? ( bv_8_89_n61 ) : ( n1558 ) ;
assign n1560 =  ( n1493 ) ? ( bv_8_71_n252 ) : ( n1559 ) ;
assign n1561 =  ( n1491 ) ? ( bv_8_240_n63 ) : ( n1560 ) ;
assign n1562 =  ( n1489 ) ? ( bv_8_173_n307 ) : ( n1561 ) ;
assign n1563 =  ( n1487 ) ? ( bv_8_212_n171 ) : ( n1562 ) ;
assign n1564 =  ( n1485 ) ? ( bv_8_162_n343 ) : ( n1563 ) ;
assign n1565 =  ( n1483 ) ? ( bv_8_175_n302 ) : ( n1564 ) ;
assign n1566 =  ( n1481 ) ? ( bv_8_156_n279 ) : ( n1565 ) ;
assign n1567 =  ( n1479 ) ? ( bv_8_164_n335 ) : ( n1566 ) ;
assign n1568 =  ( n1477 ) ? ( bv_8_114_n494 ) : ( n1567 ) ;
assign n1569 =  ( n1475 ) ? ( bv_8_192_n242 ) : ( n1568 ) ;
assign n1570 =  ( n1473 ) ? ( bv_8_183_n273 ) : ( n1569 ) ;
assign n1571 =  ( n1471 ) ? ( bv_8_253_n11 ) : ( n1570 ) ;
assign n1572 =  ( n1469 ) ? ( bv_8_147_n392 ) : ( n1571 ) ;
assign n1573 =  ( n1467 ) ? ( bv_8_38_n444 ) : ( n1572 ) ;
assign n1574 =  ( n1465 ) ? ( bv_8_54_n616 ) : ( n1573 ) ;
assign n1575 =  ( n1463 ) ? ( bv_8_63_n489 ) : ( n1574 ) ;
assign n1576 =  ( n1461 ) ? ( bv_8_247_n35 ) : ( n1575 ) ;
assign n1577 =  ( n1459 ) ? ( bv_8_204_n177 ) : ( n1576 ) ;
assign n1578 =  ( n1457 ) ? ( bv_8_52_n619 ) : ( n1577 ) ;
assign n1579 =  ( n1455 ) ? ( bv_8_165_n69 ) : ( n1578 ) ;
assign n1580 =  ( n1453 ) ? ( bv_8_229_n107 ) : ( n1579 ) ;
assign n1581 =  ( n1451 ) ? ( bv_8_241_n59 ) : ( n1580 ) ;
assign n1582 =  ( n1449 ) ? ( bv_8_113_n180 ) : ( n1581 ) ;
assign n1583 =  ( n1447 ) ? ( bv_8_216_n157 ) : ( n1582 ) ;
assign n1584 =  ( n1445 ) ? ( bv_8_49_n309 ) : ( n1583 ) ;
assign n1585 =  ( n1443 ) ? ( bv_8_21_n89 ) : ( n1584 ) ;
assign n1586 =  ( n1441 ) ? ( bv_8_4_n516 ) : ( n1585 ) ;
assign n1587 =  ( n1439 ) ? ( bv_8_199_n216 ) : ( n1586 ) ;
assign n1588 =  ( n1437 ) ? ( bv_8_35_n696 ) : ( n1587 ) ;
assign n1589 =  ( n1435 ) ? ( bv_8_195_n232 ) : ( n1588 ) ;
assign n1590 =  ( n1433 ) ? ( bv_8_24_n448 ) : ( n1589 ) ;
assign n1591 =  ( n1431 ) ? ( bv_8_150_n201 ) : ( n1590 ) ;
assign n1592 =  ( n1429 ) ? ( bv_8_5_n492 ) : ( n1591 ) ;
assign n1593 =  ( n1427 ) ? ( bv_8_154_n368 ) : ( n1592 ) ;
assign n1594 =  ( n1425 ) ? ( bv_8_7_n105 ) : ( n1593 ) ;
assign n1595 =  ( n1423 ) ? ( bv_8_18_n628 ) : ( n1594 ) ;
assign n1596 =  ( n1421 ) ? ( bv_8_128_n450 ) : ( n1595 ) ;
assign n1597 =  ( n1419 ) ? ( bv_8_226_n119 ) : ( n1596 ) ;
assign n1598 =  ( n1417 ) ? ( bv_8_235_n83 ) : ( n1597 ) ;
assign n1599 =  ( n1415 ) ? ( bv_8_39_n132 ) : ( n1598 ) ;
assign n1600 =  ( n1413 ) ? ( bv_8_178_n292 ) : ( n1599 ) ;
assign n1601 =  ( n1411 ) ? ( bv_8_117_n484 ) : ( n1600 ) ;
assign n1602 =  ( n1409 ) ? ( bv_8_9_n57 ) : ( n1601 ) ;
assign n1603 =  ( n1407 ) ? ( bv_8_131_n440 ) : ( n1602 ) ;
assign n1604 =  ( n1405 ) ? ( bv_8_44_n5 ) : ( n1603 ) ;
assign n1605 =  ( n1403 ) ? ( bv_8_26_n53 ) : ( n1604 ) ;
assign n1606 =  ( n1401 ) ? ( bv_8_27_n642 ) : ( n1605 ) ;
assign n1607 =  ( n1399 ) ? ( bv_8_110_n294 ) : ( n1606 ) ;
assign n1608 =  ( n1397 ) ? ( bv_8_90_n25 ) : ( n1607 ) ;
assign n1609 =  ( n1395 ) ? ( bv_8_160_n350 ) : ( n1608 ) ;
assign n1610 =  ( n1393 ) ? ( bv_8_82_n578 ) : ( n1609 ) ;
assign n1611 =  ( n1391 ) ? ( bv_8_59_n382 ) : ( n1610 ) ;
assign n1612 =  ( n1389 ) ? ( bv_8_214_n164 ) : ( n1611 ) ;
assign n1613 =  ( n1387 ) ? ( bv_8_179_n289 ) : ( n1612 ) ;
assign n1614 =  ( n1385 ) ? ( bv_8_41_n29 ) : ( n1613 ) ;
assign n1615 =  ( n1383 ) ? ( bv_8_227_n115 ) : ( n1614 ) ;
assign n1616 =  ( n1381 ) ? ( bv_8_47_n652 ) : ( n1615 ) ;
assign n1617 =  ( n1379 ) ? ( bv_8_132_n41 ) : ( n1616 ) ;
assign n1618 =  ( n1377 ) ? ( bv_8_83_n575 ) : ( n1617 ) ;
assign n1619 =  ( n1375 ) ? ( bv_8_209_n182 ) : ( n1618 ) ;
assign n1620 =  ( n1373 ) ? ( bv_8_0_n580 ) : ( n1619 ) ;
assign n1621 =  ( n1371 ) ? ( bv_8_237_n75 ) : ( n1620 ) ;
assign n1622 =  ( n1369 ) ? ( bv_8_32_n463 ) : ( n1621 ) ;
assign n1623 =  ( n1367 ) ? ( bv_8_252_n15 ) : ( n1622 ) ;
assign n1624 =  ( n1365 ) ? ( bv_8_177_n283 ) : ( n1623 ) ;
assign n1625 =  ( n1363 ) ? ( bv_8_91_n555 ) : ( n1624 ) ;
assign n1626 =  ( n1361 ) ? ( bv_8_106_n155 ) : ( n1625 ) ;
assign n1627 =  ( n1359 ) ? ( bv_8_203_n203 ) : ( n1626 ) ;
assign n1628 =  ( n1357 ) ? ( bv_8_190_n250 ) : ( n1627 ) ;
assign n1629 =  ( n1355 ) ? ( bv_8_57_n312 ) : ( n1628 ) ;
assign n1630 =  ( n1353 ) ? ( bv_8_74_n237 ) : ( n1629 ) ;
assign n1631 =  ( n1351 ) ? ( bv_8_76_n596 ) : ( n1630 ) ;
assign n1632 =  ( n1349 ) ? ( bv_8_88_n562 ) : ( n1631 ) ;
assign n1633 =  ( n1347 ) ? ( bv_8_207_n188 ) : ( n1632 ) ;
assign n1634 =  ( n1345 ) ? ( bv_8_208_n37 ) : ( n1633 ) ;
assign n1635 =  ( n1343 ) ? ( bv_8_239_n67 ) : ( n1634 ) ;
assign n1636 =  ( n1341 ) ? ( bv_8_170_n77 ) : ( n1635 ) ;
assign n1637 =  ( n1339 ) ? ( bv_8_251_n19 ) : ( n1636 ) ;
assign n1638 =  ( n1337 ) ? ( bv_8_67_n318 ) : ( n1637 ) ;
assign n1639 =  ( n1335 ) ? ( bv_8_77_n593 ) : ( n1638 ) ;
assign n1640 =  ( n1333 ) ? ( bv_8_51_n101 ) : ( n1639 ) ;
assign n1641 =  ( n1331 ) ? ( bv_8_133_n434 ) : ( n1640 ) ;
assign n1642 =  ( n1329 ) ? ( bv_8_69_n612 ) : ( n1641 ) ;
assign n1643 =  ( n1327 ) ? ( bv_8_249_n27 ) : ( n1642 ) ;
assign n1644 =  ( n1325 ) ? ( bv_8_2_n751 ) : ( n1643 ) ;
assign n1645 =  ( n1323 ) ? ( bv_8_127_n453 ) : ( n1644 ) ;
assign n1646 =  ( n1321 ) ? ( bv_8_80_n73 ) : ( n1645 ) ;
assign n1647 =  ( n1319 ) ? ( bv_8_60_n93 ) : ( n1646 ) ;
assign n1648 =  ( n1317 ) ? ( bv_8_159_n323 ) : ( n1647 ) ;
assign n1649 =  ( n1315 ) ? ( bv_8_168_n13 ) : ( n1648 ) ;
assign n1650 =  ( n1313 ) ? ( bv_8_81_n582 ) : ( n1649 ) ;
assign n1651 =  ( n1311 ) ? ( bv_8_163_n339 ) : ( n1650 ) ;
assign n1652 =  ( n1309 ) ? ( bv_8_64_n573 ) : ( n1651 ) ;
assign n1653 =  ( n1307 ) ? ( bv_8_143_n403 ) : ( n1652 ) ;
assign n1654 =  ( n1305 ) ? ( bv_8_146_n337 ) : ( n1653 ) ;
assign n1655 =  ( n1303 ) ? ( bv_8_157_n359 ) : ( n1654 ) ;
assign n1656 =  ( n1301 ) ? ( bv_8_56_n230 ) : ( n1655 ) ;
assign n1657 =  ( n1299 ) ? ( bv_8_245_n43 ) : ( n1656 ) ;
assign n1658 =  ( n1297 ) ? ( bv_8_188_n257 ) : ( n1657 ) ;
assign n1659 =  ( n1295 ) ? ( bv_8_182_n277 ) : ( n1658 ) ;
assign n1660 =  ( n1293 ) ? ( bv_8_218_n150 ) : ( n1659 ) ;
assign n1661 =  ( n1291 ) ? ( bv_8_33_n486 ) : ( n1660 ) ;
assign n1662 =  ( n1289 ) ? ( bv_8_16_n248 ) : ( n1661 ) ;
assign n1663 =  ( n1287 ) ? ( bv_8_255_n3 ) : ( n1662 ) ;
assign n1664 =  ( n1285 ) ? ( bv_8_243_n51 ) : ( n1663 ) ;
assign n1665 =  ( n1283 ) ? ( bv_8_210_n113 ) : ( n1664 ) ;
assign n1666 =  ( n1281 ) ? ( bv_8_205_n196 ) : ( n1665 ) ;
assign n1667 =  ( n1279 ) ? ( bv_8_12_n333 ) : ( n1666 ) ;
assign n1668 =  ( n1277 ) ? ( bv_8_19_n588 ) : ( n1667 ) ;
assign n1669 =  ( n1275 ) ? ( bv_8_236_n79 ) : ( n1668 ) ;
assign n1670 =  ( n1273 ) ? ( bv_8_95_n545 ) : ( n1669 ) ;
assign n1671 =  ( n1271 ) ? ( bv_8_151_n218 ) : ( n1670 ) ;
assign n1672 =  ( n1269 ) ? ( bv_8_68_n390 ) : ( n1671 ) ;
assign n1673 =  ( n1267 ) ? ( bv_8_23_n144 ) : ( n1672 ) ;
assign n1674 =  ( n1265 ) ? ( bv_8_196_n228 ) : ( n1673 ) ;
assign n1675 =  ( n1263 ) ? ( bv_8_167_n325 ) : ( n1674 ) ;
assign n1676 =  ( n1261 ) ? ( bv_8_126_n456 ) : ( n1675 ) ;
assign n1677 =  ( n1259 ) ? ( bv_8_61_n634 ) : ( n1676 ) ;
assign n1678 =  ( n1257 ) ? ( bv_8_100_n348 ) : ( n1677 ) ;
assign n1679 =  ( n1255 ) ? ( bv_8_93_n498 ) : ( n1678 ) ;
assign n1680 =  ( n1253 ) ? ( bv_8_25_n399 ) : ( n1679 ) ;
assign n1681 =  ( n1251 ) ? ( bv_8_115_n222 ) : ( n1680 ) ;
assign n1682 =  ( n1249 ) ? ( bv_8_96_n542 ) : ( n1681 ) ;
assign n1683 =  ( n1247 ) ? ( bv_8_129_n446 ) : ( n1682 ) ;
assign n1684 =  ( n1245 ) ? ( bv_8_79_n538 ) : ( n1683 ) ;
assign n1685 =  ( n1243 ) ? ( bv_8_220_n142 ) : ( n1684 ) ;
assign n1686 =  ( n1241 ) ? ( bv_8_34_n117 ) : ( n1685 ) ;
assign n1687 =  ( n1239 ) ? ( bv_8_42_n672 ) : ( n1686 ) ;
assign n1688 =  ( n1237 ) ? ( bv_8_144_n173 ) : ( n1687 ) ;
assign n1689 =  ( n1235 ) ? ( bv_8_136_n425 ) : ( n1688 ) ;
assign n1690 =  ( n1233 ) ? ( bv_8_70_n609 ) : ( n1689 ) ;
assign n1691 =  ( n1231 ) ? ( bv_8_238_n71 ) : ( n1690 ) ;
assign n1692 =  ( n1229 ) ? ( bv_8_184_n270 ) : ( n1691 ) ;
assign n1693 =  ( n1227 ) ? ( bv_8_20_n341 ) : ( n1692 ) ;
assign n1694 =  ( n1225 ) ? ( bv_8_222_n134 ) : ( n1693 ) ;
assign n1695 =  ( n1223 ) ? ( bv_8_94_n548 ) : ( n1694 ) ;
assign n1696 =  ( n1221 ) ? ( bv_8_11_n379 ) : ( n1695 ) ;
assign n1697 =  ( n1219 ) ? ( bv_8_219_n146 ) : ( n1696 ) ;
assign n1698 =  ( n1217 ) ? ( bv_8_224_n126 ) : ( n1697 ) ;
assign n1699 =  ( n1215 ) ? ( bv_8_50_n408 ) : ( n1698 ) ;
assign n1700 =  ( n1213 ) ? ( bv_8_58_n136 ) : ( n1699 ) ;
assign n1701 =  ( n1211 ) ? ( bv_8_10_n655 ) : ( n1700 ) ;
assign n1702 =  ( n1209 ) ? ( bv_8_73_n275 ) : ( n1701 ) ;
assign n1703 =  ( n1207 ) ? ( bv_8_6_n169 ) : ( n1702 ) ;
assign n1704 =  ( n1205 ) ? ( bv_8_36_n645 ) : ( n1703 ) ;
assign n1705 =  ( n1203 ) ? ( bv_8_92_n234 ) : ( n1704 ) ;
assign n1706 =  ( n1201 ) ? ( bv_8_194_n159 ) : ( n1705 ) ;
assign n1707 =  ( n1199 ) ? ( bv_8_211_n175 ) : ( n1706 ) ;
assign n1708 =  ( n1197 ) ? ( bv_8_172_n268 ) : ( n1707 ) ;
assign n1709 =  ( n1195 ) ? ( bv_8_98_n536 ) : ( n1708 ) ;
assign n1710 =  ( n1193 ) ? ( bv_8_145_n397 ) : ( n1709 ) ;
assign n1711 =  ( n1191 ) ? ( bv_8_149_n384 ) : ( n1710 ) ;
assign n1712 =  ( n1189 ) ? ( bv_8_228_n111 ) : ( n1711 ) ;
assign n1713 =  ( n1187 ) ? ( bv_8_121_n470 ) : ( n1712 ) ;
assign n1714 =  ( n1185 ) ? ( bv_8_231_n99 ) : ( n1713 ) ;
assign n1715 =  ( n1183 ) ? ( bv_8_200_n213 ) : ( n1714 ) ;
assign n1716 =  ( n1181 ) ? ( bv_8_55_n650 ) : ( n1715 ) ;
assign n1717 =  ( n1179 ) ? ( bv_8_109_n9 ) : ( n1716 ) ;
assign n1718 =  ( n1177 ) ? ( bv_8_141_n410 ) : ( n1717 ) ;
assign n1719 =  ( n1175 ) ? ( bv_8_213_n167 ) : ( n1718 ) ;
assign n1720 =  ( n1173 ) ? ( bv_8_78_n590 ) : ( n1719 ) ;
assign n1721 =  ( n1171 ) ? ( bv_8_169_n109 ) : ( n1720 ) ;
assign n1722 =  ( n1169 ) ? ( bv_8_108_n510 ) : ( n1721 ) ;
assign n1723 =  ( n1167 ) ? ( bv_8_86_n567 ) : ( n1722 ) ;
assign n1724 =  ( n1165 ) ? ( bv_8_244_n47 ) : ( n1723 ) ;
assign n1725 =  ( n1163 ) ? ( bv_8_234_n87 ) : ( n1724 ) ;
assign n1726 =  ( n1161 ) ? ( bv_8_101_n49 ) : ( n1725 ) ;
assign n1727 =  ( n1159 ) ? ( bv_8_122_n416 ) : ( n1726 ) ;
assign n1728 =  ( n1157 ) ? ( bv_8_174_n152 ) : ( n1727 ) ;
assign n1729 =  ( n1155 ) ? ( bv_8_8_n669 ) : ( n1728 ) ;
assign n1730 =  ( n1153 ) ? ( bv_8_186_n263 ) : ( n1729 ) ;
assign n1731 =  ( n1151 ) ? ( bv_8_120_n474 ) : ( n1730 ) ;
assign n1732 =  ( n1149 ) ? ( bv_8_37_n506 ) : ( n1731 ) ;
assign n1733 =  ( n1147 ) ? ( bv_8_46_n429 ) : ( n1732 ) ;
assign n1734 =  ( n1145 ) ? ( bv_8_28_n162 ) : ( n1733 ) ;
assign n1735 =  ( n1143 ) ? ( bv_8_166_n328 ) : ( n1734 ) ;
assign n1736 =  ( n1141 ) ? ( bv_8_180_n285 ) : ( n1735 ) ;
assign n1737 =  ( n1139 ) ? ( bv_8_198_n220 ) : ( n1736 ) ;
assign n1738 =  ( n1137 ) ? ( bv_8_232_n95 ) : ( n1737 ) ;
assign n1739 =  ( n1135 ) ? ( bv_8_221_n138 ) : ( n1738 ) ;
assign n1740 =  ( n1133 ) ? ( bv_8_116_n345 ) : ( n1739 ) ;
assign n1741 =  ( n1131 ) ? ( bv_8_31_n705 ) : ( n1740 ) ;
assign n1742 =  ( n1129 ) ? ( bv_8_75_n503 ) : ( n1741 ) ;
assign n1743 =  ( n1127 ) ? ( bv_8_189_n254 ) : ( n1742 ) ;
assign n1744 =  ( n1125 ) ? ( bv_8_139_n297 ) : ( n1743 ) ;
assign n1745 =  ( n1123 ) ? ( bv_8_138_n418 ) : ( n1744 ) ;
assign n1746 =  ( n1121 ) ? ( bv_8_112_n482 ) : ( n1745 ) ;
assign n1747 =  ( n1119 ) ? ( bv_8_62_n205 ) : ( n1746 ) ;
assign n1748 =  ( n1117 ) ? ( bv_8_181_n281 ) : ( n1747 ) ;
assign n1749 =  ( n1115 ) ? ( bv_8_102_n527 ) : ( n1748 ) ;
assign n1750 =  ( n1113 ) ? ( bv_8_72_n330 ) : ( n1749 ) ;
assign n1751 =  ( n1111 ) ? ( bv_8_3_n65 ) : ( n1750 ) ;
assign n1752 =  ( n1109 ) ? ( bv_8_246_n39 ) : ( n1751 ) ;
assign n1753 =  ( n1107 ) ? ( bv_8_14_n648 ) : ( n1752 ) ;
assign n1754 =  ( n1105 ) ? ( bv_8_97_n198 ) : ( n1753 ) ;
assign n1755 =  ( n1103 ) ? ( bv_8_53_n436 ) : ( n1754 ) ;
assign n1756 =  ( n1101 ) ? ( bv_8_87_n226 ) : ( n1755 ) ;
assign n1757 =  ( n1099 ) ? ( bv_8_185_n266 ) : ( n1756 ) ;
assign n1758 =  ( n1097 ) ? ( bv_8_134_n431 ) : ( n1757 ) ;
assign n1759 =  ( n1095 ) ? ( bv_8_193_n239 ) : ( n1758 ) ;
assign n1760 =  ( n1093 ) ? ( bv_8_29_n625 ) : ( n1759 ) ;
assign n1761 =  ( n1091 ) ? ( bv_8_158_n355 ) : ( n1760 ) ;
assign n1762 =  ( n1089 ) ? ( bv_8_225_n123 ) : ( n1761 ) ;
assign n1763 =  ( n1087 ) ? ( bv_8_248_n31 ) : ( n1762 ) ;
assign n1764 =  ( n1085 ) ? ( bv_8_152_n374 ) : ( n1763 ) ;
assign n1765 =  ( n1083 ) ? ( bv_8_17_n525 ) : ( n1764 ) ;
assign n1766 =  ( n1081 ) ? ( bv_8_105_n148 ) : ( n1765 ) ;
assign n1767 =  ( n1079 ) ? ( bv_8_217_n128 ) : ( n1766 ) ;
assign n1768 =  ( n1077 ) ? ( bv_8_142_n406 ) : ( n1767 ) ;
assign n1769 =  ( n1075 ) ? ( bv_8_148_n388 ) : ( n1768 ) ;
assign n1770 =  ( n1073 ) ? ( bv_8_155_n364 ) : ( n1769 ) ;
assign n1771 =  ( n1071 ) ? ( bv_8_30_n21 ) : ( n1770 ) ;
assign n1772 =  ( n1069 ) ? ( bv_8_135_n81 ) : ( n1771 ) ;
assign n1773 =  ( n1067 ) ? ( bv_8_233_n91 ) : ( n1772 ) ;
assign n1774 =  ( n1065 ) ? ( bv_8_206_n192 ) : ( n1773 ) ;
assign n1775 =  ( n1063 ) ? ( bv_8_85_n423 ) : ( n1774 ) ;
assign n1776 =  ( n1061 ) ? ( bv_8_40_n366 ) : ( n1775 ) ;
assign n1777 =  ( n1059 ) ? ( bv_8_223_n130 ) : ( n1776 ) ;
assign n1778 =  ( n1057 ) ? ( bv_8_140_n376 ) : ( n1777 ) ;
assign n1779 =  ( n1055 ) ? ( bv_8_161_n211 ) : ( n1778 ) ;
assign n1780 =  ( n1053 ) ? ( bv_8_137_n421 ) : ( n1779 ) ;
assign n1781 =  ( n1051 ) ? ( bv_8_13_n194 ) : ( n1780 ) ;
assign n1782 =  ( n1049 ) ? ( bv_8_191_n246 ) : ( n1781 ) ;
assign n1783 =  ( n1047 ) ? ( bv_8_230_n103 ) : ( n1782 ) ;
assign n1784 =  ( n1045 ) ? ( bv_8_66_n466 ) : ( n1783 ) ;
assign n1785 =  ( n1043 ) ? ( bv_8_104_n520 ) : ( n1784 ) ;
assign n1786 =  ( n1041 ) ? ( bv_8_65_n623 ) : ( n1785 ) ;
assign n1787 =  ( n1039 ) ? ( bv_8_153_n140 ) : ( n1786 ) ;
assign n1788 =  ( n1037 ) ? ( bv_8_45_n97 ) : ( n1787 ) ;
assign n1789 =  ( n1035 ) ? ( bv_8_15_n190 ) : ( n1788 ) ;
assign n1790 =  ( n1033 ) ? ( bv_8_176_n299 ) : ( n1789 ) ;
assign n1791 =  ( n1031 ) ? ( bv_8_84_n386 ) : ( n1790 ) ;
assign n1792 =  ( n1029 ) ? ( bv_8_187_n260 ) : ( n1791 ) ;
assign n1793 =  ( n1027 ) ? ( bv_8_22_n357 ) : ( n1792 ) ;
assign n1794 =  ( n1025 ) ^ ( n1793 )  ;
assign n1795 = state_in[87:80] ;
assign n1796 =  ( n1795 ) == ( bv_8_255_n3 )  ;
assign n1797 = state_in[87:80] ;
assign n1798 =  ( n1797 ) == ( bv_8_254_n7 )  ;
assign n1799 = state_in[87:80] ;
assign n1800 =  ( n1799 ) == ( bv_8_253_n11 )  ;
assign n1801 = state_in[87:80] ;
assign n1802 =  ( n1801 ) == ( bv_8_252_n15 )  ;
assign n1803 = state_in[87:80] ;
assign n1804 =  ( n1803 ) == ( bv_8_251_n19 )  ;
assign n1805 = state_in[87:80] ;
assign n1806 =  ( n1805 ) == ( bv_8_250_n23 )  ;
assign n1807 = state_in[87:80] ;
assign n1808 =  ( n1807 ) == ( bv_8_249_n27 )  ;
assign n1809 = state_in[87:80] ;
assign n1810 =  ( n1809 ) == ( bv_8_248_n31 )  ;
assign n1811 = state_in[87:80] ;
assign n1812 =  ( n1811 ) == ( bv_8_247_n35 )  ;
assign n1813 = state_in[87:80] ;
assign n1814 =  ( n1813 ) == ( bv_8_246_n39 )  ;
assign n1815 = state_in[87:80] ;
assign n1816 =  ( n1815 ) == ( bv_8_245_n43 )  ;
assign n1817 = state_in[87:80] ;
assign n1818 =  ( n1817 ) == ( bv_8_244_n47 )  ;
assign n1819 = state_in[87:80] ;
assign n1820 =  ( n1819 ) == ( bv_8_243_n51 )  ;
assign n1821 = state_in[87:80] ;
assign n1822 =  ( n1821 ) == ( bv_8_242_n55 )  ;
assign n1823 = state_in[87:80] ;
assign n1824 =  ( n1823 ) == ( bv_8_241_n59 )  ;
assign n1825 = state_in[87:80] ;
assign n1826 =  ( n1825 ) == ( bv_8_240_n63 )  ;
assign n1827 = state_in[87:80] ;
assign n1828 =  ( n1827 ) == ( bv_8_239_n67 )  ;
assign n1829 = state_in[87:80] ;
assign n1830 =  ( n1829 ) == ( bv_8_238_n71 )  ;
assign n1831 = state_in[87:80] ;
assign n1832 =  ( n1831 ) == ( bv_8_237_n75 )  ;
assign n1833 = state_in[87:80] ;
assign n1834 =  ( n1833 ) == ( bv_8_236_n79 )  ;
assign n1835 = state_in[87:80] ;
assign n1836 =  ( n1835 ) == ( bv_8_235_n83 )  ;
assign n1837 = state_in[87:80] ;
assign n1838 =  ( n1837 ) == ( bv_8_234_n87 )  ;
assign n1839 = state_in[87:80] ;
assign n1840 =  ( n1839 ) == ( bv_8_233_n91 )  ;
assign n1841 = state_in[87:80] ;
assign n1842 =  ( n1841 ) == ( bv_8_232_n95 )  ;
assign n1843 = state_in[87:80] ;
assign n1844 =  ( n1843 ) == ( bv_8_231_n99 )  ;
assign n1845 = state_in[87:80] ;
assign n1846 =  ( n1845 ) == ( bv_8_230_n103 )  ;
assign n1847 = state_in[87:80] ;
assign n1848 =  ( n1847 ) == ( bv_8_229_n107 )  ;
assign n1849 = state_in[87:80] ;
assign n1850 =  ( n1849 ) == ( bv_8_228_n111 )  ;
assign n1851 = state_in[87:80] ;
assign n1852 =  ( n1851 ) == ( bv_8_227_n115 )  ;
assign n1853 = state_in[87:80] ;
assign n1854 =  ( n1853 ) == ( bv_8_226_n119 )  ;
assign n1855 = state_in[87:80] ;
assign n1856 =  ( n1855 ) == ( bv_8_225_n123 )  ;
assign n1857 = state_in[87:80] ;
assign n1858 =  ( n1857 ) == ( bv_8_224_n126 )  ;
assign n1859 = state_in[87:80] ;
assign n1860 =  ( n1859 ) == ( bv_8_223_n130 )  ;
assign n1861 = state_in[87:80] ;
assign n1862 =  ( n1861 ) == ( bv_8_222_n134 )  ;
assign n1863 = state_in[87:80] ;
assign n1864 =  ( n1863 ) == ( bv_8_221_n138 )  ;
assign n1865 = state_in[87:80] ;
assign n1866 =  ( n1865 ) == ( bv_8_220_n142 )  ;
assign n1867 = state_in[87:80] ;
assign n1868 =  ( n1867 ) == ( bv_8_219_n146 )  ;
assign n1869 = state_in[87:80] ;
assign n1870 =  ( n1869 ) == ( bv_8_218_n150 )  ;
assign n1871 = state_in[87:80] ;
assign n1872 =  ( n1871 ) == ( bv_8_217_n128 )  ;
assign n1873 = state_in[87:80] ;
assign n1874 =  ( n1873 ) == ( bv_8_216_n157 )  ;
assign n1875 = state_in[87:80] ;
assign n1876 =  ( n1875 ) == ( bv_8_215_n45 )  ;
assign n1877 = state_in[87:80] ;
assign n1878 =  ( n1877 ) == ( bv_8_214_n164 )  ;
assign n1879 = state_in[87:80] ;
assign n1880 =  ( n1879 ) == ( bv_8_213_n167 )  ;
assign n1881 = state_in[87:80] ;
assign n1882 =  ( n1881 ) == ( bv_8_212_n171 )  ;
assign n1883 = state_in[87:80] ;
assign n1884 =  ( n1883 ) == ( bv_8_211_n175 )  ;
assign n1885 = state_in[87:80] ;
assign n1886 =  ( n1885 ) == ( bv_8_210_n113 )  ;
assign n1887 = state_in[87:80] ;
assign n1888 =  ( n1887 ) == ( bv_8_209_n182 )  ;
assign n1889 = state_in[87:80] ;
assign n1890 =  ( n1889 ) == ( bv_8_208_n37 )  ;
assign n1891 = state_in[87:80] ;
assign n1892 =  ( n1891 ) == ( bv_8_207_n188 )  ;
assign n1893 = state_in[87:80] ;
assign n1894 =  ( n1893 ) == ( bv_8_206_n192 )  ;
assign n1895 = state_in[87:80] ;
assign n1896 =  ( n1895 ) == ( bv_8_205_n196 )  ;
assign n1897 = state_in[87:80] ;
assign n1898 =  ( n1897 ) == ( bv_8_204_n177 )  ;
assign n1899 = state_in[87:80] ;
assign n1900 =  ( n1899 ) == ( bv_8_203_n203 )  ;
assign n1901 = state_in[87:80] ;
assign n1902 =  ( n1901 ) == ( bv_8_202_n207 )  ;
assign n1903 = state_in[87:80] ;
assign n1904 =  ( n1903 ) == ( bv_8_201_n85 )  ;
assign n1905 = state_in[87:80] ;
assign n1906 =  ( n1905 ) == ( bv_8_200_n213 )  ;
assign n1907 = state_in[87:80] ;
assign n1908 =  ( n1907 ) == ( bv_8_199_n216 )  ;
assign n1909 = state_in[87:80] ;
assign n1910 =  ( n1909 ) == ( bv_8_198_n220 )  ;
assign n1911 = state_in[87:80] ;
assign n1912 =  ( n1911 ) == ( bv_8_197_n224 )  ;
assign n1913 = state_in[87:80] ;
assign n1914 =  ( n1913 ) == ( bv_8_196_n228 )  ;
assign n1915 = state_in[87:80] ;
assign n1916 =  ( n1915 ) == ( bv_8_195_n232 )  ;
assign n1917 = state_in[87:80] ;
assign n1918 =  ( n1917 ) == ( bv_8_194_n159 )  ;
assign n1919 = state_in[87:80] ;
assign n1920 =  ( n1919 ) == ( bv_8_193_n239 )  ;
assign n1921 = state_in[87:80] ;
assign n1922 =  ( n1921 ) == ( bv_8_192_n242 )  ;
assign n1923 = state_in[87:80] ;
assign n1924 =  ( n1923 ) == ( bv_8_191_n246 )  ;
assign n1925 = state_in[87:80] ;
assign n1926 =  ( n1925 ) == ( bv_8_190_n250 )  ;
assign n1927 = state_in[87:80] ;
assign n1928 =  ( n1927 ) == ( bv_8_189_n254 )  ;
assign n1929 = state_in[87:80] ;
assign n1930 =  ( n1929 ) == ( bv_8_188_n257 )  ;
assign n1931 = state_in[87:80] ;
assign n1932 =  ( n1931 ) == ( bv_8_187_n260 )  ;
assign n1933 = state_in[87:80] ;
assign n1934 =  ( n1933 ) == ( bv_8_186_n263 )  ;
assign n1935 = state_in[87:80] ;
assign n1936 =  ( n1935 ) == ( bv_8_185_n266 )  ;
assign n1937 = state_in[87:80] ;
assign n1938 =  ( n1937 ) == ( bv_8_184_n270 )  ;
assign n1939 = state_in[87:80] ;
assign n1940 =  ( n1939 ) == ( bv_8_183_n273 )  ;
assign n1941 = state_in[87:80] ;
assign n1942 =  ( n1941 ) == ( bv_8_182_n277 )  ;
assign n1943 = state_in[87:80] ;
assign n1944 =  ( n1943 ) == ( bv_8_181_n281 )  ;
assign n1945 = state_in[87:80] ;
assign n1946 =  ( n1945 ) == ( bv_8_180_n285 )  ;
assign n1947 = state_in[87:80] ;
assign n1948 =  ( n1947 ) == ( bv_8_179_n289 )  ;
assign n1949 = state_in[87:80] ;
assign n1950 =  ( n1949 ) == ( bv_8_178_n292 )  ;
assign n1951 = state_in[87:80] ;
assign n1952 =  ( n1951 ) == ( bv_8_177_n283 )  ;
assign n1953 = state_in[87:80] ;
assign n1954 =  ( n1953 ) == ( bv_8_176_n299 )  ;
assign n1955 = state_in[87:80] ;
assign n1956 =  ( n1955 ) == ( bv_8_175_n302 )  ;
assign n1957 = state_in[87:80] ;
assign n1958 =  ( n1957 ) == ( bv_8_174_n152 )  ;
assign n1959 = state_in[87:80] ;
assign n1960 =  ( n1959 ) == ( bv_8_173_n307 )  ;
assign n1961 = state_in[87:80] ;
assign n1962 =  ( n1961 ) == ( bv_8_172_n268 )  ;
assign n1963 = state_in[87:80] ;
assign n1964 =  ( n1963 ) == ( bv_8_171_n314 )  ;
assign n1965 = state_in[87:80] ;
assign n1966 =  ( n1965 ) == ( bv_8_170_n77 )  ;
assign n1967 = state_in[87:80] ;
assign n1968 =  ( n1967 ) == ( bv_8_169_n109 )  ;
assign n1969 = state_in[87:80] ;
assign n1970 =  ( n1969 ) == ( bv_8_168_n13 )  ;
assign n1971 = state_in[87:80] ;
assign n1972 =  ( n1971 ) == ( bv_8_167_n325 )  ;
assign n1973 = state_in[87:80] ;
assign n1974 =  ( n1973 ) == ( bv_8_166_n328 )  ;
assign n1975 = state_in[87:80] ;
assign n1976 =  ( n1975 ) == ( bv_8_165_n69 )  ;
assign n1977 = state_in[87:80] ;
assign n1978 =  ( n1977 ) == ( bv_8_164_n335 )  ;
assign n1979 = state_in[87:80] ;
assign n1980 =  ( n1979 ) == ( bv_8_163_n339 )  ;
assign n1981 = state_in[87:80] ;
assign n1982 =  ( n1981 ) == ( bv_8_162_n343 )  ;
assign n1983 = state_in[87:80] ;
assign n1984 =  ( n1983 ) == ( bv_8_161_n211 )  ;
assign n1985 = state_in[87:80] ;
assign n1986 =  ( n1985 ) == ( bv_8_160_n350 )  ;
assign n1987 = state_in[87:80] ;
assign n1988 =  ( n1987 ) == ( bv_8_159_n323 )  ;
assign n1989 = state_in[87:80] ;
assign n1990 =  ( n1989 ) == ( bv_8_158_n355 )  ;
assign n1991 = state_in[87:80] ;
assign n1992 =  ( n1991 ) == ( bv_8_157_n359 )  ;
assign n1993 = state_in[87:80] ;
assign n1994 =  ( n1993 ) == ( bv_8_156_n279 )  ;
assign n1995 = state_in[87:80] ;
assign n1996 =  ( n1995 ) == ( bv_8_155_n364 )  ;
assign n1997 = state_in[87:80] ;
assign n1998 =  ( n1997 ) == ( bv_8_154_n368 )  ;
assign n1999 = state_in[87:80] ;
assign n2000 =  ( n1999 ) == ( bv_8_153_n140 )  ;
assign n2001 = state_in[87:80] ;
assign n2002 =  ( n2001 ) == ( bv_8_152_n374 )  ;
assign n2003 = state_in[87:80] ;
assign n2004 =  ( n2003 ) == ( bv_8_151_n218 )  ;
assign n2005 = state_in[87:80] ;
assign n2006 =  ( n2005 ) == ( bv_8_150_n201 )  ;
assign n2007 = state_in[87:80] ;
assign n2008 =  ( n2007 ) == ( bv_8_149_n384 )  ;
assign n2009 = state_in[87:80] ;
assign n2010 =  ( n2009 ) == ( bv_8_148_n388 )  ;
assign n2011 = state_in[87:80] ;
assign n2012 =  ( n2011 ) == ( bv_8_147_n392 )  ;
assign n2013 = state_in[87:80] ;
assign n2014 =  ( n2013 ) == ( bv_8_146_n337 )  ;
assign n2015 = state_in[87:80] ;
assign n2016 =  ( n2015 ) == ( bv_8_145_n397 )  ;
assign n2017 = state_in[87:80] ;
assign n2018 =  ( n2017 ) == ( bv_8_144_n173 )  ;
assign n2019 = state_in[87:80] ;
assign n2020 =  ( n2019 ) == ( bv_8_143_n403 )  ;
assign n2021 = state_in[87:80] ;
assign n2022 =  ( n2021 ) == ( bv_8_142_n406 )  ;
assign n2023 = state_in[87:80] ;
assign n2024 =  ( n2023 ) == ( bv_8_141_n410 )  ;
assign n2025 = state_in[87:80] ;
assign n2026 =  ( n2025 ) == ( bv_8_140_n376 )  ;
assign n2027 = state_in[87:80] ;
assign n2028 =  ( n2027 ) == ( bv_8_139_n297 )  ;
assign n2029 = state_in[87:80] ;
assign n2030 =  ( n2029 ) == ( bv_8_138_n418 )  ;
assign n2031 = state_in[87:80] ;
assign n2032 =  ( n2031 ) == ( bv_8_137_n421 )  ;
assign n2033 = state_in[87:80] ;
assign n2034 =  ( n2033 ) == ( bv_8_136_n425 )  ;
assign n2035 = state_in[87:80] ;
assign n2036 =  ( n2035 ) == ( bv_8_135_n81 )  ;
assign n2037 = state_in[87:80] ;
assign n2038 =  ( n2037 ) == ( bv_8_134_n431 )  ;
assign n2039 = state_in[87:80] ;
assign n2040 =  ( n2039 ) == ( bv_8_133_n434 )  ;
assign n2041 = state_in[87:80] ;
assign n2042 =  ( n2041 ) == ( bv_8_132_n41 )  ;
assign n2043 = state_in[87:80] ;
assign n2044 =  ( n2043 ) == ( bv_8_131_n440 )  ;
assign n2045 = state_in[87:80] ;
assign n2046 =  ( n2045 ) == ( bv_8_130_n33 )  ;
assign n2047 = state_in[87:80] ;
assign n2048 =  ( n2047 ) == ( bv_8_129_n446 )  ;
assign n2049 = state_in[87:80] ;
assign n2050 =  ( n2049 ) == ( bv_8_128_n450 )  ;
assign n2051 = state_in[87:80] ;
assign n2052 =  ( n2051 ) == ( bv_8_127_n453 )  ;
assign n2053 = state_in[87:80] ;
assign n2054 =  ( n2053 ) == ( bv_8_126_n456 )  ;
assign n2055 = state_in[87:80] ;
assign n2056 =  ( n2055 ) == ( bv_8_125_n459 )  ;
assign n2057 = state_in[87:80] ;
assign n2058 =  ( n2057 ) == ( bv_8_124_n184 )  ;
assign n2059 = state_in[87:80] ;
assign n2060 =  ( n2059 ) == ( bv_8_123_n17 )  ;
assign n2061 = state_in[87:80] ;
assign n2062 =  ( n2061 ) == ( bv_8_122_n416 )  ;
assign n2063 = state_in[87:80] ;
assign n2064 =  ( n2063 ) == ( bv_8_121_n470 )  ;
assign n2065 = state_in[87:80] ;
assign n2066 =  ( n2065 ) == ( bv_8_120_n474 )  ;
assign n2067 = state_in[87:80] ;
assign n2068 =  ( n2067 ) == ( bv_8_119_n472 )  ;
assign n2069 = state_in[87:80] ;
assign n2070 =  ( n2069 ) == ( bv_8_118_n480 )  ;
assign n2071 = state_in[87:80] ;
assign n2072 =  ( n2071 ) == ( bv_8_117_n484 )  ;
assign n2073 = state_in[87:80] ;
assign n2074 =  ( n2073 ) == ( bv_8_116_n345 )  ;
assign n2075 = state_in[87:80] ;
assign n2076 =  ( n2075 ) == ( bv_8_115_n222 )  ;
assign n2077 = state_in[87:80] ;
assign n2078 =  ( n2077 ) == ( bv_8_114_n494 )  ;
assign n2079 = state_in[87:80] ;
assign n2080 =  ( n2079 ) == ( bv_8_113_n180 )  ;
assign n2081 = state_in[87:80] ;
assign n2082 =  ( n2081 ) == ( bv_8_112_n482 )  ;
assign n2083 = state_in[87:80] ;
assign n2084 =  ( n2083 ) == ( bv_8_111_n244 )  ;
assign n2085 = state_in[87:80] ;
assign n2086 =  ( n2085 ) == ( bv_8_110_n294 )  ;
assign n2087 = state_in[87:80] ;
assign n2088 =  ( n2087 ) == ( bv_8_109_n9 )  ;
assign n2089 = state_in[87:80] ;
assign n2090 =  ( n2089 ) == ( bv_8_108_n510 )  ;
assign n2091 = state_in[87:80] ;
assign n2092 =  ( n2091 ) == ( bv_8_107_n370 )  ;
assign n2093 = state_in[87:80] ;
assign n2094 =  ( n2093 ) == ( bv_8_106_n155 )  ;
assign n2095 = state_in[87:80] ;
assign n2096 =  ( n2095 ) == ( bv_8_105_n148 )  ;
assign n2097 = state_in[87:80] ;
assign n2098 =  ( n2097 ) == ( bv_8_104_n520 )  ;
assign n2099 = state_in[87:80] ;
assign n2100 =  ( n2099 ) == ( bv_8_103_n523 )  ;
assign n2101 = state_in[87:80] ;
assign n2102 =  ( n2101 ) == ( bv_8_102_n527 )  ;
assign n2103 = state_in[87:80] ;
assign n2104 =  ( n2103 ) == ( bv_8_101_n49 )  ;
assign n2105 = state_in[87:80] ;
assign n2106 =  ( n2105 ) == ( bv_8_100_n348 )  ;
assign n2107 = state_in[87:80] ;
assign n2108 =  ( n2107 ) == ( bv_8_99_n476 )  ;
assign n2109 = state_in[87:80] ;
assign n2110 =  ( n2109 ) == ( bv_8_98_n536 )  ;
assign n2111 = state_in[87:80] ;
assign n2112 =  ( n2111 ) == ( bv_8_97_n198 )  ;
assign n2113 = state_in[87:80] ;
assign n2114 =  ( n2113 ) == ( bv_8_96_n542 )  ;
assign n2115 = state_in[87:80] ;
assign n2116 =  ( n2115 ) == ( bv_8_95_n545 )  ;
assign n2117 = state_in[87:80] ;
assign n2118 =  ( n2117 ) == ( bv_8_94_n548 )  ;
assign n2119 = state_in[87:80] ;
assign n2120 =  ( n2119 ) == ( bv_8_93_n498 )  ;
assign n2121 = state_in[87:80] ;
assign n2122 =  ( n2121 ) == ( bv_8_92_n234 )  ;
assign n2123 = state_in[87:80] ;
assign n2124 =  ( n2123 ) == ( bv_8_91_n555 )  ;
assign n2125 = state_in[87:80] ;
assign n2126 =  ( n2125 ) == ( bv_8_90_n25 )  ;
assign n2127 = state_in[87:80] ;
assign n2128 =  ( n2127 ) == ( bv_8_89_n61 )  ;
assign n2129 = state_in[87:80] ;
assign n2130 =  ( n2129 ) == ( bv_8_88_n562 )  ;
assign n2131 = state_in[87:80] ;
assign n2132 =  ( n2131 ) == ( bv_8_87_n226 )  ;
assign n2133 = state_in[87:80] ;
assign n2134 =  ( n2133 ) == ( bv_8_86_n567 )  ;
assign n2135 = state_in[87:80] ;
assign n2136 =  ( n2135 ) == ( bv_8_85_n423 )  ;
assign n2137 = state_in[87:80] ;
assign n2138 =  ( n2137 ) == ( bv_8_84_n386 )  ;
assign n2139 = state_in[87:80] ;
assign n2140 =  ( n2139 ) == ( bv_8_83_n575 )  ;
assign n2141 = state_in[87:80] ;
assign n2142 =  ( n2141 ) == ( bv_8_82_n578 )  ;
assign n2143 = state_in[87:80] ;
assign n2144 =  ( n2143 ) == ( bv_8_81_n582 )  ;
assign n2145 = state_in[87:80] ;
assign n2146 =  ( n2145 ) == ( bv_8_80_n73 )  ;
assign n2147 = state_in[87:80] ;
assign n2148 =  ( n2147 ) == ( bv_8_79_n538 )  ;
assign n2149 = state_in[87:80] ;
assign n2150 =  ( n2149 ) == ( bv_8_78_n590 )  ;
assign n2151 = state_in[87:80] ;
assign n2152 =  ( n2151 ) == ( bv_8_77_n593 )  ;
assign n2153 = state_in[87:80] ;
assign n2154 =  ( n2153 ) == ( bv_8_76_n596 )  ;
assign n2155 = state_in[87:80] ;
assign n2156 =  ( n2155 ) == ( bv_8_75_n503 )  ;
assign n2157 = state_in[87:80] ;
assign n2158 =  ( n2157 ) == ( bv_8_74_n237 )  ;
assign n2159 = state_in[87:80] ;
assign n2160 =  ( n2159 ) == ( bv_8_73_n275 )  ;
assign n2161 = state_in[87:80] ;
assign n2162 =  ( n2161 ) == ( bv_8_72_n330 )  ;
assign n2163 = state_in[87:80] ;
assign n2164 =  ( n2163 ) == ( bv_8_71_n252 )  ;
assign n2165 = state_in[87:80] ;
assign n2166 =  ( n2165 ) == ( bv_8_70_n609 )  ;
assign n2167 = state_in[87:80] ;
assign n2168 =  ( n2167 ) == ( bv_8_69_n612 )  ;
assign n2169 = state_in[87:80] ;
assign n2170 =  ( n2169 ) == ( bv_8_68_n390 )  ;
assign n2171 = state_in[87:80] ;
assign n2172 =  ( n2171 ) == ( bv_8_67_n318 )  ;
assign n2173 = state_in[87:80] ;
assign n2174 =  ( n2173 ) == ( bv_8_66_n466 )  ;
assign n2175 = state_in[87:80] ;
assign n2176 =  ( n2175 ) == ( bv_8_65_n623 )  ;
assign n2177 = state_in[87:80] ;
assign n2178 =  ( n2177 ) == ( bv_8_64_n573 )  ;
assign n2179 = state_in[87:80] ;
assign n2180 =  ( n2179 ) == ( bv_8_63_n489 )  ;
assign n2181 = state_in[87:80] ;
assign n2182 =  ( n2181 ) == ( bv_8_62_n205 )  ;
assign n2183 = state_in[87:80] ;
assign n2184 =  ( n2183 ) == ( bv_8_61_n634 )  ;
assign n2185 = state_in[87:80] ;
assign n2186 =  ( n2185 ) == ( bv_8_60_n93 )  ;
assign n2187 = state_in[87:80] ;
assign n2188 =  ( n2187 ) == ( bv_8_59_n382 )  ;
assign n2189 = state_in[87:80] ;
assign n2190 =  ( n2189 ) == ( bv_8_58_n136 )  ;
assign n2191 = state_in[87:80] ;
assign n2192 =  ( n2191 ) == ( bv_8_57_n312 )  ;
assign n2193 = state_in[87:80] ;
assign n2194 =  ( n2193 ) == ( bv_8_56_n230 )  ;
assign n2195 = state_in[87:80] ;
assign n2196 =  ( n2195 ) == ( bv_8_55_n650 )  ;
assign n2197 = state_in[87:80] ;
assign n2198 =  ( n2197 ) == ( bv_8_54_n616 )  ;
assign n2199 = state_in[87:80] ;
assign n2200 =  ( n2199 ) == ( bv_8_53_n436 )  ;
assign n2201 = state_in[87:80] ;
assign n2202 =  ( n2201 ) == ( bv_8_52_n619 )  ;
assign n2203 = state_in[87:80] ;
assign n2204 =  ( n2203 ) == ( bv_8_51_n101 )  ;
assign n2205 = state_in[87:80] ;
assign n2206 =  ( n2205 ) == ( bv_8_50_n408 )  ;
assign n2207 = state_in[87:80] ;
assign n2208 =  ( n2207 ) == ( bv_8_49_n309 )  ;
assign n2209 = state_in[87:80] ;
assign n2210 =  ( n2209 ) == ( bv_8_48_n660 )  ;
assign n2211 = state_in[87:80] ;
assign n2212 =  ( n2211 ) == ( bv_8_47_n652 )  ;
assign n2213 = state_in[87:80] ;
assign n2214 =  ( n2213 ) == ( bv_8_46_n429 )  ;
assign n2215 = state_in[87:80] ;
assign n2216 =  ( n2215 ) == ( bv_8_45_n97 )  ;
assign n2217 = state_in[87:80] ;
assign n2218 =  ( n2217 ) == ( bv_8_44_n5 )  ;
assign n2219 = state_in[87:80] ;
assign n2220 =  ( n2219 ) == ( bv_8_43_n121 )  ;
assign n2221 = state_in[87:80] ;
assign n2222 =  ( n2221 ) == ( bv_8_42_n672 )  ;
assign n2223 = state_in[87:80] ;
assign n2224 =  ( n2223 ) == ( bv_8_41_n29 )  ;
assign n2225 = state_in[87:80] ;
assign n2226 =  ( n2225 ) == ( bv_8_40_n366 )  ;
assign n2227 = state_in[87:80] ;
assign n2228 =  ( n2227 ) == ( bv_8_39_n132 )  ;
assign n2229 = state_in[87:80] ;
assign n2230 =  ( n2229 ) == ( bv_8_38_n444 )  ;
assign n2231 = state_in[87:80] ;
assign n2232 =  ( n2231 ) == ( bv_8_37_n506 )  ;
assign n2233 = state_in[87:80] ;
assign n2234 =  ( n2233 ) == ( bv_8_36_n645 )  ;
assign n2235 = state_in[87:80] ;
assign n2236 =  ( n2235 ) == ( bv_8_35_n696 )  ;
assign n2237 = state_in[87:80] ;
assign n2238 =  ( n2237 ) == ( bv_8_34_n117 )  ;
assign n2239 = state_in[87:80] ;
assign n2240 =  ( n2239 ) == ( bv_8_33_n486 )  ;
assign n2241 = state_in[87:80] ;
assign n2242 =  ( n2241 ) == ( bv_8_32_n463 )  ;
assign n2243 = state_in[87:80] ;
assign n2244 =  ( n2243 ) == ( bv_8_31_n705 )  ;
assign n2245 = state_in[87:80] ;
assign n2246 =  ( n2245 ) == ( bv_8_30_n21 )  ;
assign n2247 = state_in[87:80] ;
assign n2248 =  ( n2247 ) == ( bv_8_29_n625 )  ;
assign n2249 = state_in[87:80] ;
assign n2250 =  ( n2249 ) == ( bv_8_28_n162 )  ;
assign n2251 = state_in[87:80] ;
assign n2252 =  ( n2251 ) == ( bv_8_27_n642 )  ;
assign n2253 = state_in[87:80] ;
assign n2254 =  ( n2253 ) == ( bv_8_26_n53 )  ;
assign n2255 = state_in[87:80] ;
assign n2256 =  ( n2255 ) == ( bv_8_25_n399 )  ;
assign n2257 = state_in[87:80] ;
assign n2258 =  ( n2257 ) == ( bv_8_24_n448 )  ;
assign n2259 = state_in[87:80] ;
assign n2260 =  ( n2259 ) == ( bv_8_23_n144 )  ;
assign n2261 = state_in[87:80] ;
assign n2262 =  ( n2261 ) == ( bv_8_22_n357 )  ;
assign n2263 = state_in[87:80] ;
assign n2264 =  ( n2263 ) == ( bv_8_21_n89 )  ;
assign n2265 = state_in[87:80] ;
assign n2266 =  ( n2265 ) == ( bv_8_20_n341 )  ;
assign n2267 = state_in[87:80] ;
assign n2268 =  ( n2267 ) == ( bv_8_19_n588 )  ;
assign n2269 = state_in[87:80] ;
assign n2270 =  ( n2269 ) == ( bv_8_18_n628 )  ;
assign n2271 = state_in[87:80] ;
assign n2272 =  ( n2271 ) == ( bv_8_17_n525 )  ;
assign n2273 = state_in[87:80] ;
assign n2274 =  ( n2273 ) == ( bv_8_16_n248 )  ;
assign n2275 = state_in[87:80] ;
assign n2276 =  ( n2275 ) == ( bv_8_15_n190 )  ;
assign n2277 = state_in[87:80] ;
assign n2278 =  ( n2277 ) == ( bv_8_14_n648 )  ;
assign n2279 = state_in[87:80] ;
assign n2280 =  ( n2279 ) == ( bv_8_13_n194 )  ;
assign n2281 = state_in[87:80] ;
assign n2282 =  ( n2281 ) == ( bv_8_12_n333 )  ;
assign n2283 = state_in[87:80] ;
assign n2284 =  ( n2283 ) == ( bv_8_11_n379 )  ;
assign n2285 = state_in[87:80] ;
assign n2286 =  ( n2285 ) == ( bv_8_10_n655 )  ;
assign n2287 = state_in[87:80] ;
assign n2288 =  ( n2287 ) == ( bv_8_9_n57 )  ;
assign n2289 = state_in[87:80] ;
assign n2290 =  ( n2289 ) == ( bv_8_8_n669 )  ;
assign n2291 = state_in[87:80] ;
assign n2292 =  ( n2291 ) == ( bv_8_7_n105 )  ;
assign n2293 = state_in[87:80] ;
assign n2294 =  ( n2293 ) == ( bv_8_6_n169 )  ;
assign n2295 = state_in[87:80] ;
assign n2296 =  ( n2295 ) == ( bv_8_5_n492 )  ;
assign n2297 = state_in[87:80] ;
assign n2298 =  ( n2297 ) == ( bv_8_4_n516 )  ;
assign n2299 = state_in[87:80] ;
assign n2300 =  ( n2299 ) == ( bv_8_3_n65 )  ;
assign n2301 = state_in[87:80] ;
assign n2302 =  ( n2301 ) == ( bv_8_2_n751 )  ;
assign n2303 = state_in[87:80] ;
assign n2304 =  ( n2303 ) == ( bv_8_1_n287 )  ;
assign n2305 = state_in[87:80] ;
assign n2306 =  ( n2305 ) == ( bv_8_0_n580 )  ;
assign n2307 =  ( n2306 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n2308 =  ( n2304 ) ? ( bv_8_248_n31 ) : ( n2307 ) ;
assign n2309 =  ( n2302 ) ? ( bv_8_238_n71 ) : ( n2308 ) ;
assign n2310 =  ( n2300 ) ? ( bv_8_246_n39 ) : ( n2309 ) ;
assign n2311 =  ( n2298 ) ? ( bv_8_255_n3 ) : ( n2310 ) ;
assign n2312 =  ( n2296 ) ? ( bv_8_214_n164 ) : ( n2311 ) ;
assign n2313 =  ( n2294 ) ? ( bv_8_222_n134 ) : ( n2312 ) ;
assign n2314 =  ( n2292 ) ? ( bv_8_145_n397 ) : ( n2313 ) ;
assign n2315 =  ( n2290 ) ? ( bv_8_96_n542 ) : ( n2314 ) ;
assign n2316 =  ( n2288 ) ? ( bv_8_2_n751 ) : ( n2315 ) ;
assign n2317 =  ( n2286 ) ? ( bv_8_206_n192 ) : ( n2316 ) ;
assign n2318 =  ( n2284 ) ? ( bv_8_86_n567 ) : ( n2317 ) ;
assign n2319 =  ( n2282 ) ? ( bv_8_231_n99 ) : ( n2318 ) ;
assign n2320 =  ( n2280 ) ? ( bv_8_181_n281 ) : ( n2319 ) ;
assign n2321 =  ( n2278 ) ? ( bv_8_77_n593 ) : ( n2320 ) ;
assign n2322 =  ( n2276 ) ? ( bv_8_236_n79 ) : ( n2321 ) ;
assign n2323 =  ( n2274 ) ? ( bv_8_143_n403 ) : ( n2322 ) ;
assign n2324 =  ( n2272 ) ? ( bv_8_31_n705 ) : ( n2323 ) ;
assign n2325 =  ( n2270 ) ? ( bv_8_137_n421 ) : ( n2324 ) ;
assign n2326 =  ( n2268 ) ? ( bv_8_250_n23 ) : ( n2325 ) ;
assign n2327 =  ( n2266 ) ? ( bv_8_239_n67 ) : ( n2326 ) ;
assign n2328 =  ( n2264 ) ? ( bv_8_178_n292 ) : ( n2327 ) ;
assign n2329 =  ( n2262 ) ? ( bv_8_142_n406 ) : ( n2328 ) ;
assign n2330 =  ( n2260 ) ? ( bv_8_251_n19 ) : ( n2329 ) ;
assign n2331 =  ( n2258 ) ? ( bv_8_65_n623 ) : ( n2330 ) ;
assign n2332 =  ( n2256 ) ? ( bv_8_179_n289 ) : ( n2331 ) ;
assign n2333 =  ( n2254 ) ? ( bv_8_95_n545 ) : ( n2332 ) ;
assign n2334 =  ( n2252 ) ? ( bv_8_69_n612 ) : ( n2333 ) ;
assign n2335 =  ( n2250 ) ? ( bv_8_35_n696 ) : ( n2334 ) ;
assign n2336 =  ( n2248 ) ? ( bv_8_83_n575 ) : ( n2335 ) ;
assign n2337 =  ( n2246 ) ? ( bv_8_228_n111 ) : ( n2336 ) ;
assign n2338 =  ( n2244 ) ? ( bv_8_155_n364 ) : ( n2337 ) ;
assign n2339 =  ( n2242 ) ? ( bv_8_117_n484 ) : ( n2338 ) ;
assign n2340 =  ( n2240 ) ? ( bv_8_225_n123 ) : ( n2339 ) ;
assign n2341 =  ( n2238 ) ? ( bv_8_61_n634 ) : ( n2340 ) ;
assign n2342 =  ( n2236 ) ? ( bv_8_76_n596 ) : ( n2341 ) ;
assign n2343 =  ( n2234 ) ? ( bv_8_108_n510 ) : ( n2342 ) ;
assign n2344 =  ( n2232 ) ? ( bv_8_126_n456 ) : ( n2343 ) ;
assign n2345 =  ( n2230 ) ? ( bv_8_245_n43 ) : ( n2344 ) ;
assign n2346 =  ( n2228 ) ? ( bv_8_131_n440 ) : ( n2345 ) ;
assign n2347 =  ( n2226 ) ? ( bv_8_104_n520 ) : ( n2346 ) ;
assign n2348 =  ( n2224 ) ? ( bv_8_81_n582 ) : ( n2347 ) ;
assign n2349 =  ( n2222 ) ? ( bv_8_209_n182 ) : ( n2348 ) ;
assign n2350 =  ( n2220 ) ? ( bv_8_249_n27 ) : ( n2349 ) ;
assign n2351 =  ( n2218 ) ? ( bv_8_226_n119 ) : ( n2350 ) ;
assign n2352 =  ( n2216 ) ? ( bv_8_171_n314 ) : ( n2351 ) ;
assign n2353 =  ( n2214 ) ? ( bv_8_98_n536 ) : ( n2352 ) ;
assign n2354 =  ( n2212 ) ? ( bv_8_42_n672 ) : ( n2353 ) ;
assign n2355 =  ( n2210 ) ? ( bv_8_8_n669 ) : ( n2354 ) ;
assign n2356 =  ( n2208 ) ? ( bv_8_149_n384 ) : ( n2355 ) ;
assign n2357 =  ( n2206 ) ? ( bv_8_70_n609 ) : ( n2356 ) ;
assign n2358 =  ( n2204 ) ? ( bv_8_157_n359 ) : ( n2357 ) ;
assign n2359 =  ( n2202 ) ? ( bv_8_48_n660 ) : ( n2358 ) ;
assign n2360 =  ( n2200 ) ? ( bv_8_55_n650 ) : ( n2359 ) ;
assign n2361 =  ( n2198 ) ? ( bv_8_10_n655 ) : ( n2360 ) ;
assign n2362 =  ( n2196 ) ? ( bv_8_47_n652 ) : ( n2361 ) ;
assign n2363 =  ( n2194 ) ? ( bv_8_14_n648 ) : ( n2362 ) ;
assign n2364 =  ( n2192 ) ? ( bv_8_36_n645 ) : ( n2363 ) ;
assign n2365 =  ( n2190 ) ? ( bv_8_27_n642 ) : ( n2364 ) ;
assign n2366 =  ( n2188 ) ? ( bv_8_223_n130 ) : ( n2365 ) ;
assign n2367 =  ( n2186 ) ? ( bv_8_205_n196 ) : ( n2366 ) ;
assign n2368 =  ( n2184 ) ? ( bv_8_78_n590 ) : ( n2367 ) ;
assign n2369 =  ( n2182 ) ? ( bv_8_127_n453 ) : ( n2368 ) ;
assign n2370 =  ( n2180 ) ? ( bv_8_234_n87 ) : ( n2369 ) ;
assign n2371 =  ( n2178 ) ? ( bv_8_18_n628 ) : ( n2370 ) ;
assign n2372 =  ( n2176 ) ? ( bv_8_29_n625 ) : ( n2371 ) ;
assign n2373 =  ( n2174 ) ? ( bv_8_88_n562 ) : ( n2372 ) ;
assign n2374 =  ( n2172 ) ? ( bv_8_52_n619 ) : ( n2373 ) ;
assign n2375 =  ( n2170 ) ? ( bv_8_54_n616 ) : ( n2374 ) ;
assign n2376 =  ( n2168 ) ? ( bv_8_220_n142 ) : ( n2375 ) ;
assign n2377 =  ( n2166 ) ? ( bv_8_180_n285 ) : ( n2376 ) ;
assign n2378 =  ( n2164 ) ? ( bv_8_91_n555 ) : ( n2377 ) ;
assign n2379 =  ( n2162 ) ? ( bv_8_164_n335 ) : ( n2378 ) ;
assign n2380 =  ( n2160 ) ? ( bv_8_118_n480 ) : ( n2379 ) ;
assign n2381 =  ( n2158 ) ? ( bv_8_183_n273 ) : ( n2380 ) ;
assign n2382 =  ( n2156 ) ? ( bv_8_125_n459 ) : ( n2381 ) ;
assign n2383 =  ( n2154 ) ? ( bv_8_82_n578 ) : ( n2382 ) ;
assign n2384 =  ( n2152 ) ? ( bv_8_221_n138 ) : ( n2383 ) ;
assign n2385 =  ( n2150 ) ? ( bv_8_94_n548 ) : ( n2384 ) ;
assign n2386 =  ( n2148 ) ? ( bv_8_19_n588 ) : ( n2385 ) ;
assign n2387 =  ( n2146 ) ? ( bv_8_166_n328 ) : ( n2386 ) ;
assign n2388 =  ( n2144 ) ? ( bv_8_185_n266 ) : ( n2387 ) ;
assign n2389 =  ( n2142 ) ? ( bv_8_0_n580 ) : ( n2388 ) ;
assign n2390 =  ( n2140 ) ? ( bv_8_193_n239 ) : ( n2389 ) ;
assign n2391 =  ( n2138 ) ? ( bv_8_64_n573 ) : ( n2390 ) ;
assign n2392 =  ( n2136 ) ? ( bv_8_227_n115 ) : ( n2391 ) ;
assign n2393 =  ( n2134 ) ? ( bv_8_121_n470 ) : ( n2392 ) ;
assign n2394 =  ( n2132 ) ? ( bv_8_182_n277 ) : ( n2393 ) ;
assign n2395 =  ( n2130 ) ? ( bv_8_212_n171 ) : ( n2394 ) ;
assign n2396 =  ( n2128 ) ? ( bv_8_141_n410 ) : ( n2395 ) ;
assign n2397 =  ( n2126 ) ? ( bv_8_103_n523 ) : ( n2396 ) ;
assign n2398 =  ( n2124 ) ? ( bv_8_114_n494 ) : ( n2397 ) ;
assign n2399 =  ( n2122 ) ? ( bv_8_148_n388 ) : ( n2398 ) ;
assign n2400 =  ( n2120 ) ? ( bv_8_152_n374 ) : ( n2399 ) ;
assign n2401 =  ( n2118 ) ? ( bv_8_176_n299 ) : ( n2400 ) ;
assign n2402 =  ( n2116 ) ? ( bv_8_133_n434 ) : ( n2401 ) ;
assign n2403 =  ( n2114 ) ? ( bv_8_187_n260 ) : ( n2402 ) ;
assign n2404 =  ( n2112 ) ? ( bv_8_197_n224 ) : ( n2403 ) ;
assign n2405 =  ( n2110 ) ? ( bv_8_79_n538 ) : ( n2404 ) ;
assign n2406 =  ( n2108 ) ? ( bv_8_237_n75 ) : ( n2405 ) ;
assign n2407 =  ( n2106 ) ? ( bv_8_134_n431 ) : ( n2406 ) ;
assign n2408 =  ( n2104 ) ? ( bv_8_154_n368 ) : ( n2407 ) ;
assign n2409 =  ( n2102 ) ? ( bv_8_102_n527 ) : ( n2408 ) ;
assign n2410 =  ( n2100 ) ? ( bv_8_17_n525 ) : ( n2409 ) ;
assign n2411 =  ( n2098 ) ? ( bv_8_138_n418 ) : ( n2410 ) ;
assign n2412 =  ( n2096 ) ? ( bv_8_233_n91 ) : ( n2411 ) ;
assign n2413 =  ( n2094 ) ? ( bv_8_4_n516 ) : ( n2412 ) ;
assign n2414 =  ( n2092 ) ? ( bv_8_254_n7 ) : ( n2413 ) ;
assign n2415 =  ( n2090 ) ? ( bv_8_160_n350 ) : ( n2414 ) ;
assign n2416 =  ( n2088 ) ? ( bv_8_120_n474 ) : ( n2415 ) ;
assign n2417 =  ( n2086 ) ? ( bv_8_37_n506 ) : ( n2416 ) ;
assign n2418 =  ( n2084 ) ? ( bv_8_75_n503 ) : ( n2417 ) ;
assign n2419 =  ( n2082 ) ? ( bv_8_162_n343 ) : ( n2418 ) ;
assign n2420 =  ( n2080 ) ? ( bv_8_93_n498 ) : ( n2419 ) ;
assign n2421 =  ( n2078 ) ? ( bv_8_128_n450 ) : ( n2420 ) ;
assign n2422 =  ( n2076 ) ? ( bv_8_5_n492 ) : ( n2421 ) ;
assign n2423 =  ( n2074 ) ? ( bv_8_63_n489 ) : ( n2422 ) ;
assign n2424 =  ( n2072 ) ? ( bv_8_33_n486 ) : ( n2423 ) ;
assign n2425 =  ( n2070 ) ? ( bv_8_112_n482 ) : ( n2424 ) ;
assign n2426 =  ( n2068 ) ? ( bv_8_241_n59 ) : ( n2425 ) ;
assign n2427 =  ( n2066 ) ? ( bv_8_99_n476 ) : ( n2426 ) ;
assign n2428 =  ( n2064 ) ? ( bv_8_119_n472 ) : ( n2427 ) ;
assign n2429 =  ( n2062 ) ? ( bv_8_175_n302 ) : ( n2428 ) ;
assign n2430 =  ( n2060 ) ? ( bv_8_66_n466 ) : ( n2429 ) ;
assign n2431 =  ( n2058 ) ? ( bv_8_32_n463 ) : ( n2430 ) ;
assign n2432 =  ( n2056 ) ? ( bv_8_229_n107 ) : ( n2431 ) ;
assign n2433 =  ( n2054 ) ? ( bv_8_253_n11 ) : ( n2432 ) ;
assign n2434 =  ( n2052 ) ? ( bv_8_191_n246 ) : ( n2433 ) ;
assign n2435 =  ( n2050 ) ? ( bv_8_129_n446 ) : ( n2434 ) ;
assign n2436 =  ( n2048 ) ? ( bv_8_24_n448 ) : ( n2435 ) ;
assign n2437 =  ( n2046 ) ? ( bv_8_38_n444 ) : ( n2436 ) ;
assign n2438 =  ( n2044 ) ? ( bv_8_195_n232 ) : ( n2437 ) ;
assign n2439 =  ( n2042 ) ? ( bv_8_190_n250 ) : ( n2438 ) ;
assign n2440 =  ( n2040 ) ? ( bv_8_53_n436 ) : ( n2439 ) ;
assign n2441 =  ( n2038 ) ? ( bv_8_136_n425 ) : ( n2440 ) ;
assign n2442 =  ( n2036 ) ? ( bv_8_46_n429 ) : ( n2441 ) ;
assign n2443 =  ( n2034 ) ? ( bv_8_147_n392 ) : ( n2442 ) ;
assign n2444 =  ( n2032 ) ? ( bv_8_85_n423 ) : ( n2443 ) ;
assign n2445 =  ( n2030 ) ? ( bv_8_252_n15 ) : ( n2444 ) ;
assign n2446 =  ( n2028 ) ? ( bv_8_122_n416 ) : ( n2445 ) ;
assign n2447 =  ( n2026 ) ? ( bv_8_200_n213 ) : ( n2446 ) ;
assign n2448 =  ( n2024 ) ? ( bv_8_186_n263 ) : ( n2447 ) ;
assign n2449 =  ( n2022 ) ? ( bv_8_50_n408 ) : ( n2448 ) ;
assign n2450 =  ( n2020 ) ? ( bv_8_230_n103 ) : ( n2449 ) ;
assign n2451 =  ( n2018 ) ? ( bv_8_192_n242 ) : ( n2450 ) ;
assign n2452 =  ( n2016 ) ? ( bv_8_25_n399 ) : ( n2451 ) ;
assign n2453 =  ( n2014 ) ? ( bv_8_158_n355 ) : ( n2452 ) ;
assign n2454 =  ( n2012 ) ? ( bv_8_163_n339 ) : ( n2453 ) ;
assign n2455 =  ( n2010 ) ? ( bv_8_68_n390 ) : ( n2454 ) ;
assign n2456 =  ( n2008 ) ? ( bv_8_84_n386 ) : ( n2455 ) ;
assign n2457 =  ( n2006 ) ? ( bv_8_59_n382 ) : ( n2456 ) ;
assign n2458 =  ( n2004 ) ? ( bv_8_11_n379 ) : ( n2457 ) ;
assign n2459 =  ( n2002 ) ? ( bv_8_140_n376 ) : ( n2458 ) ;
assign n2460 =  ( n2000 ) ? ( bv_8_199_n216 ) : ( n2459 ) ;
assign n2461 =  ( n1998 ) ? ( bv_8_107_n370 ) : ( n2460 ) ;
assign n2462 =  ( n1996 ) ? ( bv_8_40_n366 ) : ( n2461 ) ;
assign n2463 =  ( n1994 ) ? ( bv_8_167_n325 ) : ( n2462 ) ;
assign n2464 =  ( n1992 ) ? ( bv_8_188_n257 ) : ( n2463 ) ;
assign n2465 =  ( n1990 ) ? ( bv_8_22_n357 ) : ( n2464 ) ;
assign n2466 =  ( n1988 ) ? ( bv_8_173_n307 ) : ( n2465 ) ;
assign n2467 =  ( n1986 ) ? ( bv_8_219_n146 ) : ( n2466 ) ;
assign n2468 =  ( n1984 ) ? ( bv_8_100_n348 ) : ( n2467 ) ;
assign n2469 =  ( n1982 ) ? ( bv_8_116_n345 ) : ( n2468 ) ;
assign n2470 =  ( n1980 ) ? ( bv_8_20_n341 ) : ( n2469 ) ;
assign n2471 =  ( n1978 ) ? ( bv_8_146_n337 ) : ( n2470 ) ;
assign n2472 =  ( n1976 ) ? ( bv_8_12_n333 ) : ( n2471 ) ;
assign n2473 =  ( n1974 ) ? ( bv_8_72_n330 ) : ( n2472 ) ;
assign n2474 =  ( n1972 ) ? ( bv_8_184_n270 ) : ( n2473 ) ;
assign n2475 =  ( n1970 ) ? ( bv_8_159_n323 ) : ( n2474 ) ;
assign n2476 =  ( n1968 ) ? ( bv_8_189_n254 ) : ( n2475 ) ;
assign n2477 =  ( n1966 ) ? ( bv_8_67_n318 ) : ( n2476 ) ;
assign n2478 =  ( n1964 ) ? ( bv_8_196_n228 ) : ( n2477 ) ;
assign n2479 =  ( n1962 ) ? ( bv_8_57_n312 ) : ( n2478 ) ;
assign n2480 =  ( n1960 ) ? ( bv_8_49_n309 ) : ( n2479 ) ;
assign n2481 =  ( n1958 ) ? ( bv_8_211_n175 ) : ( n2480 ) ;
assign n2482 =  ( n1956 ) ? ( bv_8_242_n55 ) : ( n2481 ) ;
assign n2483 =  ( n1954 ) ? ( bv_8_213_n167 ) : ( n2482 ) ;
assign n2484 =  ( n1952 ) ? ( bv_8_139_n297 ) : ( n2483 ) ;
assign n2485 =  ( n1950 ) ? ( bv_8_110_n294 ) : ( n2484 ) ;
assign n2486 =  ( n1948 ) ? ( bv_8_218_n150 ) : ( n2485 ) ;
assign n2487 =  ( n1946 ) ? ( bv_8_1_n287 ) : ( n2486 ) ;
assign n2488 =  ( n1944 ) ? ( bv_8_177_n283 ) : ( n2487 ) ;
assign n2489 =  ( n1942 ) ? ( bv_8_156_n279 ) : ( n2488 ) ;
assign n2490 =  ( n1940 ) ? ( bv_8_73_n275 ) : ( n2489 ) ;
assign n2491 =  ( n1938 ) ? ( bv_8_216_n157 ) : ( n2490 ) ;
assign n2492 =  ( n1936 ) ? ( bv_8_172_n268 ) : ( n2491 ) ;
assign n2493 =  ( n1934 ) ? ( bv_8_243_n51 ) : ( n2492 ) ;
assign n2494 =  ( n1932 ) ? ( bv_8_207_n188 ) : ( n2493 ) ;
assign n2495 =  ( n1930 ) ? ( bv_8_202_n207 ) : ( n2494 ) ;
assign n2496 =  ( n1928 ) ? ( bv_8_244_n47 ) : ( n2495 ) ;
assign n2497 =  ( n1926 ) ? ( bv_8_71_n252 ) : ( n2496 ) ;
assign n2498 =  ( n1924 ) ? ( bv_8_16_n248 ) : ( n2497 ) ;
assign n2499 =  ( n1922 ) ? ( bv_8_111_n244 ) : ( n2498 ) ;
assign n2500 =  ( n1920 ) ? ( bv_8_240_n63 ) : ( n2499 ) ;
assign n2501 =  ( n1918 ) ? ( bv_8_74_n237 ) : ( n2500 ) ;
assign n2502 =  ( n1916 ) ? ( bv_8_92_n234 ) : ( n2501 ) ;
assign n2503 =  ( n1914 ) ? ( bv_8_56_n230 ) : ( n2502 ) ;
assign n2504 =  ( n1912 ) ? ( bv_8_87_n226 ) : ( n2503 ) ;
assign n2505 =  ( n1910 ) ? ( bv_8_115_n222 ) : ( n2504 ) ;
assign n2506 =  ( n1908 ) ? ( bv_8_151_n218 ) : ( n2505 ) ;
assign n2507 =  ( n1906 ) ? ( bv_8_203_n203 ) : ( n2506 ) ;
assign n2508 =  ( n1904 ) ? ( bv_8_161_n211 ) : ( n2507 ) ;
assign n2509 =  ( n1902 ) ? ( bv_8_232_n95 ) : ( n2508 ) ;
assign n2510 =  ( n1900 ) ? ( bv_8_62_n205 ) : ( n2509 ) ;
assign n2511 =  ( n1898 ) ? ( bv_8_150_n201 ) : ( n2510 ) ;
assign n2512 =  ( n1896 ) ? ( bv_8_97_n198 ) : ( n2511 ) ;
assign n2513 =  ( n1894 ) ? ( bv_8_13_n194 ) : ( n2512 ) ;
assign n2514 =  ( n1892 ) ? ( bv_8_15_n190 ) : ( n2513 ) ;
assign n2515 =  ( n1890 ) ? ( bv_8_224_n126 ) : ( n2514 ) ;
assign n2516 =  ( n1888 ) ? ( bv_8_124_n184 ) : ( n2515 ) ;
assign n2517 =  ( n1886 ) ? ( bv_8_113_n180 ) : ( n2516 ) ;
assign n2518 =  ( n1884 ) ? ( bv_8_204_n177 ) : ( n2517 ) ;
assign n2519 =  ( n1882 ) ? ( bv_8_144_n173 ) : ( n2518 ) ;
assign n2520 =  ( n1880 ) ? ( bv_8_6_n169 ) : ( n2519 ) ;
assign n2521 =  ( n1878 ) ? ( bv_8_247_n35 ) : ( n2520 ) ;
assign n2522 =  ( n1876 ) ? ( bv_8_28_n162 ) : ( n2521 ) ;
assign n2523 =  ( n1874 ) ? ( bv_8_194_n159 ) : ( n2522 ) ;
assign n2524 =  ( n1872 ) ? ( bv_8_106_n155 ) : ( n2523 ) ;
assign n2525 =  ( n1870 ) ? ( bv_8_174_n152 ) : ( n2524 ) ;
assign n2526 =  ( n1868 ) ? ( bv_8_105_n148 ) : ( n2525 ) ;
assign n2527 =  ( n1866 ) ? ( bv_8_23_n144 ) : ( n2526 ) ;
assign n2528 =  ( n1864 ) ? ( bv_8_153_n140 ) : ( n2527 ) ;
assign n2529 =  ( n1862 ) ? ( bv_8_58_n136 ) : ( n2528 ) ;
assign n2530 =  ( n1860 ) ? ( bv_8_39_n132 ) : ( n2529 ) ;
assign n2531 =  ( n1858 ) ? ( bv_8_217_n128 ) : ( n2530 ) ;
assign n2532 =  ( n1856 ) ? ( bv_8_235_n83 ) : ( n2531 ) ;
assign n2533 =  ( n1854 ) ? ( bv_8_43_n121 ) : ( n2532 ) ;
assign n2534 =  ( n1852 ) ? ( bv_8_34_n117 ) : ( n2533 ) ;
assign n2535 =  ( n1850 ) ? ( bv_8_210_n113 ) : ( n2534 ) ;
assign n2536 =  ( n1848 ) ? ( bv_8_169_n109 ) : ( n2535 ) ;
assign n2537 =  ( n1846 ) ? ( bv_8_7_n105 ) : ( n2536 ) ;
assign n2538 =  ( n1844 ) ? ( bv_8_51_n101 ) : ( n2537 ) ;
assign n2539 =  ( n1842 ) ? ( bv_8_45_n97 ) : ( n2538 ) ;
assign n2540 =  ( n1840 ) ? ( bv_8_60_n93 ) : ( n2539 ) ;
assign n2541 =  ( n1838 ) ? ( bv_8_21_n89 ) : ( n2540 ) ;
assign n2542 =  ( n1836 ) ? ( bv_8_201_n85 ) : ( n2541 ) ;
assign n2543 =  ( n1834 ) ? ( bv_8_135_n81 ) : ( n2542 ) ;
assign n2544 =  ( n1832 ) ? ( bv_8_170_n77 ) : ( n2543 ) ;
assign n2545 =  ( n1830 ) ? ( bv_8_80_n73 ) : ( n2544 ) ;
assign n2546 =  ( n1828 ) ? ( bv_8_165_n69 ) : ( n2545 ) ;
assign n2547 =  ( n1826 ) ? ( bv_8_3_n65 ) : ( n2546 ) ;
assign n2548 =  ( n1824 ) ? ( bv_8_89_n61 ) : ( n2547 ) ;
assign n2549 =  ( n1822 ) ? ( bv_8_9_n57 ) : ( n2548 ) ;
assign n2550 =  ( n1820 ) ? ( bv_8_26_n53 ) : ( n2549 ) ;
assign n2551 =  ( n1818 ) ? ( bv_8_101_n49 ) : ( n2550 ) ;
assign n2552 =  ( n1816 ) ? ( bv_8_215_n45 ) : ( n2551 ) ;
assign n2553 =  ( n1814 ) ? ( bv_8_132_n41 ) : ( n2552 ) ;
assign n2554 =  ( n1812 ) ? ( bv_8_208_n37 ) : ( n2553 ) ;
assign n2555 =  ( n1810 ) ? ( bv_8_130_n33 ) : ( n2554 ) ;
assign n2556 =  ( n1808 ) ? ( bv_8_41_n29 ) : ( n2555 ) ;
assign n2557 =  ( n1806 ) ? ( bv_8_90_n25 ) : ( n2556 ) ;
assign n2558 =  ( n1804 ) ? ( bv_8_30_n21 ) : ( n2557 ) ;
assign n2559 =  ( n1802 ) ? ( bv_8_123_n17 ) : ( n2558 ) ;
assign n2560 =  ( n1800 ) ? ( bv_8_168_n13 ) : ( n2559 ) ;
assign n2561 =  ( n1798 ) ? ( bv_8_109_n9 ) : ( n2560 ) ;
assign n2562 =  ( n1796 ) ? ( bv_8_44_n5 ) : ( n2561 ) ;
assign n2563 =  ( n1794 ) ^ ( n2562 )  ;
assign n2564 = state_in[47:40] ;
assign n2565 =  ( n2564 ) == ( bv_8_255_n3 )  ;
assign n2566 = state_in[47:40] ;
assign n2567 =  ( n2566 ) == ( bv_8_254_n7 )  ;
assign n2568 = state_in[47:40] ;
assign n2569 =  ( n2568 ) == ( bv_8_253_n11 )  ;
assign n2570 = state_in[47:40] ;
assign n2571 =  ( n2570 ) == ( bv_8_252_n15 )  ;
assign n2572 = state_in[47:40] ;
assign n2573 =  ( n2572 ) == ( bv_8_251_n19 )  ;
assign n2574 = state_in[47:40] ;
assign n2575 =  ( n2574 ) == ( bv_8_250_n23 )  ;
assign n2576 = state_in[47:40] ;
assign n2577 =  ( n2576 ) == ( bv_8_249_n27 )  ;
assign n2578 = state_in[47:40] ;
assign n2579 =  ( n2578 ) == ( bv_8_248_n31 )  ;
assign n2580 = state_in[47:40] ;
assign n2581 =  ( n2580 ) == ( bv_8_247_n35 )  ;
assign n2582 = state_in[47:40] ;
assign n2583 =  ( n2582 ) == ( bv_8_246_n39 )  ;
assign n2584 = state_in[47:40] ;
assign n2585 =  ( n2584 ) == ( bv_8_245_n43 )  ;
assign n2586 = state_in[47:40] ;
assign n2587 =  ( n2586 ) == ( bv_8_244_n47 )  ;
assign n2588 = state_in[47:40] ;
assign n2589 =  ( n2588 ) == ( bv_8_243_n51 )  ;
assign n2590 = state_in[47:40] ;
assign n2591 =  ( n2590 ) == ( bv_8_242_n55 )  ;
assign n2592 = state_in[47:40] ;
assign n2593 =  ( n2592 ) == ( bv_8_241_n59 )  ;
assign n2594 = state_in[47:40] ;
assign n2595 =  ( n2594 ) == ( bv_8_240_n63 )  ;
assign n2596 = state_in[47:40] ;
assign n2597 =  ( n2596 ) == ( bv_8_239_n67 )  ;
assign n2598 = state_in[47:40] ;
assign n2599 =  ( n2598 ) == ( bv_8_238_n71 )  ;
assign n2600 = state_in[47:40] ;
assign n2601 =  ( n2600 ) == ( bv_8_237_n75 )  ;
assign n2602 = state_in[47:40] ;
assign n2603 =  ( n2602 ) == ( bv_8_236_n79 )  ;
assign n2604 = state_in[47:40] ;
assign n2605 =  ( n2604 ) == ( bv_8_235_n83 )  ;
assign n2606 = state_in[47:40] ;
assign n2607 =  ( n2606 ) == ( bv_8_234_n87 )  ;
assign n2608 = state_in[47:40] ;
assign n2609 =  ( n2608 ) == ( bv_8_233_n91 )  ;
assign n2610 = state_in[47:40] ;
assign n2611 =  ( n2610 ) == ( bv_8_232_n95 )  ;
assign n2612 = state_in[47:40] ;
assign n2613 =  ( n2612 ) == ( bv_8_231_n99 )  ;
assign n2614 = state_in[47:40] ;
assign n2615 =  ( n2614 ) == ( bv_8_230_n103 )  ;
assign n2616 = state_in[47:40] ;
assign n2617 =  ( n2616 ) == ( bv_8_229_n107 )  ;
assign n2618 = state_in[47:40] ;
assign n2619 =  ( n2618 ) == ( bv_8_228_n111 )  ;
assign n2620 = state_in[47:40] ;
assign n2621 =  ( n2620 ) == ( bv_8_227_n115 )  ;
assign n2622 = state_in[47:40] ;
assign n2623 =  ( n2622 ) == ( bv_8_226_n119 )  ;
assign n2624 = state_in[47:40] ;
assign n2625 =  ( n2624 ) == ( bv_8_225_n123 )  ;
assign n2626 = state_in[47:40] ;
assign n2627 =  ( n2626 ) == ( bv_8_224_n126 )  ;
assign n2628 = state_in[47:40] ;
assign n2629 =  ( n2628 ) == ( bv_8_223_n130 )  ;
assign n2630 = state_in[47:40] ;
assign n2631 =  ( n2630 ) == ( bv_8_222_n134 )  ;
assign n2632 = state_in[47:40] ;
assign n2633 =  ( n2632 ) == ( bv_8_221_n138 )  ;
assign n2634 = state_in[47:40] ;
assign n2635 =  ( n2634 ) == ( bv_8_220_n142 )  ;
assign n2636 = state_in[47:40] ;
assign n2637 =  ( n2636 ) == ( bv_8_219_n146 )  ;
assign n2638 = state_in[47:40] ;
assign n2639 =  ( n2638 ) == ( bv_8_218_n150 )  ;
assign n2640 = state_in[47:40] ;
assign n2641 =  ( n2640 ) == ( bv_8_217_n128 )  ;
assign n2642 = state_in[47:40] ;
assign n2643 =  ( n2642 ) == ( bv_8_216_n157 )  ;
assign n2644 = state_in[47:40] ;
assign n2645 =  ( n2644 ) == ( bv_8_215_n45 )  ;
assign n2646 = state_in[47:40] ;
assign n2647 =  ( n2646 ) == ( bv_8_214_n164 )  ;
assign n2648 = state_in[47:40] ;
assign n2649 =  ( n2648 ) == ( bv_8_213_n167 )  ;
assign n2650 = state_in[47:40] ;
assign n2651 =  ( n2650 ) == ( bv_8_212_n171 )  ;
assign n2652 = state_in[47:40] ;
assign n2653 =  ( n2652 ) == ( bv_8_211_n175 )  ;
assign n2654 = state_in[47:40] ;
assign n2655 =  ( n2654 ) == ( bv_8_210_n113 )  ;
assign n2656 = state_in[47:40] ;
assign n2657 =  ( n2656 ) == ( bv_8_209_n182 )  ;
assign n2658 = state_in[47:40] ;
assign n2659 =  ( n2658 ) == ( bv_8_208_n37 )  ;
assign n2660 = state_in[47:40] ;
assign n2661 =  ( n2660 ) == ( bv_8_207_n188 )  ;
assign n2662 = state_in[47:40] ;
assign n2663 =  ( n2662 ) == ( bv_8_206_n192 )  ;
assign n2664 = state_in[47:40] ;
assign n2665 =  ( n2664 ) == ( bv_8_205_n196 )  ;
assign n2666 = state_in[47:40] ;
assign n2667 =  ( n2666 ) == ( bv_8_204_n177 )  ;
assign n2668 = state_in[47:40] ;
assign n2669 =  ( n2668 ) == ( bv_8_203_n203 )  ;
assign n2670 = state_in[47:40] ;
assign n2671 =  ( n2670 ) == ( bv_8_202_n207 )  ;
assign n2672 = state_in[47:40] ;
assign n2673 =  ( n2672 ) == ( bv_8_201_n85 )  ;
assign n2674 = state_in[47:40] ;
assign n2675 =  ( n2674 ) == ( bv_8_200_n213 )  ;
assign n2676 = state_in[47:40] ;
assign n2677 =  ( n2676 ) == ( bv_8_199_n216 )  ;
assign n2678 = state_in[47:40] ;
assign n2679 =  ( n2678 ) == ( bv_8_198_n220 )  ;
assign n2680 = state_in[47:40] ;
assign n2681 =  ( n2680 ) == ( bv_8_197_n224 )  ;
assign n2682 = state_in[47:40] ;
assign n2683 =  ( n2682 ) == ( bv_8_196_n228 )  ;
assign n2684 = state_in[47:40] ;
assign n2685 =  ( n2684 ) == ( bv_8_195_n232 )  ;
assign n2686 = state_in[47:40] ;
assign n2687 =  ( n2686 ) == ( bv_8_194_n159 )  ;
assign n2688 = state_in[47:40] ;
assign n2689 =  ( n2688 ) == ( bv_8_193_n239 )  ;
assign n2690 = state_in[47:40] ;
assign n2691 =  ( n2690 ) == ( bv_8_192_n242 )  ;
assign n2692 = state_in[47:40] ;
assign n2693 =  ( n2692 ) == ( bv_8_191_n246 )  ;
assign n2694 = state_in[47:40] ;
assign n2695 =  ( n2694 ) == ( bv_8_190_n250 )  ;
assign n2696 = state_in[47:40] ;
assign n2697 =  ( n2696 ) == ( bv_8_189_n254 )  ;
assign n2698 = state_in[47:40] ;
assign n2699 =  ( n2698 ) == ( bv_8_188_n257 )  ;
assign n2700 = state_in[47:40] ;
assign n2701 =  ( n2700 ) == ( bv_8_187_n260 )  ;
assign n2702 = state_in[47:40] ;
assign n2703 =  ( n2702 ) == ( bv_8_186_n263 )  ;
assign n2704 = state_in[47:40] ;
assign n2705 =  ( n2704 ) == ( bv_8_185_n266 )  ;
assign n2706 = state_in[47:40] ;
assign n2707 =  ( n2706 ) == ( bv_8_184_n270 )  ;
assign n2708 = state_in[47:40] ;
assign n2709 =  ( n2708 ) == ( bv_8_183_n273 )  ;
assign n2710 = state_in[47:40] ;
assign n2711 =  ( n2710 ) == ( bv_8_182_n277 )  ;
assign n2712 = state_in[47:40] ;
assign n2713 =  ( n2712 ) == ( bv_8_181_n281 )  ;
assign n2714 = state_in[47:40] ;
assign n2715 =  ( n2714 ) == ( bv_8_180_n285 )  ;
assign n2716 = state_in[47:40] ;
assign n2717 =  ( n2716 ) == ( bv_8_179_n289 )  ;
assign n2718 = state_in[47:40] ;
assign n2719 =  ( n2718 ) == ( bv_8_178_n292 )  ;
assign n2720 = state_in[47:40] ;
assign n2721 =  ( n2720 ) == ( bv_8_177_n283 )  ;
assign n2722 = state_in[47:40] ;
assign n2723 =  ( n2722 ) == ( bv_8_176_n299 )  ;
assign n2724 = state_in[47:40] ;
assign n2725 =  ( n2724 ) == ( bv_8_175_n302 )  ;
assign n2726 = state_in[47:40] ;
assign n2727 =  ( n2726 ) == ( bv_8_174_n152 )  ;
assign n2728 = state_in[47:40] ;
assign n2729 =  ( n2728 ) == ( bv_8_173_n307 )  ;
assign n2730 = state_in[47:40] ;
assign n2731 =  ( n2730 ) == ( bv_8_172_n268 )  ;
assign n2732 = state_in[47:40] ;
assign n2733 =  ( n2732 ) == ( bv_8_171_n314 )  ;
assign n2734 = state_in[47:40] ;
assign n2735 =  ( n2734 ) == ( bv_8_170_n77 )  ;
assign n2736 = state_in[47:40] ;
assign n2737 =  ( n2736 ) == ( bv_8_169_n109 )  ;
assign n2738 = state_in[47:40] ;
assign n2739 =  ( n2738 ) == ( bv_8_168_n13 )  ;
assign n2740 = state_in[47:40] ;
assign n2741 =  ( n2740 ) == ( bv_8_167_n325 )  ;
assign n2742 = state_in[47:40] ;
assign n2743 =  ( n2742 ) == ( bv_8_166_n328 )  ;
assign n2744 = state_in[47:40] ;
assign n2745 =  ( n2744 ) == ( bv_8_165_n69 )  ;
assign n2746 = state_in[47:40] ;
assign n2747 =  ( n2746 ) == ( bv_8_164_n335 )  ;
assign n2748 = state_in[47:40] ;
assign n2749 =  ( n2748 ) == ( bv_8_163_n339 )  ;
assign n2750 = state_in[47:40] ;
assign n2751 =  ( n2750 ) == ( bv_8_162_n343 )  ;
assign n2752 = state_in[47:40] ;
assign n2753 =  ( n2752 ) == ( bv_8_161_n211 )  ;
assign n2754 = state_in[47:40] ;
assign n2755 =  ( n2754 ) == ( bv_8_160_n350 )  ;
assign n2756 = state_in[47:40] ;
assign n2757 =  ( n2756 ) == ( bv_8_159_n323 )  ;
assign n2758 = state_in[47:40] ;
assign n2759 =  ( n2758 ) == ( bv_8_158_n355 )  ;
assign n2760 = state_in[47:40] ;
assign n2761 =  ( n2760 ) == ( bv_8_157_n359 )  ;
assign n2762 = state_in[47:40] ;
assign n2763 =  ( n2762 ) == ( bv_8_156_n279 )  ;
assign n2764 = state_in[47:40] ;
assign n2765 =  ( n2764 ) == ( bv_8_155_n364 )  ;
assign n2766 = state_in[47:40] ;
assign n2767 =  ( n2766 ) == ( bv_8_154_n368 )  ;
assign n2768 = state_in[47:40] ;
assign n2769 =  ( n2768 ) == ( bv_8_153_n140 )  ;
assign n2770 = state_in[47:40] ;
assign n2771 =  ( n2770 ) == ( bv_8_152_n374 )  ;
assign n2772 = state_in[47:40] ;
assign n2773 =  ( n2772 ) == ( bv_8_151_n218 )  ;
assign n2774 = state_in[47:40] ;
assign n2775 =  ( n2774 ) == ( bv_8_150_n201 )  ;
assign n2776 = state_in[47:40] ;
assign n2777 =  ( n2776 ) == ( bv_8_149_n384 )  ;
assign n2778 = state_in[47:40] ;
assign n2779 =  ( n2778 ) == ( bv_8_148_n388 )  ;
assign n2780 = state_in[47:40] ;
assign n2781 =  ( n2780 ) == ( bv_8_147_n392 )  ;
assign n2782 = state_in[47:40] ;
assign n2783 =  ( n2782 ) == ( bv_8_146_n337 )  ;
assign n2784 = state_in[47:40] ;
assign n2785 =  ( n2784 ) == ( bv_8_145_n397 )  ;
assign n2786 = state_in[47:40] ;
assign n2787 =  ( n2786 ) == ( bv_8_144_n173 )  ;
assign n2788 = state_in[47:40] ;
assign n2789 =  ( n2788 ) == ( bv_8_143_n403 )  ;
assign n2790 = state_in[47:40] ;
assign n2791 =  ( n2790 ) == ( bv_8_142_n406 )  ;
assign n2792 = state_in[47:40] ;
assign n2793 =  ( n2792 ) == ( bv_8_141_n410 )  ;
assign n2794 = state_in[47:40] ;
assign n2795 =  ( n2794 ) == ( bv_8_140_n376 )  ;
assign n2796 = state_in[47:40] ;
assign n2797 =  ( n2796 ) == ( bv_8_139_n297 )  ;
assign n2798 = state_in[47:40] ;
assign n2799 =  ( n2798 ) == ( bv_8_138_n418 )  ;
assign n2800 = state_in[47:40] ;
assign n2801 =  ( n2800 ) == ( bv_8_137_n421 )  ;
assign n2802 = state_in[47:40] ;
assign n2803 =  ( n2802 ) == ( bv_8_136_n425 )  ;
assign n2804 = state_in[47:40] ;
assign n2805 =  ( n2804 ) == ( bv_8_135_n81 )  ;
assign n2806 = state_in[47:40] ;
assign n2807 =  ( n2806 ) == ( bv_8_134_n431 )  ;
assign n2808 = state_in[47:40] ;
assign n2809 =  ( n2808 ) == ( bv_8_133_n434 )  ;
assign n2810 = state_in[47:40] ;
assign n2811 =  ( n2810 ) == ( bv_8_132_n41 )  ;
assign n2812 = state_in[47:40] ;
assign n2813 =  ( n2812 ) == ( bv_8_131_n440 )  ;
assign n2814 = state_in[47:40] ;
assign n2815 =  ( n2814 ) == ( bv_8_130_n33 )  ;
assign n2816 = state_in[47:40] ;
assign n2817 =  ( n2816 ) == ( bv_8_129_n446 )  ;
assign n2818 = state_in[47:40] ;
assign n2819 =  ( n2818 ) == ( bv_8_128_n450 )  ;
assign n2820 = state_in[47:40] ;
assign n2821 =  ( n2820 ) == ( bv_8_127_n453 )  ;
assign n2822 = state_in[47:40] ;
assign n2823 =  ( n2822 ) == ( bv_8_126_n456 )  ;
assign n2824 = state_in[47:40] ;
assign n2825 =  ( n2824 ) == ( bv_8_125_n459 )  ;
assign n2826 = state_in[47:40] ;
assign n2827 =  ( n2826 ) == ( bv_8_124_n184 )  ;
assign n2828 = state_in[47:40] ;
assign n2829 =  ( n2828 ) == ( bv_8_123_n17 )  ;
assign n2830 = state_in[47:40] ;
assign n2831 =  ( n2830 ) == ( bv_8_122_n416 )  ;
assign n2832 = state_in[47:40] ;
assign n2833 =  ( n2832 ) == ( bv_8_121_n470 )  ;
assign n2834 = state_in[47:40] ;
assign n2835 =  ( n2834 ) == ( bv_8_120_n474 )  ;
assign n2836 = state_in[47:40] ;
assign n2837 =  ( n2836 ) == ( bv_8_119_n472 )  ;
assign n2838 = state_in[47:40] ;
assign n2839 =  ( n2838 ) == ( bv_8_118_n480 )  ;
assign n2840 = state_in[47:40] ;
assign n2841 =  ( n2840 ) == ( bv_8_117_n484 )  ;
assign n2842 = state_in[47:40] ;
assign n2843 =  ( n2842 ) == ( bv_8_116_n345 )  ;
assign n2844 = state_in[47:40] ;
assign n2845 =  ( n2844 ) == ( bv_8_115_n222 )  ;
assign n2846 = state_in[47:40] ;
assign n2847 =  ( n2846 ) == ( bv_8_114_n494 )  ;
assign n2848 = state_in[47:40] ;
assign n2849 =  ( n2848 ) == ( bv_8_113_n180 )  ;
assign n2850 = state_in[47:40] ;
assign n2851 =  ( n2850 ) == ( bv_8_112_n482 )  ;
assign n2852 = state_in[47:40] ;
assign n2853 =  ( n2852 ) == ( bv_8_111_n244 )  ;
assign n2854 = state_in[47:40] ;
assign n2855 =  ( n2854 ) == ( bv_8_110_n294 )  ;
assign n2856 = state_in[47:40] ;
assign n2857 =  ( n2856 ) == ( bv_8_109_n9 )  ;
assign n2858 = state_in[47:40] ;
assign n2859 =  ( n2858 ) == ( bv_8_108_n510 )  ;
assign n2860 = state_in[47:40] ;
assign n2861 =  ( n2860 ) == ( bv_8_107_n370 )  ;
assign n2862 = state_in[47:40] ;
assign n2863 =  ( n2862 ) == ( bv_8_106_n155 )  ;
assign n2864 = state_in[47:40] ;
assign n2865 =  ( n2864 ) == ( bv_8_105_n148 )  ;
assign n2866 = state_in[47:40] ;
assign n2867 =  ( n2866 ) == ( bv_8_104_n520 )  ;
assign n2868 = state_in[47:40] ;
assign n2869 =  ( n2868 ) == ( bv_8_103_n523 )  ;
assign n2870 = state_in[47:40] ;
assign n2871 =  ( n2870 ) == ( bv_8_102_n527 )  ;
assign n2872 = state_in[47:40] ;
assign n2873 =  ( n2872 ) == ( bv_8_101_n49 )  ;
assign n2874 = state_in[47:40] ;
assign n2875 =  ( n2874 ) == ( bv_8_100_n348 )  ;
assign n2876 = state_in[47:40] ;
assign n2877 =  ( n2876 ) == ( bv_8_99_n476 )  ;
assign n2878 = state_in[47:40] ;
assign n2879 =  ( n2878 ) == ( bv_8_98_n536 )  ;
assign n2880 = state_in[47:40] ;
assign n2881 =  ( n2880 ) == ( bv_8_97_n198 )  ;
assign n2882 = state_in[47:40] ;
assign n2883 =  ( n2882 ) == ( bv_8_96_n542 )  ;
assign n2884 = state_in[47:40] ;
assign n2885 =  ( n2884 ) == ( bv_8_95_n545 )  ;
assign n2886 = state_in[47:40] ;
assign n2887 =  ( n2886 ) == ( bv_8_94_n548 )  ;
assign n2888 = state_in[47:40] ;
assign n2889 =  ( n2888 ) == ( bv_8_93_n498 )  ;
assign n2890 = state_in[47:40] ;
assign n2891 =  ( n2890 ) == ( bv_8_92_n234 )  ;
assign n2892 = state_in[47:40] ;
assign n2893 =  ( n2892 ) == ( bv_8_91_n555 )  ;
assign n2894 = state_in[47:40] ;
assign n2895 =  ( n2894 ) == ( bv_8_90_n25 )  ;
assign n2896 = state_in[47:40] ;
assign n2897 =  ( n2896 ) == ( bv_8_89_n61 )  ;
assign n2898 = state_in[47:40] ;
assign n2899 =  ( n2898 ) == ( bv_8_88_n562 )  ;
assign n2900 = state_in[47:40] ;
assign n2901 =  ( n2900 ) == ( bv_8_87_n226 )  ;
assign n2902 = state_in[47:40] ;
assign n2903 =  ( n2902 ) == ( bv_8_86_n567 )  ;
assign n2904 = state_in[47:40] ;
assign n2905 =  ( n2904 ) == ( bv_8_85_n423 )  ;
assign n2906 = state_in[47:40] ;
assign n2907 =  ( n2906 ) == ( bv_8_84_n386 )  ;
assign n2908 = state_in[47:40] ;
assign n2909 =  ( n2908 ) == ( bv_8_83_n575 )  ;
assign n2910 = state_in[47:40] ;
assign n2911 =  ( n2910 ) == ( bv_8_82_n578 )  ;
assign n2912 = state_in[47:40] ;
assign n2913 =  ( n2912 ) == ( bv_8_81_n582 )  ;
assign n2914 = state_in[47:40] ;
assign n2915 =  ( n2914 ) == ( bv_8_80_n73 )  ;
assign n2916 = state_in[47:40] ;
assign n2917 =  ( n2916 ) == ( bv_8_79_n538 )  ;
assign n2918 = state_in[47:40] ;
assign n2919 =  ( n2918 ) == ( bv_8_78_n590 )  ;
assign n2920 = state_in[47:40] ;
assign n2921 =  ( n2920 ) == ( bv_8_77_n593 )  ;
assign n2922 = state_in[47:40] ;
assign n2923 =  ( n2922 ) == ( bv_8_76_n596 )  ;
assign n2924 = state_in[47:40] ;
assign n2925 =  ( n2924 ) == ( bv_8_75_n503 )  ;
assign n2926 = state_in[47:40] ;
assign n2927 =  ( n2926 ) == ( bv_8_74_n237 )  ;
assign n2928 = state_in[47:40] ;
assign n2929 =  ( n2928 ) == ( bv_8_73_n275 )  ;
assign n2930 = state_in[47:40] ;
assign n2931 =  ( n2930 ) == ( bv_8_72_n330 )  ;
assign n2932 = state_in[47:40] ;
assign n2933 =  ( n2932 ) == ( bv_8_71_n252 )  ;
assign n2934 = state_in[47:40] ;
assign n2935 =  ( n2934 ) == ( bv_8_70_n609 )  ;
assign n2936 = state_in[47:40] ;
assign n2937 =  ( n2936 ) == ( bv_8_69_n612 )  ;
assign n2938 = state_in[47:40] ;
assign n2939 =  ( n2938 ) == ( bv_8_68_n390 )  ;
assign n2940 = state_in[47:40] ;
assign n2941 =  ( n2940 ) == ( bv_8_67_n318 )  ;
assign n2942 = state_in[47:40] ;
assign n2943 =  ( n2942 ) == ( bv_8_66_n466 )  ;
assign n2944 = state_in[47:40] ;
assign n2945 =  ( n2944 ) == ( bv_8_65_n623 )  ;
assign n2946 = state_in[47:40] ;
assign n2947 =  ( n2946 ) == ( bv_8_64_n573 )  ;
assign n2948 = state_in[47:40] ;
assign n2949 =  ( n2948 ) == ( bv_8_63_n489 )  ;
assign n2950 = state_in[47:40] ;
assign n2951 =  ( n2950 ) == ( bv_8_62_n205 )  ;
assign n2952 = state_in[47:40] ;
assign n2953 =  ( n2952 ) == ( bv_8_61_n634 )  ;
assign n2954 = state_in[47:40] ;
assign n2955 =  ( n2954 ) == ( bv_8_60_n93 )  ;
assign n2956 = state_in[47:40] ;
assign n2957 =  ( n2956 ) == ( bv_8_59_n382 )  ;
assign n2958 = state_in[47:40] ;
assign n2959 =  ( n2958 ) == ( bv_8_58_n136 )  ;
assign n2960 = state_in[47:40] ;
assign n2961 =  ( n2960 ) == ( bv_8_57_n312 )  ;
assign n2962 = state_in[47:40] ;
assign n2963 =  ( n2962 ) == ( bv_8_56_n230 )  ;
assign n2964 = state_in[47:40] ;
assign n2965 =  ( n2964 ) == ( bv_8_55_n650 )  ;
assign n2966 = state_in[47:40] ;
assign n2967 =  ( n2966 ) == ( bv_8_54_n616 )  ;
assign n2968 = state_in[47:40] ;
assign n2969 =  ( n2968 ) == ( bv_8_53_n436 )  ;
assign n2970 = state_in[47:40] ;
assign n2971 =  ( n2970 ) == ( bv_8_52_n619 )  ;
assign n2972 = state_in[47:40] ;
assign n2973 =  ( n2972 ) == ( bv_8_51_n101 )  ;
assign n2974 = state_in[47:40] ;
assign n2975 =  ( n2974 ) == ( bv_8_50_n408 )  ;
assign n2976 = state_in[47:40] ;
assign n2977 =  ( n2976 ) == ( bv_8_49_n309 )  ;
assign n2978 = state_in[47:40] ;
assign n2979 =  ( n2978 ) == ( bv_8_48_n660 )  ;
assign n2980 = state_in[47:40] ;
assign n2981 =  ( n2980 ) == ( bv_8_47_n652 )  ;
assign n2982 = state_in[47:40] ;
assign n2983 =  ( n2982 ) == ( bv_8_46_n429 )  ;
assign n2984 = state_in[47:40] ;
assign n2985 =  ( n2984 ) == ( bv_8_45_n97 )  ;
assign n2986 = state_in[47:40] ;
assign n2987 =  ( n2986 ) == ( bv_8_44_n5 )  ;
assign n2988 = state_in[47:40] ;
assign n2989 =  ( n2988 ) == ( bv_8_43_n121 )  ;
assign n2990 = state_in[47:40] ;
assign n2991 =  ( n2990 ) == ( bv_8_42_n672 )  ;
assign n2992 = state_in[47:40] ;
assign n2993 =  ( n2992 ) == ( bv_8_41_n29 )  ;
assign n2994 = state_in[47:40] ;
assign n2995 =  ( n2994 ) == ( bv_8_40_n366 )  ;
assign n2996 = state_in[47:40] ;
assign n2997 =  ( n2996 ) == ( bv_8_39_n132 )  ;
assign n2998 = state_in[47:40] ;
assign n2999 =  ( n2998 ) == ( bv_8_38_n444 )  ;
assign n3000 = state_in[47:40] ;
assign n3001 =  ( n3000 ) == ( bv_8_37_n506 )  ;
assign n3002 = state_in[47:40] ;
assign n3003 =  ( n3002 ) == ( bv_8_36_n645 )  ;
assign n3004 = state_in[47:40] ;
assign n3005 =  ( n3004 ) == ( bv_8_35_n696 )  ;
assign n3006 = state_in[47:40] ;
assign n3007 =  ( n3006 ) == ( bv_8_34_n117 )  ;
assign n3008 = state_in[47:40] ;
assign n3009 =  ( n3008 ) == ( bv_8_33_n486 )  ;
assign n3010 = state_in[47:40] ;
assign n3011 =  ( n3010 ) == ( bv_8_32_n463 )  ;
assign n3012 = state_in[47:40] ;
assign n3013 =  ( n3012 ) == ( bv_8_31_n705 )  ;
assign n3014 = state_in[47:40] ;
assign n3015 =  ( n3014 ) == ( bv_8_30_n21 )  ;
assign n3016 = state_in[47:40] ;
assign n3017 =  ( n3016 ) == ( bv_8_29_n625 )  ;
assign n3018 = state_in[47:40] ;
assign n3019 =  ( n3018 ) == ( bv_8_28_n162 )  ;
assign n3020 = state_in[47:40] ;
assign n3021 =  ( n3020 ) == ( bv_8_27_n642 )  ;
assign n3022 = state_in[47:40] ;
assign n3023 =  ( n3022 ) == ( bv_8_26_n53 )  ;
assign n3024 = state_in[47:40] ;
assign n3025 =  ( n3024 ) == ( bv_8_25_n399 )  ;
assign n3026 = state_in[47:40] ;
assign n3027 =  ( n3026 ) == ( bv_8_24_n448 )  ;
assign n3028 = state_in[47:40] ;
assign n3029 =  ( n3028 ) == ( bv_8_23_n144 )  ;
assign n3030 = state_in[47:40] ;
assign n3031 =  ( n3030 ) == ( bv_8_22_n357 )  ;
assign n3032 = state_in[47:40] ;
assign n3033 =  ( n3032 ) == ( bv_8_21_n89 )  ;
assign n3034 = state_in[47:40] ;
assign n3035 =  ( n3034 ) == ( bv_8_20_n341 )  ;
assign n3036 = state_in[47:40] ;
assign n3037 =  ( n3036 ) == ( bv_8_19_n588 )  ;
assign n3038 = state_in[47:40] ;
assign n3039 =  ( n3038 ) == ( bv_8_18_n628 )  ;
assign n3040 = state_in[47:40] ;
assign n3041 =  ( n3040 ) == ( bv_8_17_n525 )  ;
assign n3042 = state_in[47:40] ;
assign n3043 =  ( n3042 ) == ( bv_8_16_n248 )  ;
assign n3044 = state_in[47:40] ;
assign n3045 =  ( n3044 ) == ( bv_8_15_n190 )  ;
assign n3046 = state_in[47:40] ;
assign n3047 =  ( n3046 ) == ( bv_8_14_n648 )  ;
assign n3048 = state_in[47:40] ;
assign n3049 =  ( n3048 ) == ( bv_8_13_n194 )  ;
assign n3050 = state_in[47:40] ;
assign n3051 =  ( n3050 ) == ( bv_8_12_n333 )  ;
assign n3052 = state_in[47:40] ;
assign n3053 =  ( n3052 ) == ( bv_8_11_n379 )  ;
assign n3054 = state_in[47:40] ;
assign n3055 =  ( n3054 ) == ( bv_8_10_n655 )  ;
assign n3056 = state_in[47:40] ;
assign n3057 =  ( n3056 ) == ( bv_8_9_n57 )  ;
assign n3058 = state_in[47:40] ;
assign n3059 =  ( n3058 ) == ( bv_8_8_n669 )  ;
assign n3060 = state_in[47:40] ;
assign n3061 =  ( n3060 ) == ( bv_8_7_n105 )  ;
assign n3062 = state_in[47:40] ;
assign n3063 =  ( n3062 ) == ( bv_8_6_n169 )  ;
assign n3064 = state_in[47:40] ;
assign n3065 =  ( n3064 ) == ( bv_8_5_n492 )  ;
assign n3066 = state_in[47:40] ;
assign n3067 =  ( n3066 ) == ( bv_8_4_n516 )  ;
assign n3068 = state_in[47:40] ;
assign n3069 =  ( n3068 ) == ( bv_8_3_n65 )  ;
assign n3070 = state_in[47:40] ;
assign n3071 =  ( n3070 ) == ( bv_8_2_n751 )  ;
assign n3072 = state_in[47:40] ;
assign n3073 =  ( n3072 ) == ( bv_8_1_n287 )  ;
assign n3074 = state_in[47:40] ;
assign n3075 =  ( n3074 ) == ( bv_8_0_n580 )  ;
assign n3076 =  ( n3075 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n3077 =  ( n3073 ) ? ( bv_8_124_n184 ) : ( n3076 ) ;
assign n3078 =  ( n3071 ) ? ( bv_8_119_n472 ) : ( n3077 ) ;
assign n3079 =  ( n3069 ) ? ( bv_8_123_n17 ) : ( n3078 ) ;
assign n3080 =  ( n3067 ) ? ( bv_8_242_n55 ) : ( n3079 ) ;
assign n3081 =  ( n3065 ) ? ( bv_8_107_n370 ) : ( n3080 ) ;
assign n3082 =  ( n3063 ) ? ( bv_8_111_n244 ) : ( n3081 ) ;
assign n3083 =  ( n3061 ) ? ( bv_8_197_n224 ) : ( n3082 ) ;
assign n3084 =  ( n3059 ) ? ( bv_8_48_n660 ) : ( n3083 ) ;
assign n3085 =  ( n3057 ) ? ( bv_8_1_n287 ) : ( n3084 ) ;
assign n3086 =  ( n3055 ) ? ( bv_8_103_n523 ) : ( n3085 ) ;
assign n3087 =  ( n3053 ) ? ( bv_8_43_n121 ) : ( n3086 ) ;
assign n3088 =  ( n3051 ) ? ( bv_8_254_n7 ) : ( n3087 ) ;
assign n3089 =  ( n3049 ) ? ( bv_8_215_n45 ) : ( n3088 ) ;
assign n3090 =  ( n3047 ) ? ( bv_8_171_n314 ) : ( n3089 ) ;
assign n3091 =  ( n3045 ) ? ( bv_8_118_n480 ) : ( n3090 ) ;
assign n3092 =  ( n3043 ) ? ( bv_8_202_n207 ) : ( n3091 ) ;
assign n3093 =  ( n3041 ) ? ( bv_8_130_n33 ) : ( n3092 ) ;
assign n3094 =  ( n3039 ) ? ( bv_8_201_n85 ) : ( n3093 ) ;
assign n3095 =  ( n3037 ) ? ( bv_8_125_n459 ) : ( n3094 ) ;
assign n3096 =  ( n3035 ) ? ( bv_8_250_n23 ) : ( n3095 ) ;
assign n3097 =  ( n3033 ) ? ( bv_8_89_n61 ) : ( n3096 ) ;
assign n3098 =  ( n3031 ) ? ( bv_8_71_n252 ) : ( n3097 ) ;
assign n3099 =  ( n3029 ) ? ( bv_8_240_n63 ) : ( n3098 ) ;
assign n3100 =  ( n3027 ) ? ( bv_8_173_n307 ) : ( n3099 ) ;
assign n3101 =  ( n3025 ) ? ( bv_8_212_n171 ) : ( n3100 ) ;
assign n3102 =  ( n3023 ) ? ( bv_8_162_n343 ) : ( n3101 ) ;
assign n3103 =  ( n3021 ) ? ( bv_8_175_n302 ) : ( n3102 ) ;
assign n3104 =  ( n3019 ) ? ( bv_8_156_n279 ) : ( n3103 ) ;
assign n3105 =  ( n3017 ) ? ( bv_8_164_n335 ) : ( n3104 ) ;
assign n3106 =  ( n3015 ) ? ( bv_8_114_n494 ) : ( n3105 ) ;
assign n3107 =  ( n3013 ) ? ( bv_8_192_n242 ) : ( n3106 ) ;
assign n3108 =  ( n3011 ) ? ( bv_8_183_n273 ) : ( n3107 ) ;
assign n3109 =  ( n3009 ) ? ( bv_8_253_n11 ) : ( n3108 ) ;
assign n3110 =  ( n3007 ) ? ( bv_8_147_n392 ) : ( n3109 ) ;
assign n3111 =  ( n3005 ) ? ( bv_8_38_n444 ) : ( n3110 ) ;
assign n3112 =  ( n3003 ) ? ( bv_8_54_n616 ) : ( n3111 ) ;
assign n3113 =  ( n3001 ) ? ( bv_8_63_n489 ) : ( n3112 ) ;
assign n3114 =  ( n2999 ) ? ( bv_8_247_n35 ) : ( n3113 ) ;
assign n3115 =  ( n2997 ) ? ( bv_8_204_n177 ) : ( n3114 ) ;
assign n3116 =  ( n2995 ) ? ( bv_8_52_n619 ) : ( n3115 ) ;
assign n3117 =  ( n2993 ) ? ( bv_8_165_n69 ) : ( n3116 ) ;
assign n3118 =  ( n2991 ) ? ( bv_8_229_n107 ) : ( n3117 ) ;
assign n3119 =  ( n2989 ) ? ( bv_8_241_n59 ) : ( n3118 ) ;
assign n3120 =  ( n2987 ) ? ( bv_8_113_n180 ) : ( n3119 ) ;
assign n3121 =  ( n2985 ) ? ( bv_8_216_n157 ) : ( n3120 ) ;
assign n3122 =  ( n2983 ) ? ( bv_8_49_n309 ) : ( n3121 ) ;
assign n3123 =  ( n2981 ) ? ( bv_8_21_n89 ) : ( n3122 ) ;
assign n3124 =  ( n2979 ) ? ( bv_8_4_n516 ) : ( n3123 ) ;
assign n3125 =  ( n2977 ) ? ( bv_8_199_n216 ) : ( n3124 ) ;
assign n3126 =  ( n2975 ) ? ( bv_8_35_n696 ) : ( n3125 ) ;
assign n3127 =  ( n2973 ) ? ( bv_8_195_n232 ) : ( n3126 ) ;
assign n3128 =  ( n2971 ) ? ( bv_8_24_n448 ) : ( n3127 ) ;
assign n3129 =  ( n2969 ) ? ( bv_8_150_n201 ) : ( n3128 ) ;
assign n3130 =  ( n2967 ) ? ( bv_8_5_n492 ) : ( n3129 ) ;
assign n3131 =  ( n2965 ) ? ( bv_8_154_n368 ) : ( n3130 ) ;
assign n3132 =  ( n2963 ) ? ( bv_8_7_n105 ) : ( n3131 ) ;
assign n3133 =  ( n2961 ) ? ( bv_8_18_n628 ) : ( n3132 ) ;
assign n3134 =  ( n2959 ) ? ( bv_8_128_n450 ) : ( n3133 ) ;
assign n3135 =  ( n2957 ) ? ( bv_8_226_n119 ) : ( n3134 ) ;
assign n3136 =  ( n2955 ) ? ( bv_8_235_n83 ) : ( n3135 ) ;
assign n3137 =  ( n2953 ) ? ( bv_8_39_n132 ) : ( n3136 ) ;
assign n3138 =  ( n2951 ) ? ( bv_8_178_n292 ) : ( n3137 ) ;
assign n3139 =  ( n2949 ) ? ( bv_8_117_n484 ) : ( n3138 ) ;
assign n3140 =  ( n2947 ) ? ( bv_8_9_n57 ) : ( n3139 ) ;
assign n3141 =  ( n2945 ) ? ( bv_8_131_n440 ) : ( n3140 ) ;
assign n3142 =  ( n2943 ) ? ( bv_8_44_n5 ) : ( n3141 ) ;
assign n3143 =  ( n2941 ) ? ( bv_8_26_n53 ) : ( n3142 ) ;
assign n3144 =  ( n2939 ) ? ( bv_8_27_n642 ) : ( n3143 ) ;
assign n3145 =  ( n2937 ) ? ( bv_8_110_n294 ) : ( n3144 ) ;
assign n3146 =  ( n2935 ) ? ( bv_8_90_n25 ) : ( n3145 ) ;
assign n3147 =  ( n2933 ) ? ( bv_8_160_n350 ) : ( n3146 ) ;
assign n3148 =  ( n2931 ) ? ( bv_8_82_n578 ) : ( n3147 ) ;
assign n3149 =  ( n2929 ) ? ( bv_8_59_n382 ) : ( n3148 ) ;
assign n3150 =  ( n2927 ) ? ( bv_8_214_n164 ) : ( n3149 ) ;
assign n3151 =  ( n2925 ) ? ( bv_8_179_n289 ) : ( n3150 ) ;
assign n3152 =  ( n2923 ) ? ( bv_8_41_n29 ) : ( n3151 ) ;
assign n3153 =  ( n2921 ) ? ( bv_8_227_n115 ) : ( n3152 ) ;
assign n3154 =  ( n2919 ) ? ( bv_8_47_n652 ) : ( n3153 ) ;
assign n3155 =  ( n2917 ) ? ( bv_8_132_n41 ) : ( n3154 ) ;
assign n3156 =  ( n2915 ) ? ( bv_8_83_n575 ) : ( n3155 ) ;
assign n3157 =  ( n2913 ) ? ( bv_8_209_n182 ) : ( n3156 ) ;
assign n3158 =  ( n2911 ) ? ( bv_8_0_n580 ) : ( n3157 ) ;
assign n3159 =  ( n2909 ) ? ( bv_8_237_n75 ) : ( n3158 ) ;
assign n3160 =  ( n2907 ) ? ( bv_8_32_n463 ) : ( n3159 ) ;
assign n3161 =  ( n2905 ) ? ( bv_8_252_n15 ) : ( n3160 ) ;
assign n3162 =  ( n2903 ) ? ( bv_8_177_n283 ) : ( n3161 ) ;
assign n3163 =  ( n2901 ) ? ( bv_8_91_n555 ) : ( n3162 ) ;
assign n3164 =  ( n2899 ) ? ( bv_8_106_n155 ) : ( n3163 ) ;
assign n3165 =  ( n2897 ) ? ( bv_8_203_n203 ) : ( n3164 ) ;
assign n3166 =  ( n2895 ) ? ( bv_8_190_n250 ) : ( n3165 ) ;
assign n3167 =  ( n2893 ) ? ( bv_8_57_n312 ) : ( n3166 ) ;
assign n3168 =  ( n2891 ) ? ( bv_8_74_n237 ) : ( n3167 ) ;
assign n3169 =  ( n2889 ) ? ( bv_8_76_n596 ) : ( n3168 ) ;
assign n3170 =  ( n2887 ) ? ( bv_8_88_n562 ) : ( n3169 ) ;
assign n3171 =  ( n2885 ) ? ( bv_8_207_n188 ) : ( n3170 ) ;
assign n3172 =  ( n2883 ) ? ( bv_8_208_n37 ) : ( n3171 ) ;
assign n3173 =  ( n2881 ) ? ( bv_8_239_n67 ) : ( n3172 ) ;
assign n3174 =  ( n2879 ) ? ( bv_8_170_n77 ) : ( n3173 ) ;
assign n3175 =  ( n2877 ) ? ( bv_8_251_n19 ) : ( n3174 ) ;
assign n3176 =  ( n2875 ) ? ( bv_8_67_n318 ) : ( n3175 ) ;
assign n3177 =  ( n2873 ) ? ( bv_8_77_n593 ) : ( n3176 ) ;
assign n3178 =  ( n2871 ) ? ( bv_8_51_n101 ) : ( n3177 ) ;
assign n3179 =  ( n2869 ) ? ( bv_8_133_n434 ) : ( n3178 ) ;
assign n3180 =  ( n2867 ) ? ( bv_8_69_n612 ) : ( n3179 ) ;
assign n3181 =  ( n2865 ) ? ( bv_8_249_n27 ) : ( n3180 ) ;
assign n3182 =  ( n2863 ) ? ( bv_8_2_n751 ) : ( n3181 ) ;
assign n3183 =  ( n2861 ) ? ( bv_8_127_n453 ) : ( n3182 ) ;
assign n3184 =  ( n2859 ) ? ( bv_8_80_n73 ) : ( n3183 ) ;
assign n3185 =  ( n2857 ) ? ( bv_8_60_n93 ) : ( n3184 ) ;
assign n3186 =  ( n2855 ) ? ( bv_8_159_n323 ) : ( n3185 ) ;
assign n3187 =  ( n2853 ) ? ( bv_8_168_n13 ) : ( n3186 ) ;
assign n3188 =  ( n2851 ) ? ( bv_8_81_n582 ) : ( n3187 ) ;
assign n3189 =  ( n2849 ) ? ( bv_8_163_n339 ) : ( n3188 ) ;
assign n3190 =  ( n2847 ) ? ( bv_8_64_n573 ) : ( n3189 ) ;
assign n3191 =  ( n2845 ) ? ( bv_8_143_n403 ) : ( n3190 ) ;
assign n3192 =  ( n2843 ) ? ( bv_8_146_n337 ) : ( n3191 ) ;
assign n3193 =  ( n2841 ) ? ( bv_8_157_n359 ) : ( n3192 ) ;
assign n3194 =  ( n2839 ) ? ( bv_8_56_n230 ) : ( n3193 ) ;
assign n3195 =  ( n2837 ) ? ( bv_8_245_n43 ) : ( n3194 ) ;
assign n3196 =  ( n2835 ) ? ( bv_8_188_n257 ) : ( n3195 ) ;
assign n3197 =  ( n2833 ) ? ( bv_8_182_n277 ) : ( n3196 ) ;
assign n3198 =  ( n2831 ) ? ( bv_8_218_n150 ) : ( n3197 ) ;
assign n3199 =  ( n2829 ) ? ( bv_8_33_n486 ) : ( n3198 ) ;
assign n3200 =  ( n2827 ) ? ( bv_8_16_n248 ) : ( n3199 ) ;
assign n3201 =  ( n2825 ) ? ( bv_8_255_n3 ) : ( n3200 ) ;
assign n3202 =  ( n2823 ) ? ( bv_8_243_n51 ) : ( n3201 ) ;
assign n3203 =  ( n2821 ) ? ( bv_8_210_n113 ) : ( n3202 ) ;
assign n3204 =  ( n2819 ) ? ( bv_8_205_n196 ) : ( n3203 ) ;
assign n3205 =  ( n2817 ) ? ( bv_8_12_n333 ) : ( n3204 ) ;
assign n3206 =  ( n2815 ) ? ( bv_8_19_n588 ) : ( n3205 ) ;
assign n3207 =  ( n2813 ) ? ( bv_8_236_n79 ) : ( n3206 ) ;
assign n3208 =  ( n2811 ) ? ( bv_8_95_n545 ) : ( n3207 ) ;
assign n3209 =  ( n2809 ) ? ( bv_8_151_n218 ) : ( n3208 ) ;
assign n3210 =  ( n2807 ) ? ( bv_8_68_n390 ) : ( n3209 ) ;
assign n3211 =  ( n2805 ) ? ( bv_8_23_n144 ) : ( n3210 ) ;
assign n3212 =  ( n2803 ) ? ( bv_8_196_n228 ) : ( n3211 ) ;
assign n3213 =  ( n2801 ) ? ( bv_8_167_n325 ) : ( n3212 ) ;
assign n3214 =  ( n2799 ) ? ( bv_8_126_n456 ) : ( n3213 ) ;
assign n3215 =  ( n2797 ) ? ( bv_8_61_n634 ) : ( n3214 ) ;
assign n3216 =  ( n2795 ) ? ( bv_8_100_n348 ) : ( n3215 ) ;
assign n3217 =  ( n2793 ) ? ( bv_8_93_n498 ) : ( n3216 ) ;
assign n3218 =  ( n2791 ) ? ( bv_8_25_n399 ) : ( n3217 ) ;
assign n3219 =  ( n2789 ) ? ( bv_8_115_n222 ) : ( n3218 ) ;
assign n3220 =  ( n2787 ) ? ( bv_8_96_n542 ) : ( n3219 ) ;
assign n3221 =  ( n2785 ) ? ( bv_8_129_n446 ) : ( n3220 ) ;
assign n3222 =  ( n2783 ) ? ( bv_8_79_n538 ) : ( n3221 ) ;
assign n3223 =  ( n2781 ) ? ( bv_8_220_n142 ) : ( n3222 ) ;
assign n3224 =  ( n2779 ) ? ( bv_8_34_n117 ) : ( n3223 ) ;
assign n3225 =  ( n2777 ) ? ( bv_8_42_n672 ) : ( n3224 ) ;
assign n3226 =  ( n2775 ) ? ( bv_8_144_n173 ) : ( n3225 ) ;
assign n3227 =  ( n2773 ) ? ( bv_8_136_n425 ) : ( n3226 ) ;
assign n3228 =  ( n2771 ) ? ( bv_8_70_n609 ) : ( n3227 ) ;
assign n3229 =  ( n2769 ) ? ( bv_8_238_n71 ) : ( n3228 ) ;
assign n3230 =  ( n2767 ) ? ( bv_8_184_n270 ) : ( n3229 ) ;
assign n3231 =  ( n2765 ) ? ( bv_8_20_n341 ) : ( n3230 ) ;
assign n3232 =  ( n2763 ) ? ( bv_8_222_n134 ) : ( n3231 ) ;
assign n3233 =  ( n2761 ) ? ( bv_8_94_n548 ) : ( n3232 ) ;
assign n3234 =  ( n2759 ) ? ( bv_8_11_n379 ) : ( n3233 ) ;
assign n3235 =  ( n2757 ) ? ( bv_8_219_n146 ) : ( n3234 ) ;
assign n3236 =  ( n2755 ) ? ( bv_8_224_n126 ) : ( n3235 ) ;
assign n3237 =  ( n2753 ) ? ( bv_8_50_n408 ) : ( n3236 ) ;
assign n3238 =  ( n2751 ) ? ( bv_8_58_n136 ) : ( n3237 ) ;
assign n3239 =  ( n2749 ) ? ( bv_8_10_n655 ) : ( n3238 ) ;
assign n3240 =  ( n2747 ) ? ( bv_8_73_n275 ) : ( n3239 ) ;
assign n3241 =  ( n2745 ) ? ( bv_8_6_n169 ) : ( n3240 ) ;
assign n3242 =  ( n2743 ) ? ( bv_8_36_n645 ) : ( n3241 ) ;
assign n3243 =  ( n2741 ) ? ( bv_8_92_n234 ) : ( n3242 ) ;
assign n3244 =  ( n2739 ) ? ( bv_8_194_n159 ) : ( n3243 ) ;
assign n3245 =  ( n2737 ) ? ( bv_8_211_n175 ) : ( n3244 ) ;
assign n3246 =  ( n2735 ) ? ( bv_8_172_n268 ) : ( n3245 ) ;
assign n3247 =  ( n2733 ) ? ( bv_8_98_n536 ) : ( n3246 ) ;
assign n3248 =  ( n2731 ) ? ( bv_8_145_n397 ) : ( n3247 ) ;
assign n3249 =  ( n2729 ) ? ( bv_8_149_n384 ) : ( n3248 ) ;
assign n3250 =  ( n2727 ) ? ( bv_8_228_n111 ) : ( n3249 ) ;
assign n3251 =  ( n2725 ) ? ( bv_8_121_n470 ) : ( n3250 ) ;
assign n3252 =  ( n2723 ) ? ( bv_8_231_n99 ) : ( n3251 ) ;
assign n3253 =  ( n2721 ) ? ( bv_8_200_n213 ) : ( n3252 ) ;
assign n3254 =  ( n2719 ) ? ( bv_8_55_n650 ) : ( n3253 ) ;
assign n3255 =  ( n2717 ) ? ( bv_8_109_n9 ) : ( n3254 ) ;
assign n3256 =  ( n2715 ) ? ( bv_8_141_n410 ) : ( n3255 ) ;
assign n3257 =  ( n2713 ) ? ( bv_8_213_n167 ) : ( n3256 ) ;
assign n3258 =  ( n2711 ) ? ( bv_8_78_n590 ) : ( n3257 ) ;
assign n3259 =  ( n2709 ) ? ( bv_8_169_n109 ) : ( n3258 ) ;
assign n3260 =  ( n2707 ) ? ( bv_8_108_n510 ) : ( n3259 ) ;
assign n3261 =  ( n2705 ) ? ( bv_8_86_n567 ) : ( n3260 ) ;
assign n3262 =  ( n2703 ) ? ( bv_8_244_n47 ) : ( n3261 ) ;
assign n3263 =  ( n2701 ) ? ( bv_8_234_n87 ) : ( n3262 ) ;
assign n3264 =  ( n2699 ) ? ( bv_8_101_n49 ) : ( n3263 ) ;
assign n3265 =  ( n2697 ) ? ( bv_8_122_n416 ) : ( n3264 ) ;
assign n3266 =  ( n2695 ) ? ( bv_8_174_n152 ) : ( n3265 ) ;
assign n3267 =  ( n2693 ) ? ( bv_8_8_n669 ) : ( n3266 ) ;
assign n3268 =  ( n2691 ) ? ( bv_8_186_n263 ) : ( n3267 ) ;
assign n3269 =  ( n2689 ) ? ( bv_8_120_n474 ) : ( n3268 ) ;
assign n3270 =  ( n2687 ) ? ( bv_8_37_n506 ) : ( n3269 ) ;
assign n3271 =  ( n2685 ) ? ( bv_8_46_n429 ) : ( n3270 ) ;
assign n3272 =  ( n2683 ) ? ( bv_8_28_n162 ) : ( n3271 ) ;
assign n3273 =  ( n2681 ) ? ( bv_8_166_n328 ) : ( n3272 ) ;
assign n3274 =  ( n2679 ) ? ( bv_8_180_n285 ) : ( n3273 ) ;
assign n3275 =  ( n2677 ) ? ( bv_8_198_n220 ) : ( n3274 ) ;
assign n3276 =  ( n2675 ) ? ( bv_8_232_n95 ) : ( n3275 ) ;
assign n3277 =  ( n2673 ) ? ( bv_8_221_n138 ) : ( n3276 ) ;
assign n3278 =  ( n2671 ) ? ( bv_8_116_n345 ) : ( n3277 ) ;
assign n3279 =  ( n2669 ) ? ( bv_8_31_n705 ) : ( n3278 ) ;
assign n3280 =  ( n2667 ) ? ( bv_8_75_n503 ) : ( n3279 ) ;
assign n3281 =  ( n2665 ) ? ( bv_8_189_n254 ) : ( n3280 ) ;
assign n3282 =  ( n2663 ) ? ( bv_8_139_n297 ) : ( n3281 ) ;
assign n3283 =  ( n2661 ) ? ( bv_8_138_n418 ) : ( n3282 ) ;
assign n3284 =  ( n2659 ) ? ( bv_8_112_n482 ) : ( n3283 ) ;
assign n3285 =  ( n2657 ) ? ( bv_8_62_n205 ) : ( n3284 ) ;
assign n3286 =  ( n2655 ) ? ( bv_8_181_n281 ) : ( n3285 ) ;
assign n3287 =  ( n2653 ) ? ( bv_8_102_n527 ) : ( n3286 ) ;
assign n3288 =  ( n2651 ) ? ( bv_8_72_n330 ) : ( n3287 ) ;
assign n3289 =  ( n2649 ) ? ( bv_8_3_n65 ) : ( n3288 ) ;
assign n3290 =  ( n2647 ) ? ( bv_8_246_n39 ) : ( n3289 ) ;
assign n3291 =  ( n2645 ) ? ( bv_8_14_n648 ) : ( n3290 ) ;
assign n3292 =  ( n2643 ) ? ( bv_8_97_n198 ) : ( n3291 ) ;
assign n3293 =  ( n2641 ) ? ( bv_8_53_n436 ) : ( n3292 ) ;
assign n3294 =  ( n2639 ) ? ( bv_8_87_n226 ) : ( n3293 ) ;
assign n3295 =  ( n2637 ) ? ( bv_8_185_n266 ) : ( n3294 ) ;
assign n3296 =  ( n2635 ) ? ( bv_8_134_n431 ) : ( n3295 ) ;
assign n3297 =  ( n2633 ) ? ( bv_8_193_n239 ) : ( n3296 ) ;
assign n3298 =  ( n2631 ) ? ( bv_8_29_n625 ) : ( n3297 ) ;
assign n3299 =  ( n2629 ) ? ( bv_8_158_n355 ) : ( n3298 ) ;
assign n3300 =  ( n2627 ) ? ( bv_8_225_n123 ) : ( n3299 ) ;
assign n3301 =  ( n2625 ) ? ( bv_8_248_n31 ) : ( n3300 ) ;
assign n3302 =  ( n2623 ) ? ( bv_8_152_n374 ) : ( n3301 ) ;
assign n3303 =  ( n2621 ) ? ( bv_8_17_n525 ) : ( n3302 ) ;
assign n3304 =  ( n2619 ) ? ( bv_8_105_n148 ) : ( n3303 ) ;
assign n3305 =  ( n2617 ) ? ( bv_8_217_n128 ) : ( n3304 ) ;
assign n3306 =  ( n2615 ) ? ( bv_8_142_n406 ) : ( n3305 ) ;
assign n3307 =  ( n2613 ) ? ( bv_8_148_n388 ) : ( n3306 ) ;
assign n3308 =  ( n2611 ) ? ( bv_8_155_n364 ) : ( n3307 ) ;
assign n3309 =  ( n2609 ) ? ( bv_8_30_n21 ) : ( n3308 ) ;
assign n3310 =  ( n2607 ) ? ( bv_8_135_n81 ) : ( n3309 ) ;
assign n3311 =  ( n2605 ) ? ( bv_8_233_n91 ) : ( n3310 ) ;
assign n3312 =  ( n2603 ) ? ( bv_8_206_n192 ) : ( n3311 ) ;
assign n3313 =  ( n2601 ) ? ( bv_8_85_n423 ) : ( n3312 ) ;
assign n3314 =  ( n2599 ) ? ( bv_8_40_n366 ) : ( n3313 ) ;
assign n3315 =  ( n2597 ) ? ( bv_8_223_n130 ) : ( n3314 ) ;
assign n3316 =  ( n2595 ) ? ( bv_8_140_n376 ) : ( n3315 ) ;
assign n3317 =  ( n2593 ) ? ( bv_8_161_n211 ) : ( n3316 ) ;
assign n3318 =  ( n2591 ) ? ( bv_8_137_n421 ) : ( n3317 ) ;
assign n3319 =  ( n2589 ) ? ( bv_8_13_n194 ) : ( n3318 ) ;
assign n3320 =  ( n2587 ) ? ( bv_8_191_n246 ) : ( n3319 ) ;
assign n3321 =  ( n2585 ) ? ( bv_8_230_n103 ) : ( n3320 ) ;
assign n3322 =  ( n2583 ) ? ( bv_8_66_n466 ) : ( n3321 ) ;
assign n3323 =  ( n2581 ) ? ( bv_8_104_n520 ) : ( n3322 ) ;
assign n3324 =  ( n2579 ) ? ( bv_8_65_n623 ) : ( n3323 ) ;
assign n3325 =  ( n2577 ) ? ( bv_8_153_n140 ) : ( n3324 ) ;
assign n3326 =  ( n2575 ) ? ( bv_8_45_n97 ) : ( n3325 ) ;
assign n3327 =  ( n2573 ) ? ( bv_8_15_n190 ) : ( n3326 ) ;
assign n3328 =  ( n2571 ) ? ( bv_8_176_n299 ) : ( n3327 ) ;
assign n3329 =  ( n2569 ) ? ( bv_8_84_n386 ) : ( n3328 ) ;
assign n3330 =  ( n2567 ) ? ( bv_8_187_n260 ) : ( n3329 ) ;
assign n3331 =  ( n2565 ) ? ( bv_8_22_n357 ) : ( n3330 ) ;
assign n3332 =  ( n2563 ) ^ ( n3331 )  ;
assign n3333 = state_in[7:0] ;
assign n3334 =  ( n3333 ) == ( bv_8_255_n3 )  ;
assign n3335 = state_in[7:0] ;
assign n3336 =  ( n3335 ) == ( bv_8_254_n7 )  ;
assign n3337 = state_in[7:0] ;
assign n3338 =  ( n3337 ) == ( bv_8_253_n11 )  ;
assign n3339 = state_in[7:0] ;
assign n3340 =  ( n3339 ) == ( bv_8_252_n15 )  ;
assign n3341 = state_in[7:0] ;
assign n3342 =  ( n3341 ) == ( bv_8_251_n19 )  ;
assign n3343 = state_in[7:0] ;
assign n3344 =  ( n3343 ) == ( bv_8_250_n23 )  ;
assign n3345 = state_in[7:0] ;
assign n3346 =  ( n3345 ) == ( bv_8_249_n27 )  ;
assign n3347 = state_in[7:0] ;
assign n3348 =  ( n3347 ) == ( bv_8_248_n31 )  ;
assign n3349 = state_in[7:0] ;
assign n3350 =  ( n3349 ) == ( bv_8_247_n35 )  ;
assign n3351 = state_in[7:0] ;
assign n3352 =  ( n3351 ) == ( bv_8_246_n39 )  ;
assign n3353 = state_in[7:0] ;
assign n3354 =  ( n3353 ) == ( bv_8_245_n43 )  ;
assign n3355 = state_in[7:0] ;
assign n3356 =  ( n3355 ) == ( bv_8_244_n47 )  ;
assign n3357 = state_in[7:0] ;
assign n3358 =  ( n3357 ) == ( bv_8_243_n51 )  ;
assign n3359 = state_in[7:0] ;
assign n3360 =  ( n3359 ) == ( bv_8_242_n55 )  ;
assign n3361 = state_in[7:0] ;
assign n3362 =  ( n3361 ) == ( bv_8_241_n59 )  ;
assign n3363 = state_in[7:0] ;
assign n3364 =  ( n3363 ) == ( bv_8_240_n63 )  ;
assign n3365 = state_in[7:0] ;
assign n3366 =  ( n3365 ) == ( bv_8_239_n67 )  ;
assign n3367 = state_in[7:0] ;
assign n3368 =  ( n3367 ) == ( bv_8_238_n71 )  ;
assign n3369 = state_in[7:0] ;
assign n3370 =  ( n3369 ) == ( bv_8_237_n75 )  ;
assign n3371 = state_in[7:0] ;
assign n3372 =  ( n3371 ) == ( bv_8_236_n79 )  ;
assign n3373 = state_in[7:0] ;
assign n3374 =  ( n3373 ) == ( bv_8_235_n83 )  ;
assign n3375 = state_in[7:0] ;
assign n3376 =  ( n3375 ) == ( bv_8_234_n87 )  ;
assign n3377 = state_in[7:0] ;
assign n3378 =  ( n3377 ) == ( bv_8_233_n91 )  ;
assign n3379 = state_in[7:0] ;
assign n3380 =  ( n3379 ) == ( bv_8_232_n95 )  ;
assign n3381 = state_in[7:0] ;
assign n3382 =  ( n3381 ) == ( bv_8_231_n99 )  ;
assign n3383 = state_in[7:0] ;
assign n3384 =  ( n3383 ) == ( bv_8_230_n103 )  ;
assign n3385 = state_in[7:0] ;
assign n3386 =  ( n3385 ) == ( bv_8_229_n107 )  ;
assign n3387 = state_in[7:0] ;
assign n3388 =  ( n3387 ) == ( bv_8_228_n111 )  ;
assign n3389 = state_in[7:0] ;
assign n3390 =  ( n3389 ) == ( bv_8_227_n115 )  ;
assign n3391 = state_in[7:0] ;
assign n3392 =  ( n3391 ) == ( bv_8_226_n119 )  ;
assign n3393 = state_in[7:0] ;
assign n3394 =  ( n3393 ) == ( bv_8_225_n123 )  ;
assign n3395 = state_in[7:0] ;
assign n3396 =  ( n3395 ) == ( bv_8_224_n126 )  ;
assign n3397 = state_in[7:0] ;
assign n3398 =  ( n3397 ) == ( bv_8_223_n130 )  ;
assign n3399 = state_in[7:0] ;
assign n3400 =  ( n3399 ) == ( bv_8_222_n134 )  ;
assign n3401 = state_in[7:0] ;
assign n3402 =  ( n3401 ) == ( bv_8_221_n138 )  ;
assign n3403 = state_in[7:0] ;
assign n3404 =  ( n3403 ) == ( bv_8_220_n142 )  ;
assign n3405 = state_in[7:0] ;
assign n3406 =  ( n3405 ) == ( bv_8_219_n146 )  ;
assign n3407 = state_in[7:0] ;
assign n3408 =  ( n3407 ) == ( bv_8_218_n150 )  ;
assign n3409 = state_in[7:0] ;
assign n3410 =  ( n3409 ) == ( bv_8_217_n128 )  ;
assign n3411 = state_in[7:0] ;
assign n3412 =  ( n3411 ) == ( bv_8_216_n157 )  ;
assign n3413 = state_in[7:0] ;
assign n3414 =  ( n3413 ) == ( bv_8_215_n45 )  ;
assign n3415 = state_in[7:0] ;
assign n3416 =  ( n3415 ) == ( bv_8_214_n164 )  ;
assign n3417 = state_in[7:0] ;
assign n3418 =  ( n3417 ) == ( bv_8_213_n167 )  ;
assign n3419 = state_in[7:0] ;
assign n3420 =  ( n3419 ) == ( bv_8_212_n171 )  ;
assign n3421 = state_in[7:0] ;
assign n3422 =  ( n3421 ) == ( bv_8_211_n175 )  ;
assign n3423 = state_in[7:0] ;
assign n3424 =  ( n3423 ) == ( bv_8_210_n113 )  ;
assign n3425 = state_in[7:0] ;
assign n3426 =  ( n3425 ) == ( bv_8_209_n182 )  ;
assign n3427 = state_in[7:0] ;
assign n3428 =  ( n3427 ) == ( bv_8_208_n37 )  ;
assign n3429 = state_in[7:0] ;
assign n3430 =  ( n3429 ) == ( bv_8_207_n188 )  ;
assign n3431 = state_in[7:0] ;
assign n3432 =  ( n3431 ) == ( bv_8_206_n192 )  ;
assign n3433 = state_in[7:0] ;
assign n3434 =  ( n3433 ) == ( bv_8_205_n196 )  ;
assign n3435 = state_in[7:0] ;
assign n3436 =  ( n3435 ) == ( bv_8_204_n177 )  ;
assign n3437 = state_in[7:0] ;
assign n3438 =  ( n3437 ) == ( bv_8_203_n203 )  ;
assign n3439 = state_in[7:0] ;
assign n3440 =  ( n3439 ) == ( bv_8_202_n207 )  ;
assign n3441 = state_in[7:0] ;
assign n3442 =  ( n3441 ) == ( bv_8_201_n85 )  ;
assign n3443 = state_in[7:0] ;
assign n3444 =  ( n3443 ) == ( bv_8_200_n213 )  ;
assign n3445 = state_in[7:0] ;
assign n3446 =  ( n3445 ) == ( bv_8_199_n216 )  ;
assign n3447 = state_in[7:0] ;
assign n3448 =  ( n3447 ) == ( bv_8_198_n220 )  ;
assign n3449 = state_in[7:0] ;
assign n3450 =  ( n3449 ) == ( bv_8_197_n224 )  ;
assign n3451 = state_in[7:0] ;
assign n3452 =  ( n3451 ) == ( bv_8_196_n228 )  ;
assign n3453 = state_in[7:0] ;
assign n3454 =  ( n3453 ) == ( bv_8_195_n232 )  ;
assign n3455 = state_in[7:0] ;
assign n3456 =  ( n3455 ) == ( bv_8_194_n159 )  ;
assign n3457 = state_in[7:0] ;
assign n3458 =  ( n3457 ) == ( bv_8_193_n239 )  ;
assign n3459 = state_in[7:0] ;
assign n3460 =  ( n3459 ) == ( bv_8_192_n242 )  ;
assign n3461 = state_in[7:0] ;
assign n3462 =  ( n3461 ) == ( bv_8_191_n246 )  ;
assign n3463 = state_in[7:0] ;
assign n3464 =  ( n3463 ) == ( bv_8_190_n250 )  ;
assign n3465 = state_in[7:0] ;
assign n3466 =  ( n3465 ) == ( bv_8_189_n254 )  ;
assign n3467 = state_in[7:0] ;
assign n3468 =  ( n3467 ) == ( bv_8_188_n257 )  ;
assign n3469 = state_in[7:0] ;
assign n3470 =  ( n3469 ) == ( bv_8_187_n260 )  ;
assign n3471 = state_in[7:0] ;
assign n3472 =  ( n3471 ) == ( bv_8_186_n263 )  ;
assign n3473 = state_in[7:0] ;
assign n3474 =  ( n3473 ) == ( bv_8_185_n266 )  ;
assign n3475 = state_in[7:0] ;
assign n3476 =  ( n3475 ) == ( bv_8_184_n270 )  ;
assign n3477 = state_in[7:0] ;
assign n3478 =  ( n3477 ) == ( bv_8_183_n273 )  ;
assign n3479 = state_in[7:0] ;
assign n3480 =  ( n3479 ) == ( bv_8_182_n277 )  ;
assign n3481 = state_in[7:0] ;
assign n3482 =  ( n3481 ) == ( bv_8_181_n281 )  ;
assign n3483 = state_in[7:0] ;
assign n3484 =  ( n3483 ) == ( bv_8_180_n285 )  ;
assign n3485 = state_in[7:0] ;
assign n3486 =  ( n3485 ) == ( bv_8_179_n289 )  ;
assign n3487 = state_in[7:0] ;
assign n3488 =  ( n3487 ) == ( bv_8_178_n292 )  ;
assign n3489 = state_in[7:0] ;
assign n3490 =  ( n3489 ) == ( bv_8_177_n283 )  ;
assign n3491 = state_in[7:0] ;
assign n3492 =  ( n3491 ) == ( bv_8_176_n299 )  ;
assign n3493 = state_in[7:0] ;
assign n3494 =  ( n3493 ) == ( bv_8_175_n302 )  ;
assign n3495 = state_in[7:0] ;
assign n3496 =  ( n3495 ) == ( bv_8_174_n152 )  ;
assign n3497 = state_in[7:0] ;
assign n3498 =  ( n3497 ) == ( bv_8_173_n307 )  ;
assign n3499 = state_in[7:0] ;
assign n3500 =  ( n3499 ) == ( bv_8_172_n268 )  ;
assign n3501 = state_in[7:0] ;
assign n3502 =  ( n3501 ) == ( bv_8_171_n314 )  ;
assign n3503 = state_in[7:0] ;
assign n3504 =  ( n3503 ) == ( bv_8_170_n77 )  ;
assign n3505 = state_in[7:0] ;
assign n3506 =  ( n3505 ) == ( bv_8_169_n109 )  ;
assign n3507 = state_in[7:0] ;
assign n3508 =  ( n3507 ) == ( bv_8_168_n13 )  ;
assign n3509 = state_in[7:0] ;
assign n3510 =  ( n3509 ) == ( bv_8_167_n325 )  ;
assign n3511 = state_in[7:0] ;
assign n3512 =  ( n3511 ) == ( bv_8_166_n328 )  ;
assign n3513 = state_in[7:0] ;
assign n3514 =  ( n3513 ) == ( bv_8_165_n69 )  ;
assign n3515 = state_in[7:0] ;
assign n3516 =  ( n3515 ) == ( bv_8_164_n335 )  ;
assign n3517 = state_in[7:0] ;
assign n3518 =  ( n3517 ) == ( bv_8_163_n339 )  ;
assign n3519 = state_in[7:0] ;
assign n3520 =  ( n3519 ) == ( bv_8_162_n343 )  ;
assign n3521 = state_in[7:0] ;
assign n3522 =  ( n3521 ) == ( bv_8_161_n211 )  ;
assign n3523 = state_in[7:0] ;
assign n3524 =  ( n3523 ) == ( bv_8_160_n350 )  ;
assign n3525 = state_in[7:0] ;
assign n3526 =  ( n3525 ) == ( bv_8_159_n323 )  ;
assign n3527 = state_in[7:0] ;
assign n3528 =  ( n3527 ) == ( bv_8_158_n355 )  ;
assign n3529 = state_in[7:0] ;
assign n3530 =  ( n3529 ) == ( bv_8_157_n359 )  ;
assign n3531 = state_in[7:0] ;
assign n3532 =  ( n3531 ) == ( bv_8_156_n279 )  ;
assign n3533 = state_in[7:0] ;
assign n3534 =  ( n3533 ) == ( bv_8_155_n364 )  ;
assign n3535 = state_in[7:0] ;
assign n3536 =  ( n3535 ) == ( bv_8_154_n368 )  ;
assign n3537 = state_in[7:0] ;
assign n3538 =  ( n3537 ) == ( bv_8_153_n140 )  ;
assign n3539 = state_in[7:0] ;
assign n3540 =  ( n3539 ) == ( bv_8_152_n374 )  ;
assign n3541 = state_in[7:0] ;
assign n3542 =  ( n3541 ) == ( bv_8_151_n218 )  ;
assign n3543 = state_in[7:0] ;
assign n3544 =  ( n3543 ) == ( bv_8_150_n201 )  ;
assign n3545 = state_in[7:0] ;
assign n3546 =  ( n3545 ) == ( bv_8_149_n384 )  ;
assign n3547 = state_in[7:0] ;
assign n3548 =  ( n3547 ) == ( bv_8_148_n388 )  ;
assign n3549 = state_in[7:0] ;
assign n3550 =  ( n3549 ) == ( bv_8_147_n392 )  ;
assign n3551 = state_in[7:0] ;
assign n3552 =  ( n3551 ) == ( bv_8_146_n337 )  ;
assign n3553 = state_in[7:0] ;
assign n3554 =  ( n3553 ) == ( bv_8_145_n397 )  ;
assign n3555 = state_in[7:0] ;
assign n3556 =  ( n3555 ) == ( bv_8_144_n173 )  ;
assign n3557 = state_in[7:0] ;
assign n3558 =  ( n3557 ) == ( bv_8_143_n403 )  ;
assign n3559 = state_in[7:0] ;
assign n3560 =  ( n3559 ) == ( bv_8_142_n406 )  ;
assign n3561 = state_in[7:0] ;
assign n3562 =  ( n3561 ) == ( bv_8_141_n410 )  ;
assign n3563 = state_in[7:0] ;
assign n3564 =  ( n3563 ) == ( bv_8_140_n376 )  ;
assign n3565 = state_in[7:0] ;
assign n3566 =  ( n3565 ) == ( bv_8_139_n297 )  ;
assign n3567 = state_in[7:0] ;
assign n3568 =  ( n3567 ) == ( bv_8_138_n418 )  ;
assign n3569 = state_in[7:0] ;
assign n3570 =  ( n3569 ) == ( bv_8_137_n421 )  ;
assign n3571 = state_in[7:0] ;
assign n3572 =  ( n3571 ) == ( bv_8_136_n425 )  ;
assign n3573 = state_in[7:0] ;
assign n3574 =  ( n3573 ) == ( bv_8_135_n81 )  ;
assign n3575 = state_in[7:0] ;
assign n3576 =  ( n3575 ) == ( bv_8_134_n431 )  ;
assign n3577 = state_in[7:0] ;
assign n3578 =  ( n3577 ) == ( bv_8_133_n434 )  ;
assign n3579 = state_in[7:0] ;
assign n3580 =  ( n3579 ) == ( bv_8_132_n41 )  ;
assign n3581 = state_in[7:0] ;
assign n3582 =  ( n3581 ) == ( bv_8_131_n440 )  ;
assign n3583 = state_in[7:0] ;
assign n3584 =  ( n3583 ) == ( bv_8_130_n33 )  ;
assign n3585 = state_in[7:0] ;
assign n3586 =  ( n3585 ) == ( bv_8_129_n446 )  ;
assign n3587 = state_in[7:0] ;
assign n3588 =  ( n3587 ) == ( bv_8_128_n450 )  ;
assign n3589 = state_in[7:0] ;
assign n3590 =  ( n3589 ) == ( bv_8_127_n453 )  ;
assign n3591 = state_in[7:0] ;
assign n3592 =  ( n3591 ) == ( bv_8_126_n456 )  ;
assign n3593 = state_in[7:0] ;
assign n3594 =  ( n3593 ) == ( bv_8_125_n459 )  ;
assign n3595 = state_in[7:0] ;
assign n3596 =  ( n3595 ) == ( bv_8_124_n184 )  ;
assign n3597 = state_in[7:0] ;
assign n3598 =  ( n3597 ) == ( bv_8_123_n17 )  ;
assign n3599 = state_in[7:0] ;
assign n3600 =  ( n3599 ) == ( bv_8_122_n416 )  ;
assign n3601 = state_in[7:0] ;
assign n3602 =  ( n3601 ) == ( bv_8_121_n470 )  ;
assign n3603 = state_in[7:0] ;
assign n3604 =  ( n3603 ) == ( bv_8_120_n474 )  ;
assign n3605 = state_in[7:0] ;
assign n3606 =  ( n3605 ) == ( bv_8_119_n472 )  ;
assign n3607 = state_in[7:0] ;
assign n3608 =  ( n3607 ) == ( bv_8_118_n480 )  ;
assign n3609 = state_in[7:0] ;
assign n3610 =  ( n3609 ) == ( bv_8_117_n484 )  ;
assign n3611 = state_in[7:0] ;
assign n3612 =  ( n3611 ) == ( bv_8_116_n345 )  ;
assign n3613 = state_in[7:0] ;
assign n3614 =  ( n3613 ) == ( bv_8_115_n222 )  ;
assign n3615 = state_in[7:0] ;
assign n3616 =  ( n3615 ) == ( bv_8_114_n494 )  ;
assign n3617 = state_in[7:0] ;
assign n3618 =  ( n3617 ) == ( bv_8_113_n180 )  ;
assign n3619 = state_in[7:0] ;
assign n3620 =  ( n3619 ) == ( bv_8_112_n482 )  ;
assign n3621 = state_in[7:0] ;
assign n3622 =  ( n3621 ) == ( bv_8_111_n244 )  ;
assign n3623 = state_in[7:0] ;
assign n3624 =  ( n3623 ) == ( bv_8_110_n294 )  ;
assign n3625 = state_in[7:0] ;
assign n3626 =  ( n3625 ) == ( bv_8_109_n9 )  ;
assign n3627 = state_in[7:0] ;
assign n3628 =  ( n3627 ) == ( bv_8_108_n510 )  ;
assign n3629 = state_in[7:0] ;
assign n3630 =  ( n3629 ) == ( bv_8_107_n370 )  ;
assign n3631 = state_in[7:0] ;
assign n3632 =  ( n3631 ) == ( bv_8_106_n155 )  ;
assign n3633 = state_in[7:0] ;
assign n3634 =  ( n3633 ) == ( bv_8_105_n148 )  ;
assign n3635 = state_in[7:0] ;
assign n3636 =  ( n3635 ) == ( bv_8_104_n520 )  ;
assign n3637 = state_in[7:0] ;
assign n3638 =  ( n3637 ) == ( bv_8_103_n523 )  ;
assign n3639 = state_in[7:0] ;
assign n3640 =  ( n3639 ) == ( bv_8_102_n527 )  ;
assign n3641 = state_in[7:0] ;
assign n3642 =  ( n3641 ) == ( bv_8_101_n49 )  ;
assign n3643 = state_in[7:0] ;
assign n3644 =  ( n3643 ) == ( bv_8_100_n348 )  ;
assign n3645 = state_in[7:0] ;
assign n3646 =  ( n3645 ) == ( bv_8_99_n476 )  ;
assign n3647 = state_in[7:0] ;
assign n3648 =  ( n3647 ) == ( bv_8_98_n536 )  ;
assign n3649 = state_in[7:0] ;
assign n3650 =  ( n3649 ) == ( bv_8_97_n198 )  ;
assign n3651 = state_in[7:0] ;
assign n3652 =  ( n3651 ) == ( bv_8_96_n542 )  ;
assign n3653 = state_in[7:0] ;
assign n3654 =  ( n3653 ) == ( bv_8_95_n545 )  ;
assign n3655 = state_in[7:0] ;
assign n3656 =  ( n3655 ) == ( bv_8_94_n548 )  ;
assign n3657 = state_in[7:0] ;
assign n3658 =  ( n3657 ) == ( bv_8_93_n498 )  ;
assign n3659 = state_in[7:0] ;
assign n3660 =  ( n3659 ) == ( bv_8_92_n234 )  ;
assign n3661 = state_in[7:0] ;
assign n3662 =  ( n3661 ) == ( bv_8_91_n555 )  ;
assign n3663 = state_in[7:0] ;
assign n3664 =  ( n3663 ) == ( bv_8_90_n25 )  ;
assign n3665 = state_in[7:0] ;
assign n3666 =  ( n3665 ) == ( bv_8_89_n61 )  ;
assign n3667 = state_in[7:0] ;
assign n3668 =  ( n3667 ) == ( bv_8_88_n562 )  ;
assign n3669 = state_in[7:0] ;
assign n3670 =  ( n3669 ) == ( bv_8_87_n226 )  ;
assign n3671 = state_in[7:0] ;
assign n3672 =  ( n3671 ) == ( bv_8_86_n567 )  ;
assign n3673 = state_in[7:0] ;
assign n3674 =  ( n3673 ) == ( bv_8_85_n423 )  ;
assign n3675 = state_in[7:0] ;
assign n3676 =  ( n3675 ) == ( bv_8_84_n386 )  ;
assign n3677 = state_in[7:0] ;
assign n3678 =  ( n3677 ) == ( bv_8_83_n575 )  ;
assign n3679 = state_in[7:0] ;
assign n3680 =  ( n3679 ) == ( bv_8_82_n578 )  ;
assign n3681 = state_in[7:0] ;
assign n3682 =  ( n3681 ) == ( bv_8_81_n582 )  ;
assign n3683 = state_in[7:0] ;
assign n3684 =  ( n3683 ) == ( bv_8_80_n73 )  ;
assign n3685 = state_in[7:0] ;
assign n3686 =  ( n3685 ) == ( bv_8_79_n538 )  ;
assign n3687 = state_in[7:0] ;
assign n3688 =  ( n3687 ) == ( bv_8_78_n590 )  ;
assign n3689 = state_in[7:0] ;
assign n3690 =  ( n3689 ) == ( bv_8_77_n593 )  ;
assign n3691 = state_in[7:0] ;
assign n3692 =  ( n3691 ) == ( bv_8_76_n596 )  ;
assign n3693 = state_in[7:0] ;
assign n3694 =  ( n3693 ) == ( bv_8_75_n503 )  ;
assign n3695 = state_in[7:0] ;
assign n3696 =  ( n3695 ) == ( bv_8_74_n237 )  ;
assign n3697 = state_in[7:0] ;
assign n3698 =  ( n3697 ) == ( bv_8_73_n275 )  ;
assign n3699 = state_in[7:0] ;
assign n3700 =  ( n3699 ) == ( bv_8_72_n330 )  ;
assign n3701 = state_in[7:0] ;
assign n3702 =  ( n3701 ) == ( bv_8_71_n252 )  ;
assign n3703 = state_in[7:0] ;
assign n3704 =  ( n3703 ) == ( bv_8_70_n609 )  ;
assign n3705 = state_in[7:0] ;
assign n3706 =  ( n3705 ) == ( bv_8_69_n612 )  ;
assign n3707 = state_in[7:0] ;
assign n3708 =  ( n3707 ) == ( bv_8_68_n390 )  ;
assign n3709 = state_in[7:0] ;
assign n3710 =  ( n3709 ) == ( bv_8_67_n318 )  ;
assign n3711 = state_in[7:0] ;
assign n3712 =  ( n3711 ) == ( bv_8_66_n466 )  ;
assign n3713 = state_in[7:0] ;
assign n3714 =  ( n3713 ) == ( bv_8_65_n623 )  ;
assign n3715 = state_in[7:0] ;
assign n3716 =  ( n3715 ) == ( bv_8_64_n573 )  ;
assign n3717 = state_in[7:0] ;
assign n3718 =  ( n3717 ) == ( bv_8_63_n489 )  ;
assign n3719 = state_in[7:0] ;
assign n3720 =  ( n3719 ) == ( bv_8_62_n205 )  ;
assign n3721 = state_in[7:0] ;
assign n3722 =  ( n3721 ) == ( bv_8_61_n634 )  ;
assign n3723 = state_in[7:0] ;
assign n3724 =  ( n3723 ) == ( bv_8_60_n93 )  ;
assign n3725 = state_in[7:0] ;
assign n3726 =  ( n3725 ) == ( bv_8_59_n382 )  ;
assign n3727 = state_in[7:0] ;
assign n3728 =  ( n3727 ) == ( bv_8_58_n136 )  ;
assign n3729 = state_in[7:0] ;
assign n3730 =  ( n3729 ) == ( bv_8_57_n312 )  ;
assign n3731 = state_in[7:0] ;
assign n3732 =  ( n3731 ) == ( bv_8_56_n230 )  ;
assign n3733 = state_in[7:0] ;
assign n3734 =  ( n3733 ) == ( bv_8_55_n650 )  ;
assign n3735 = state_in[7:0] ;
assign n3736 =  ( n3735 ) == ( bv_8_54_n616 )  ;
assign n3737 = state_in[7:0] ;
assign n3738 =  ( n3737 ) == ( bv_8_53_n436 )  ;
assign n3739 = state_in[7:0] ;
assign n3740 =  ( n3739 ) == ( bv_8_52_n619 )  ;
assign n3741 = state_in[7:0] ;
assign n3742 =  ( n3741 ) == ( bv_8_51_n101 )  ;
assign n3743 = state_in[7:0] ;
assign n3744 =  ( n3743 ) == ( bv_8_50_n408 )  ;
assign n3745 = state_in[7:0] ;
assign n3746 =  ( n3745 ) == ( bv_8_49_n309 )  ;
assign n3747 = state_in[7:0] ;
assign n3748 =  ( n3747 ) == ( bv_8_48_n660 )  ;
assign n3749 = state_in[7:0] ;
assign n3750 =  ( n3749 ) == ( bv_8_47_n652 )  ;
assign n3751 = state_in[7:0] ;
assign n3752 =  ( n3751 ) == ( bv_8_46_n429 )  ;
assign n3753 = state_in[7:0] ;
assign n3754 =  ( n3753 ) == ( bv_8_45_n97 )  ;
assign n3755 = state_in[7:0] ;
assign n3756 =  ( n3755 ) == ( bv_8_44_n5 )  ;
assign n3757 = state_in[7:0] ;
assign n3758 =  ( n3757 ) == ( bv_8_43_n121 )  ;
assign n3759 = state_in[7:0] ;
assign n3760 =  ( n3759 ) == ( bv_8_42_n672 )  ;
assign n3761 = state_in[7:0] ;
assign n3762 =  ( n3761 ) == ( bv_8_41_n29 )  ;
assign n3763 = state_in[7:0] ;
assign n3764 =  ( n3763 ) == ( bv_8_40_n366 )  ;
assign n3765 = state_in[7:0] ;
assign n3766 =  ( n3765 ) == ( bv_8_39_n132 )  ;
assign n3767 = state_in[7:0] ;
assign n3768 =  ( n3767 ) == ( bv_8_38_n444 )  ;
assign n3769 = state_in[7:0] ;
assign n3770 =  ( n3769 ) == ( bv_8_37_n506 )  ;
assign n3771 = state_in[7:0] ;
assign n3772 =  ( n3771 ) == ( bv_8_36_n645 )  ;
assign n3773 = state_in[7:0] ;
assign n3774 =  ( n3773 ) == ( bv_8_35_n696 )  ;
assign n3775 = state_in[7:0] ;
assign n3776 =  ( n3775 ) == ( bv_8_34_n117 )  ;
assign n3777 = state_in[7:0] ;
assign n3778 =  ( n3777 ) == ( bv_8_33_n486 )  ;
assign n3779 = state_in[7:0] ;
assign n3780 =  ( n3779 ) == ( bv_8_32_n463 )  ;
assign n3781 = state_in[7:0] ;
assign n3782 =  ( n3781 ) == ( bv_8_31_n705 )  ;
assign n3783 = state_in[7:0] ;
assign n3784 =  ( n3783 ) == ( bv_8_30_n21 )  ;
assign n3785 = state_in[7:0] ;
assign n3786 =  ( n3785 ) == ( bv_8_29_n625 )  ;
assign n3787 = state_in[7:0] ;
assign n3788 =  ( n3787 ) == ( bv_8_28_n162 )  ;
assign n3789 = state_in[7:0] ;
assign n3790 =  ( n3789 ) == ( bv_8_27_n642 )  ;
assign n3791 = state_in[7:0] ;
assign n3792 =  ( n3791 ) == ( bv_8_26_n53 )  ;
assign n3793 = state_in[7:0] ;
assign n3794 =  ( n3793 ) == ( bv_8_25_n399 )  ;
assign n3795 = state_in[7:0] ;
assign n3796 =  ( n3795 ) == ( bv_8_24_n448 )  ;
assign n3797 = state_in[7:0] ;
assign n3798 =  ( n3797 ) == ( bv_8_23_n144 )  ;
assign n3799 = state_in[7:0] ;
assign n3800 =  ( n3799 ) == ( bv_8_22_n357 )  ;
assign n3801 = state_in[7:0] ;
assign n3802 =  ( n3801 ) == ( bv_8_21_n89 )  ;
assign n3803 = state_in[7:0] ;
assign n3804 =  ( n3803 ) == ( bv_8_20_n341 )  ;
assign n3805 = state_in[7:0] ;
assign n3806 =  ( n3805 ) == ( bv_8_19_n588 )  ;
assign n3807 = state_in[7:0] ;
assign n3808 =  ( n3807 ) == ( bv_8_18_n628 )  ;
assign n3809 = state_in[7:0] ;
assign n3810 =  ( n3809 ) == ( bv_8_17_n525 )  ;
assign n3811 = state_in[7:0] ;
assign n3812 =  ( n3811 ) == ( bv_8_16_n248 )  ;
assign n3813 = state_in[7:0] ;
assign n3814 =  ( n3813 ) == ( bv_8_15_n190 )  ;
assign n3815 = state_in[7:0] ;
assign n3816 =  ( n3815 ) == ( bv_8_14_n648 )  ;
assign n3817 = state_in[7:0] ;
assign n3818 =  ( n3817 ) == ( bv_8_13_n194 )  ;
assign n3819 = state_in[7:0] ;
assign n3820 =  ( n3819 ) == ( bv_8_12_n333 )  ;
assign n3821 = state_in[7:0] ;
assign n3822 =  ( n3821 ) == ( bv_8_11_n379 )  ;
assign n3823 = state_in[7:0] ;
assign n3824 =  ( n3823 ) == ( bv_8_10_n655 )  ;
assign n3825 = state_in[7:0] ;
assign n3826 =  ( n3825 ) == ( bv_8_9_n57 )  ;
assign n3827 = state_in[7:0] ;
assign n3828 =  ( n3827 ) == ( bv_8_8_n669 )  ;
assign n3829 = state_in[7:0] ;
assign n3830 =  ( n3829 ) == ( bv_8_7_n105 )  ;
assign n3831 = state_in[7:0] ;
assign n3832 =  ( n3831 ) == ( bv_8_6_n169 )  ;
assign n3833 = state_in[7:0] ;
assign n3834 =  ( n3833 ) == ( bv_8_5_n492 )  ;
assign n3835 = state_in[7:0] ;
assign n3836 =  ( n3835 ) == ( bv_8_4_n516 )  ;
assign n3837 = state_in[7:0] ;
assign n3838 =  ( n3837 ) == ( bv_8_3_n65 )  ;
assign n3839 = state_in[7:0] ;
assign n3840 =  ( n3839 ) == ( bv_8_2_n751 )  ;
assign n3841 = state_in[7:0] ;
assign n3842 =  ( n3841 ) == ( bv_8_1_n287 )  ;
assign n3843 = state_in[7:0] ;
assign n3844 =  ( n3843 ) == ( bv_8_0_n580 )  ;
assign n3845 =  ( n3844 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n3846 =  ( n3842 ) ? ( bv_8_124_n184 ) : ( n3845 ) ;
assign n3847 =  ( n3840 ) ? ( bv_8_119_n472 ) : ( n3846 ) ;
assign n3848 =  ( n3838 ) ? ( bv_8_123_n17 ) : ( n3847 ) ;
assign n3849 =  ( n3836 ) ? ( bv_8_242_n55 ) : ( n3848 ) ;
assign n3850 =  ( n3834 ) ? ( bv_8_107_n370 ) : ( n3849 ) ;
assign n3851 =  ( n3832 ) ? ( bv_8_111_n244 ) : ( n3850 ) ;
assign n3852 =  ( n3830 ) ? ( bv_8_197_n224 ) : ( n3851 ) ;
assign n3853 =  ( n3828 ) ? ( bv_8_48_n660 ) : ( n3852 ) ;
assign n3854 =  ( n3826 ) ? ( bv_8_1_n287 ) : ( n3853 ) ;
assign n3855 =  ( n3824 ) ? ( bv_8_103_n523 ) : ( n3854 ) ;
assign n3856 =  ( n3822 ) ? ( bv_8_43_n121 ) : ( n3855 ) ;
assign n3857 =  ( n3820 ) ? ( bv_8_254_n7 ) : ( n3856 ) ;
assign n3858 =  ( n3818 ) ? ( bv_8_215_n45 ) : ( n3857 ) ;
assign n3859 =  ( n3816 ) ? ( bv_8_171_n314 ) : ( n3858 ) ;
assign n3860 =  ( n3814 ) ? ( bv_8_118_n480 ) : ( n3859 ) ;
assign n3861 =  ( n3812 ) ? ( bv_8_202_n207 ) : ( n3860 ) ;
assign n3862 =  ( n3810 ) ? ( bv_8_130_n33 ) : ( n3861 ) ;
assign n3863 =  ( n3808 ) ? ( bv_8_201_n85 ) : ( n3862 ) ;
assign n3864 =  ( n3806 ) ? ( bv_8_125_n459 ) : ( n3863 ) ;
assign n3865 =  ( n3804 ) ? ( bv_8_250_n23 ) : ( n3864 ) ;
assign n3866 =  ( n3802 ) ? ( bv_8_89_n61 ) : ( n3865 ) ;
assign n3867 =  ( n3800 ) ? ( bv_8_71_n252 ) : ( n3866 ) ;
assign n3868 =  ( n3798 ) ? ( bv_8_240_n63 ) : ( n3867 ) ;
assign n3869 =  ( n3796 ) ? ( bv_8_173_n307 ) : ( n3868 ) ;
assign n3870 =  ( n3794 ) ? ( bv_8_212_n171 ) : ( n3869 ) ;
assign n3871 =  ( n3792 ) ? ( bv_8_162_n343 ) : ( n3870 ) ;
assign n3872 =  ( n3790 ) ? ( bv_8_175_n302 ) : ( n3871 ) ;
assign n3873 =  ( n3788 ) ? ( bv_8_156_n279 ) : ( n3872 ) ;
assign n3874 =  ( n3786 ) ? ( bv_8_164_n335 ) : ( n3873 ) ;
assign n3875 =  ( n3784 ) ? ( bv_8_114_n494 ) : ( n3874 ) ;
assign n3876 =  ( n3782 ) ? ( bv_8_192_n242 ) : ( n3875 ) ;
assign n3877 =  ( n3780 ) ? ( bv_8_183_n273 ) : ( n3876 ) ;
assign n3878 =  ( n3778 ) ? ( bv_8_253_n11 ) : ( n3877 ) ;
assign n3879 =  ( n3776 ) ? ( bv_8_147_n392 ) : ( n3878 ) ;
assign n3880 =  ( n3774 ) ? ( bv_8_38_n444 ) : ( n3879 ) ;
assign n3881 =  ( n3772 ) ? ( bv_8_54_n616 ) : ( n3880 ) ;
assign n3882 =  ( n3770 ) ? ( bv_8_63_n489 ) : ( n3881 ) ;
assign n3883 =  ( n3768 ) ? ( bv_8_247_n35 ) : ( n3882 ) ;
assign n3884 =  ( n3766 ) ? ( bv_8_204_n177 ) : ( n3883 ) ;
assign n3885 =  ( n3764 ) ? ( bv_8_52_n619 ) : ( n3884 ) ;
assign n3886 =  ( n3762 ) ? ( bv_8_165_n69 ) : ( n3885 ) ;
assign n3887 =  ( n3760 ) ? ( bv_8_229_n107 ) : ( n3886 ) ;
assign n3888 =  ( n3758 ) ? ( bv_8_241_n59 ) : ( n3887 ) ;
assign n3889 =  ( n3756 ) ? ( bv_8_113_n180 ) : ( n3888 ) ;
assign n3890 =  ( n3754 ) ? ( bv_8_216_n157 ) : ( n3889 ) ;
assign n3891 =  ( n3752 ) ? ( bv_8_49_n309 ) : ( n3890 ) ;
assign n3892 =  ( n3750 ) ? ( bv_8_21_n89 ) : ( n3891 ) ;
assign n3893 =  ( n3748 ) ? ( bv_8_4_n516 ) : ( n3892 ) ;
assign n3894 =  ( n3746 ) ? ( bv_8_199_n216 ) : ( n3893 ) ;
assign n3895 =  ( n3744 ) ? ( bv_8_35_n696 ) : ( n3894 ) ;
assign n3896 =  ( n3742 ) ? ( bv_8_195_n232 ) : ( n3895 ) ;
assign n3897 =  ( n3740 ) ? ( bv_8_24_n448 ) : ( n3896 ) ;
assign n3898 =  ( n3738 ) ? ( bv_8_150_n201 ) : ( n3897 ) ;
assign n3899 =  ( n3736 ) ? ( bv_8_5_n492 ) : ( n3898 ) ;
assign n3900 =  ( n3734 ) ? ( bv_8_154_n368 ) : ( n3899 ) ;
assign n3901 =  ( n3732 ) ? ( bv_8_7_n105 ) : ( n3900 ) ;
assign n3902 =  ( n3730 ) ? ( bv_8_18_n628 ) : ( n3901 ) ;
assign n3903 =  ( n3728 ) ? ( bv_8_128_n450 ) : ( n3902 ) ;
assign n3904 =  ( n3726 ) ? ( bv_8_226_n119 ) : ( n3903 ) ;
assign n3905 =  ( n3724 ) ? ( bv_8_235_n83 ) : ( n3904 ) ;
assign n3906 =  ( n3722 ) ? ( bv_8_39_n132 ) : ( n3905 ) ;
assign n3907 =  ( n3720 ) ? ( bv_8_178_n292 ) : ( n3906 ) ;
assign n3908 =  ( n3718 ) ? ( bv_8_117_n484 ) : ( n3907 ) ;
assign n3909 =  ( n3716 ) ? ( bv_8_9_n57 ) : ( n3908 ) ;
assign n3910 =  ( n3714 ) ? ( bv_8_131_n440 ) : ( n3909 ) ;
assign n3911 =  ( n3712 ) ? ( bv_8_44_n5 ) : ( n3910 ) ;
assign n3912 =  ( n3710 ) ? ( bv_8_26_n53 ) : ( n3911 ) ;
assign n3913 =  ( n3708 ) ? ( bv_8_27_n642 ) : ( n3912 ) ;
assign n3914 =  ( n3706 ) ? ( bv_8_110_n294 ) : ( n3913 ) ;
assign n3915 =  ( n3704 ) ? ( bv_8_90_n25 ) : ( n3914 ) ;
assign n3916 =  ( n3702 ) ? ( bv_8_160_n350 ) : ( n3915 ) ;
assign n3917 =  ( n3700 ) ? ( bv_8_82_n578 ) : ( n3916 ) ;
assign n3918 =  ( n3698 ) ? ( bv_8_59_n382 ) : ( n3917 ) ;
assign n3919 =  ( n3696 ) ? ( bv_8_214_n164 ) : ( n3918 ) ;
assign n3920 =  ( n3694 ) ? ( bv_8_179_n289 ) : ( n3919 ) ;
assign n3921 =  ( n3692 ) ? ( bv_8_41_n29 ) : ( n3920 ) ;
assign n3922 =  ( n3690 ) ? ( bv_8_227_n115 ) : ( n3921 ) ;
assign n3923 =  ( n3688 ) ? ( bv_8_47_n652 ) : ( n3922 ) ;
assign n3924 =  ( n3686 ) ? ( bv_8_132_n41 ) : ( n3923 ) ;
assign n3925 =  ( n3684 ) ? ( bv_8_83_n575 ) : ( n3924 ) ;
assign n3926 =  ( n3682 ) ? ( bv_8_209_n182 ) : ( n3925 ) ;
assign n3927 =  ( n3680 ) ? ( bv_8_0_n580 ) : ( n3926 ) ;
assign n3928 =  ( n3678 ) ? ( bv_8_237_n75 ) : ( n3927 ) ;
assign n3929 =  ( n3676 ) ? ( bv_8_32_n463 ) : ( n3928 ) ;
assign n3930 =  ( n3674 ) ? ( bv_8_252_n15 ) : ( n3929 ) ;
assign n3931 =  ( n3672 ) ? ( bv_8_177_n283 ) : ( n3930 ) ;
assign n3932 =  ( n3670 ) ? ( bv_8_91_n555 ) : ( n3931 ) ;
assign n3933 =  ( n3668 ) ? ( bv_8_106_n155 ) : ( n3932 ) ;
assign n3934 =  ( n3666 ) ? ( bv_8_203_n203 ) : ( n3933 ) ;
assign n3935 =  ( n3664 ) ? ( bv_8_190_n250 ) : ( n3934 ) ;
assign n3936 =  ( n3662 ) ? ( bv_8_57_n312 ) : ( n3935 ) ;
assign n3937 =  ( n3660 ) ? ( bv_8_74_n237 ) : ( n3936 ) ;
assign n3938 =  ( n3658 ) ? ( bv_8_76_n596 ) : ( n3937 ) ;
assign n3939 =  ( n3656 ) ? ( bv_8_88_n562 ) : ( n3938 ) ;
assign n3940 =  ( n3654 ) ? ( bv_8_207_n188 ) : ( n3939 ) ;
assign n3941 =  ( n3652 ) ? ( bv_8_208_n37 ) : ( n3940 ) ;
assign n3942 =  ( n3650 ) ? ( bv_8_239_n67 ) : ( n3941 ) ;
assign n3943 =  ( n3648 ) ? ( bv_8_170_n77 ) : ( n3942 ) ;
assign n3944 =  ( n3646 ) ? ( bv_8_251_n19 ) : ( n3943 ) ;
assign n3945 =  ( n3644 ) ? ( bv_8_67_n318 ) : ( n3944 ) ;
assign n3946 =  ( n3642 ) ? ( bv_8_77_n593 ) : ( n3945 ) ;
assign n3947 =  ( n3640 ) ? ( bv_8_51_n101 ) : ( n3946 ) ;
assign n3948 =  ( n3638 ) ? ( bv_8_133_n434 ) : ( n3947 ) ;
assign n3949 =  ( n3636 ) ? ( bv_8_69_n612 ) : ( n3948 ) ;
assign n3950 =  ( n3634 ) ? ( bv_8_249_n27 ) : ( n3949 ) ;
assign n3951 =  ( n3632 ) ? ( bv_8_2_n751 ) : ( n3950 ) ;
assign n3952 =  ( n3630 ) ? ( bv_8_127_n453 ) : ( n3951 ) ;
assign n3953 =  ( n3628 ) ? ( bv_8_80_n73 ) : ( n3952 ) ;
assign n3954 =  ( n3626 ) ? ( bv_8_60_n93 ) : ( n3953 ) ;
assign n3955 =  ( n3624 ) ? ( bv_8_159_n323 ) : ( n3954 ) ;
assign n3956 =  ( n3622 ) ? ( bv_8_168_n13 ) : ( n3955 ) ;
assign n3957 =  ( n3620 ) ? ( bv_8_81_n582 ) : ( n3956 ) ;
assign n3958 =  ( n3618 ) ? ( bv_8_163_n339 ) : ( n3957 ) ;
assign n3959 =  ( n3616 ) ? ( bv_8_64_n573 ) : ( n3958 ) ;
assign n3960 =  ( n3614 ) ? ( bv_8_143_n403 ) : ( n3959 ) ;
assign n3961 =  ( n3612 ) ? ( bv_8_146_n337 ) : ( n3960 ) ;
assign n3962 =  ( n3610 ) ? ( bv_8_157_n359 ) : ( n3961 ) ;
assign n3963 =  ( n3608 ) ? ( bv_8_56_n230 ) : ( n3962 ) ;
assign n3964 =  ( n3606 ) ? ( bv_8_245_n43 ) : ( n3963 ) ;
assign n3965 =  ( n3604 ) ? ( bv_8_188_n257 ) : ( n3964 ) ;
assign n3966 =  ( n3602 ) ? ( bv_8_182_n277 ) : ( n3965 ) ;
assign n3967 =  ( n3600 ) ? ( bv_8_218_n150 ) : ( n3966 ) ;
assign n3968 =  ( n3598 ) ? ( bv_8_33_n486 ) : ( n3967 ) ;
assign n3969 =  ( n3596 ) ? ( bv_8_16_n248 ) : ( n3968 ) ;
assign n3970 =  ( n3594 ) ? ( bv_8_255_n3 ) : ( n3969 ) ;
assign n3971 =  ( n3592 ) ? ( bv_8_243_n51 ) : ( n3970 ) ;
assign n3972 =  ( n3590 ) ? ( bv_8_210_n113 ) : ( n3971 ) ;
assign n3973 =  ( n3588 ) ? ( bv_8_205_n196 ) : ( n3972 ) ;
assign n3974 =  ( n3586 ) ? ( bv_8_12_n333 ) : ( n3973 ) ;
assign n3975 =  ( n3584 ) ? ( bv_8_19_n588 ) : ( n3974 ) ;
assign n3976 =  ( n3582 ) ? ( bv_8_236_n79 ) : ( n3975 ) ;
assign n3977 =  ( n3580 ) ? ( bv_8_95_n545 ) : ( n3976 ) ;
assign n3978 =  ( n3578 ) ? ( bv_8_151_n218 ) : ( n3977 ) ;
assign n3979 =  ( n3576 ) ? ( bv_8_68_n390 ) : ( n3978 ) ;
assign n3980 =  ( n3574 ) ? ( bv_8_23_n144 ) : ( n3979 ) ;
assign n3981 =  ( n3572 ) ? ( bv_8_196_n228 ) : ( n3980 ) ;
assign n3982 =  ( n3570 ) ? ( bv_8_167_n325 ) : ( n3981 ) ;
assign n3983 =  ( n3568 ) ? ( bv_8_126_n456 ) : ( n3982 ) ;
assign n3984 =  ( n3566 ) ? ( bv_8_61_n634 ) : ( n3983 ) ;
assign n3985 =  ( n3564 ) ? ( bv_8_100_n348 ) : ( n3984 ) ;
assign n3986 =  ( n3562 ) ? ( bv_8_93_n498 ) : ( n3985 ) ;
assign n3987 =  ( n3560 ) ? ( bv_8_25_n399 ) : ( n3986 ) ;
assign n3988 =  ( n3558 ) ? ( bv_8_115_n222 ) : ( n3987 ) ;
assign n3989 =  ( n3556 ) ? ( bv_8_96_n542 ) : ( n3988 ) ;
assign n3990 =  ( n3554 ) ? ( bv_8_129_n446 ) : ( n3989 ) ;
assign n3991 =  ( n3552 ) ? ( bv_8_79_n538 ) : ( n3990 ) ;
assign n3992 =  ( n3550 ) ? ( bv_8_220_n142 ) : ( n3991 ) ;
assign n3993 =  ( n3548 ) ? ( bv_8_34_n117 ) : ( n3992 ) ;
assign n3994 =  ( n3546 ) ? ( bv_8_42_n672 ) : ( n3993 ) ;
assign n3995 =  ( n3544 ) ? ( bv_8_144_n173 ) : ( n3994 ) ;
assign n3996 =  ( n3542 ) ? ( bv_8_136_n425 ) : ( n3995 ) ;
assign n3997 =  ( n3540 ) ? ( bv_8_70_n609 ) : ( n3996 ) ;
assign n3998 =  ( n3538 ) ? ( bv_8_238_n71 ) : ( n3997 ) ;
assign n3999 =  ( n3536 ) ? ( bv_8_184_n270 ) : ( n3998 ) ;
assign n4000 =  ( n3534 ) ? ( bv_8_20_n341 ) : ( n3999 ) ;
assign n4001 =  ( n3532 ) ? ( bv_8_222_n134 ) : ( n4000 ) ;
assign n4002 =  ( n3530 ) ? ( bv_8_94_n548 ) : ( n4001 ) ;
assign n4003 =  ( n3528 ) ? ( bv_8_11_n379 ) : ( n4002 ) ;
assign n4004 =  ( n3526 ) ? ( bv_8_219_n146 ) : ( n4003 ) ;
assign n4005 =  ( n3524 ) ? ( bv_8_224_n126 ) : ( n4004 ) ;
assign n4006 =  ( n3522 ) ? ( bv_8_50_n408 ) : ( n4005 ) ;
assign n4007 =  ( n3520 ) ? ( bv_8_58_n136 ) : ( n4006 ) ;
assign n4008 =  ( n3518 ) ? ( bv_8_10_n655 ) : ( n4007 ) ;
assign n4009 =  ( n3516 ) ? ( bv_8_73_n275 ) : ( n4008 ) ;
assign n4010 =  ( n3514 ) ? ( bv_8_6_n169 ) : ( n4009 ) ;
assign n4011 =  ( n3512 ) ? ( bv_8_36_n645 ) : ( n4010 ) ;
assign n4012 =  ( n3510 ) ? ( bv_8_92_n234 ) : ( n4011 ) ;
assign n4013 =  ( n3508 ) ? ( bv_8_194_n159 ) : ( n4012 ) ;
assign n4014 =  ( n3506 ) ? ( bv_8_211_n175 ) : ( n4013 ) ;
assign n4015 =  ( n3504 ) ? ( bv_8_172_n268 ) : ( n4014 ) ;
assign n4016 =  ( n3502 ) ? ( bv_8_98_n536 ) : ( n4015 ) ;
assign n4017 =  ( n3500 ) ? ( bv_8_145_n397 ) : ( n4016 ) ;
assign n4018 =  ( n3498 ) ? ( bv_8_149_n384 ) : ( n4017 ) ;
assign n4019 =  ( n3496 ) ? ( bv_8_228_n111 ) : ( n4018 ) ;
assign n4020 =  ( n3494 ) ? ( bv_8_121_n470 ) : ( n4019 ) ;
assign n4021 =  ( n3492 ) ? ( bv_8_231_n99 ) : ( n4020 ) ;
assign n4022 =  ( n3490 ) ? ( bv_8_200_n213 ) : ( n4021 ) ;
assign n4023 =  ( n3488 ) ? ( bv_8_55_n650 ) : ( n4022 ) ;
assign n4024 =  ( n3486 ) ? ( bv_8_109_n9 ) : ( n4023 ) ;
assign n4025 =  ( n3484 ) ? ( bv_8_141_n410 ) : ( n4024 ) ;
assign n4026 =  ( n3482 ) ? ( bv_8_213_n167 ) : ( n4025 ) ;
assign n4027 =  ( n3480 ) ? ( bv_8_78_n590 ) : ( n4026 ) ;
assign n4028 =  ( n3478 ) ? ( bv_8_169_n109 ) : ( n4027 ) ;
assign n4029 =  ( n3476 ) ? ( bv_8_108_n510 ) : ( n4028 ) ;
assign n4030 =  ( n3474 ) ? ( bv_8_86_n567 ) : ( n4029 ) ;
assign n4031 =  ( n3472 ) ? ( bv_8_244_n47 ) : ( n4030 ) ;
assign n4032 =  ( n3470 ) ? ( bv_8_234_n87 ) : ( n4031 ) ;
assign n4033 =  ( n3468 ) ? ( bv_8_101_n49 ) : ( n4032 ) ;
assign n4034 =  ( n3466 ) ? ( bv_8_122_n416 ) : ( n4033 ) ;
assign n4035 =  ( n3464 ) ? ( bv_8_174_n152 ) : ( n4034 ) ;
assign n4036 =  ( n3462 ) ? ( bv_8_8_n669 ) : ( n4035 ) ;
assign n4037 =  ( n3460 ) ? ( bv_8_186_n263 ) : ( n4036 ) ;
assign n4038 =  ( n3458 ) ? ( bv_8_120_n474 ) : ( n4037 ) ;
assign n4039 =  ( n3456 ) ? ( bv_8_37_n506 ) : ( n4038 ) ;
assign n4040 =  ( n3454 ) ? ( bv_8_46_n429 ) : ( n4039 ) ;
assign n4041 =  ( n3452 ) ? ( bv_8_28_n162 ) : ( n4040 ) ;
assign n4042 =  ( n3450 ) ? ( bv_8_166_n328 ) : ( n4041 ) ;
assign n4043 =  ( n3448 ) ? ( bv_8_180_n285 ) : ( n4042 ) ;
assign n4044 =  ( n3446 ) ? ( bv_8_198_n220 ) : ( n4043 ) ;
assign n4045 =  ( n3444 ) ? ( bv_8_232_n95 ) : ( n4044 ) ;
assign n4046 =  ( n3442 ) ? ( bv_8_221_n138 ) : ( n4045 ) ;
assign n4047 =  ( n3440 ) ? ( bv_8_116_n345 ) : ( n4046 ) ;
assign n4048 =  ( n3438 ) ? ( bv_8_31_n705 ) : ( n4047 ) ;
assign n4049 =  ( n3436 ) ? ( bv_8_75_n503 ) : ( n4048 ) ;
assign n4050 =  ( n3434 ) ? ( bv_8_189_n254 ) : ( n4049 ) ;
assign n4051 =  ( n3432 ) ? ( bv_8_139_n297 ) : ( n4050 ) ;
assign n4052 =  ( n3430 ) ? ( bv_8_138_n418 ) : ( n4051 ) ;
assign n4053 =  ( n3428 ) ? ( bv_8_112_n482 ) : ( n4052 ) ;
assign n4054 =  ( n3426 ) ? ( bv_8_62_n205 ) : ( n4053 ) ;
assign n4055 =  ( n3424 ) ? ( bv_8_181_n281 ) : ( n4054 ) ;
assign n4056 =  ( n3422 ) ? ( bv_8_102_n527 ) : ( n4055 ) ;
assign n4057 =  ( n3420 ) ? ( bv_8_72_n330 ) : ( n4056 ) ;
assign n4058 =  ( n3418 ) ? ( bv_8_3_n65 ) : ( n4057 ) ;
assign n4059 =  ( n3416 ) ? ( bv_8_246_n39 ) : ( n4058 ) ;
assign n4060 =  ( n3414 ) ? ( bv_8_14_n648 ) : ( n4059 ) ;
assign n4061 =  ( n3412 ) ? ( bv_8_97_n198 ) : ( n4060 ) ;
assign n4062 =  ( n3410 ) ? ( bv_8_53_n436 ) : ( n4061 ) ;
assign n4063 =  ( n3408 ) ? ( bv_8_87_n226 ) : ( n4062 ) ;
assign n4064 =  ( n3406 ) ? ( bv_8_185_n266 ) : ( n4063 ) ;
assign n4065 =  ( n3404 ) ? ( bv_8_134_n431 ) : ( n4064 ) ;
assign n4066 =  ( n3402 ) ? ( bv_8_193_n239 ) : ( n4065 ) ;
assign n4067 =  ( n3400 ) ? ( bv_8_29_n625 ) : ( n4066 ) ;
assign n4068 =  ( n3398 ) ? ( bv_8_158_n355 ) : ( n4067 ) ;
assign n4069 =  ( n3396 ) ? ( bv_8_225_n123 ) : ( n4068 ) ;
assign n4070 =  ( n3394 ) ? ( bv_8_248_n31 ) : ( n4069 ) ;
assign n4071 =  ( n3392 ) ? ( bv_8_152_n374 ) : ( n4070 ) ;
assign n4072 =  ( n3390 ) ? ( bv_8_17_n525 ) : ( n4071 ) ;
assign n4073 =  ( n3388 ) ? ( bv_8_105_n148 ) : ( n4072 ) ;
assign n4074 =  ( n3386 ) ? ( bv_8_217_n128 ) : ( n4073 ) ;
assign n4075 =  ( n3384 ) ? ( bv_8_142_n406 ) : ( n4074 ) ;
assign n4076 =  ( n3382 ) ? ( bv_8_148_n388 ) : ( n4075 ) ;
assign n4077 =  ( n3380 ) ? ( bv_8_155_n364 ) : ( n4076 ) ;
assign n4078 =  ( n3378 ) ? ( bv_8_30_n21 ) : ( n4077 ) ;
assign n4079 =  ( n3376 ) ? ( bv_8_135_n81 ) : ( n4078 ) ;
assign n4080 =  ( n3374 ) ? ( bv_8_233_n91 ) : ( n4079 ) ;
assign n4081 =  ( n3372 ) ? ( bv_8_206_n192 ) : ( n4080 ) ;
assign n4082 =  ( n3370 ) ? ( bv_8_85_n423 ) : ( n4081 ) ;
assign n4083 =  ( n3368 ) ? ( bv_8_40_n366 ) : ( n4082 ) ;
assign n4084 =  ( n3366 ) ? ( bv_8_223_n130 ) : ( n4083 ) ;
assign n4085 =  ( n3364 ) ? ( bv_8_140_n376 ) : ( n4084 ) ;
assign n4086 =  ( n3362 ) ? ( bv_8_161_n211 ) : ( n4085 ) ;
assign n4087 =  ( n3360 ) ? ( bv_8_137_n421 ) : ( n4086 ) ;
assign n4088 =  ( n3358 ) ? ( bv_8_13_n194 ) : ( n4087 ) ;
assign n4089 =  ( n3356 ) ? ( bv_8_191_n246 ) : ( n4088 ) ;
assign n4090 =  ( n3354 ) ? ( bv_8_230_n103 ) : ( n4089 ) ;
assign n4091 =  ( n3352 ) ? ( bv_8_66_n466 ) : ( n4090 ) ;
assign n4092 =  ( n3350 ) ? ( bv_8_104_n520 ) : ( n4091 ) ;
assign n4093 =  ( n3348 ) ? ( bv_8_65_n623 ) : ( n4092 ) ;
assign n4094 =  ( n3346 ) ? ( bv_8_153_n140 ) : ( n4093 ) ;
assign n4095 =  ( n3344 ) ? ( bv_8_45_n97 ) : ( n4094 ) ;
assign n4096 =  ( n3342 ) ? ( bv_8_15_n190 ) : ( n4095 ) ;
assign n4097 =  ( n3340 ) ? ( bv_8_176_n299 ) : ( n4096 ) ;
assign n4098 =  ( n3338 ) ? ( bv_8_84_n386 ) : ( n4097 ) ;
assign n4099 =  ( n3336 ) ? ( bv_8_187_n260 ) : ( n4098 ) ;
assign n4100 =  ( n3334 ) ? ( bv_8_22_n357 ) : ( n4099 ) ;
assign n4101 =  ( n3332 ) ^ ( n4100 )  ;
assign n4102 = key[127:120] ;
assign n4103 =  ( n4101 ) ^ ( n4102 )  ;
assign n4104 = state_in[127:120] ;
assign n4105 =  ( n4104 ) == ( bv_8_255_n3 )  ;
assign n4106 = state_in[127:120] ;
assign n4107 =  ( n4106 ) == ( bv_8_254_n7 )  ;
assign n4108 = state_in[127:120] ;
assign n4109 =  ( n4108 ) == ( bv_8_253_n11 )  ;
assign n4110 = state_in[127:120] ;
assign n4111 =  ( n4110 ) == ( bv_8_252_n15 )  ;
assign n4112 = state_in[127:120] ;
assign n4113 =  ( n4112 ) == ( bv_8_251_n19 )  ;
assign n4114 = state_in[127:120] ;
assign n4115 =  ( n4114 ) == ( bv_8_250_n23 )  ;
assign n4116 = state_in[127:120] ;
assign n4117 =  ( n4116 ) == ( bv_8_249_n27 )  ;
assign n4118 = state_in[127:120] ;
assign n4119 =  ( n4118 ) == ( bv_8_248_n31 )  ;
assign n4120 = state_in[127:120] ;
assign n4121 =  ( n4120 ) == ( bv_8_247_n35 )  ;
assign n4122 = state_in[127:120] ;
assign n4123 =  ( n4122 ) == ( bv_8_246_n39 )  ;
assign n4124 = state_in[127:120] ;
assign n4125 =  ( n4124 ) == ( bv_8_245_n43 )  ;
assign n4126 = state_in[127:120] ;
assign n4127 =  ( n4126 ) == ( bv_8_244_n47 )  ;
assign n4128 = state_in[127:120] ;
assign n4129 =  ( n4128 ) == ( bv_8_243_n51 )  ;
assign n4130 = state_in[127:120] ;
assign n4131 =  ( n4130 ) == ( bv_8_242_n55 )  ;
assign n4132 = state_in[127:120] ;
assign n4133 =  ( n4132 ) == ( bv_8_241_n59 )  ;
assign n4134 = state_in[127:120] ;
assign n4135 =  ( n4134 ) == ( bv_8_240_n63 )  ;
assign n4136 = state_in[127:120] ;
assign n4137 =  ( n4136 ) == ( bv_8_239_n67 )  ;
assign n4138 = state_in[127:120] ;
assign n4139 =  ( n4138 ) == ( bv_8_238_n71 )  ;
assign n4140 = state_in[127:120] ;
assign n4141 =  ( n4140 ) == ( bv_8_237_n75 )  ;
assign n4142 = state_in[127:120] ;
assign n4143 =  ( n4142 ) == ( bv_8_236_n79 )  ;
assign n4144 = state_in[127:120] ;
assign n4145 =  ( n4144 ) == ( bv_8_235_n83 )  ;
assign n4146 = state_in[127:120] ;
assign n4147 =  ( n4146 ) == ( bv_8_234_n87 )  ;
assign n4148 = state_in[127:120] ;
assign n4149 =  ( n4148 ) == ( bv_8_233_n91 )  ;
assign n4150 = state_in[127:120] ;
assign n4151 =  ( n4150 ) == ( bv_8_232_n95 )  ;
assign n4152 = state_in[127:120] ;
assign n4153 =  ( n4152 ) == ( bv_8_231_n99 )  ;
assign n4154 = state_in[127:120] ;
assign n4155 =  ( n4154 ) == ( bv_8_230_n103 )  ;
assign n4156 = state_in[127:120] ;
assign n4157 =  ( n4156 ) == ( bv_8_229_n107 )  ;
assign n4158 = state_in[127:120] ;
assign n4159 =  ( n4158 ) == ( bv_8_228_n111 )  ;
assign n4160 = state_in[127:120] ;
assign n4161 =  ( n4160 ) == ( bv_8_227_n115 )  ;
assign n4162 = state_in[127:120] ;
assign n4163 =  ( n4162 ) == ( bv_8_226_n119 )  ;
assign n4164 = state_in[127:120] ;
assign n4165 =  ( n4164 ) == ( bv_8_225_n123 )  ;
assign n4166 = state_in[127:120] ;
assign n4167 =  ( n4166 ) == ( bv_8_224_n126 )  ;
assign n4168 = state_in[127:120] ;
assign n4169 =  ( n4168 ) == ( bv_8_223_n130 )  ;
assign n4170 = state_in[127:120] ;
assign n4171 =  ( n4170 ) == ( bv_8_222_n134 )  ;
assign n4172 = state_in[127:120] ;
assign n4173 =  ( n4172 ) == ( bv_8_221_n138 )  ;
assign n4174 = state_in[127:120] ;
assign n4175 =  ( n4174 ) == ( bv_8_220_n142 )  ;
assign n4176 = state_in[127:120] ;
assign n4177 =  ( n4176 ) == ( bv_8_219_n146 )  ;
assign n4178 = state_in[127:120] ;
assign n4179 =  ( n4178 ) == ( bv_8_218_n150 )  ;
assign n4180 = state_in[127:120] ;
assign n4181 =  ( n4180 ) == ( bv_8_217_n128 )  ;
assign n4182 = state_in[127:120] ;
assign n4183 =  ( n4182 ) == ( bv_8_216_n157 )  ;
assign n4184 = state_in[127:120] ;
assign n4185 =  ( n4184 ) == ( bv_8_215_n45 )  ;
assign n4186 = state_in[127:120] ;
assign n4187 =  ( n4186 ) == ( bv_8_214_n164 )  ;
assign n4188 = state_in[127:120] ;
assign n4189 =  ( n4188 ) == ( bv_8_213_n167 )  ;
assign n4190 = state_in[127:120] ;
assign n4191 =  ( n4190 ) == ( bv_8_212_n171 )  ;
assign n4192 = state_in[127:120] ;
assign n4193 =  ( n4192 ) == ( bv_8_211_n175 )  ;
assign n4194 = state_in[127:120] ;
assign n4195 =  ( n4194 ) == ( bv_8_210_n113 )  ;
assign n4196 = state_in[127:120] ;
assign n4197 =  ( n4196 ) == ( bv_8_209_n182 )  ;
assign n4198 = state_in[127:120] ;
assign n4199 =  ( n4198 ) == ( bv_8_208_n37 )  ;
assign n4200 = state_in[127:120] ;
assign n4201 =  ( n4200 ) == ( bv_8_207_n188 )  ;
assign n4202 = state_in[127:120] ;
assign n4203 =  ( n4202 ) == ( bv_8_206_n192 )  ;
assign n4204 = state_in[127:120] ;
assign n4205 =  ( n4204 ) == ( bv_8_205_n196 )  ;
assign n4206 = state_in[127:120] ;
assign n4207 =  ( n4206 ) == ( bv_8_204_n177 )  ;
assign n4208 = state_in[127:120] ;
assign n4209 =  ( n4208 ) == ( bv_8_203_n203 )  ;
assign n4210 = state_in[127:120] ;
assign n4211 =  ( n4210 ) == ( bv_8_202_n207 )  ;
assign n4212 = state_in[127:120] ;
assign n4213 =  ( n4212 ) == ( bv_8_201_n85 )  ;
assign n4214 = state_in[127:120] ;
assign n4215 =  ( n4214 ) == ( bv_8_200_n213 )  ;
assign n4216 = state_in[127:120] ;
assign n4217 =  ( n4216 ) == ( bv_8_199_n216 )  ;
assign n4218 = state_in[127:120] ;
assign n4219 =  ( n4218 ) == ( bv_8_198_n220 )  ;
assign n4220 = state_in[127:120] ;
assign n4221 =  ( n4220 ) == ( bv_8_197_n224 )  ;
assign n4222 = state_in[127:120] ;
assign n4223 =  ( n4222 ) == ( bv_8_196_n228 )  ;
assign n4224 = state_in[127:120] ;
assign n4225 =  ( n4224 ) == ( bv_8_195_n232 )  ;
assign n4226 = state_in[127:120] ;
assign n4227 =  ( n4226 ) == ( bv_8_194_n159 )  ;
assign n4228 = state_in[127:120] ;
assign n4229 =  ( n4228 ) == ( bv_8_193_n239 )  ;
assign n4230 = state_in[127:120] ;
assign n4231 =  ( n4230 ) == ( bv_8_192_n242 )  ;
assign n4232 = state_in[127:120] ;
assign n4233 =  ( n4232 ) == ( bv_8_191_n246 )  ;
assign n4234 = state_in[127:120] ;
assign n4235 =  ( n4234 ) == ( bv_8_190_n250 )  ;
assign n4236 = state_in[127:120] ;
assign n4237 =  ( n4236 ) == ( bv_8_189_n254 )  ;
assign n4238 = state_in[127:120] ;
assign n4239 =  ( n4238 ) == ( bv_8_188_n257 )  ;
assign n4240 = state_in[127:120] ;
assign n4241 =  ( n4240 ) == ( bv_8_187_n260 )  ;
assign n4242 = state_in[127:120] ;
assign n4243 =  ( n4242 ) == ( bv_8_186_n263 )  ;
assign n4244 = state_in[127:120] ;
assign n4245 =  ( n4244 ) == ( bv_8_185_n266 )  ;
assign n4246 = state_in[127:120] ;
assign n4247 =  ( n4246 ) == ( bv_8_184_n270 )  ;
assign n4248 = state_in[127:120] ;
assign n4249 =  ( n4248 ) == ( bv_8_183_n273 )  ;
assign n4250 = state_in[127:120] ;
assign n4251 =  ( n4250 ) == ( bv_8_182_n277 )  ;
assign n4252 = state_in[127:120] ;
assign n4253 =  ( n4252 ) == ( bv_8_181_n281 )  ;
assign n4254 = state_in[127:120] ;
assign n4255 =  ( n4254 ) == ( bv_8_180_n285 )  ;
assign n4256 = state_in[127:120] ;
assign n4257 =  ( n4256 ) == ( bv_8_179_n289 )  ;
assign n4258 = state_in[127:120] ;
assign n4259 =  ( n4258 ) == ( bv_8_178_n292 )  ;
assign n4260 = state_in[127:120] ;
assign n4261 =  ( n4260 ) == ( bv_8_177_n283 )  ;
assign n4262 = state_in[127:120] ;
assign n4263 =  ( n4262 ) == ( bv_8_176_n299 )  ;
assign n4264 = state_in[127:120] ;
assign n4265 =  ( n4264 ) == ( bv_8_175_n302 )  ;
assign n4266 = state_in[127:120] ;
assign n4267 =  ( n4266 ) == ( bv_8_174_n152 )  ;
assign n4268 = state_in[127:120] ;
assign n4269 =  ( n4268 ) == ( bv_8_173_n307 )  ;
assign n4270 = state_in[127:120] ;
assign n4271 =  ( n4270 ) == ( bv_8_172_n268 )  ;
assign n4272 = state_in[127:120] ;
assign n4273 =  ( n4272 ) == ( bv_8_171_n314 )  ;
assign n4274 = state_in[127:120] ;
assign n4275 =  ( n4274 ) == ( bv_8_170_n77 )  ;
assign n4276 = state_in[127:120] ;
assign n4277 =  ( n4276 ) == ( bv_8_169_n109 )  ;
assign n4278 = state_in[127:120] ;
assign n4279 =  ( n4278 ) == ( bv_8_168_n13 )  ;
assign n4280 = state_in[127:120] ;
assign n4281 =  ( n4280 ) == ( bv_8_167_n325 )  ;
assign n4282 = state_in[127:120] ;
assign n4283 =  ( n4282 ) == ( bv_8_166_n328 )  ;
assign n4284 = state_in[127:120] ;
assign n4285 =  ( n4284 ) == ( bv_8_165_n69 )  ;
assign n4286 = state_in[127:120] ;
assign n4287 =  ( n4286 ) == ( bv_8_164_n335 )  ;
assign n4288 = state_in[127:120] ;
assign n4289 =  ( n4288 ) == ( bv_8_163_n339 )  ;
assign n4290 = state_in[127:120] ;
assign n4291 =  ( n4290 ) == ( bv_8_162_n343 )  ;
assign n4292 = state_in[127:120] ;
assign n4293 =  ( n4292 ) == ( bv_8_161_n211 )  ;
assign n4294 = state_in[127:120] ;
assign n4295 =  ( n4294 ) == ( bv_8_160_n350 )  ;
assign n4296 = state_in[127:120] ;
assign n4297 =  ( n4296 ) == ( bv_8_159_n323 )  ;
assign n4298 = state_in[127:120] ;
assign n4299 =  ( n4298 ) == ( bv_8_158_n355 )  ;
assign n4300 = state_in[127:120] ;
assign n4301 =  ( n4300 ) == ( bv_8_157_n359 )  ;
assign n4302 = state_in[127:120] ;
assign n4303 =  ( n4302 ) == ( bv_8_156_n279 )  ;
assign n4304 = state_in[127:120] ;
assign n4305 =  ( n4304 ) == ( bv_8_155_n364 )  ;
assign n4306 = state_in[127:120] ;
assign n4307 =  ( n4306 ) == ( bv_8_154_n368 )  ;
assign n4308 = state_in[127:120] ;
assign n4309 =  ( n4308 ) == ( bv_8_153_n140 )  ;
assign n4310 = state_in[127:120] ;
assign n4311 =  ( n4310 ) == ( bv_8_152_n374 )  ;
assign n4312 = state_in[127:120] ;
assign n4313 =  ( n4312 ) == ( bv_8_151_n218 )  ;
assign n4314 = state_in[127:120] ;
assign n4315 =  ( n4314 ) == ( bv_8_150_n201 )  ;
assign n4316 = state_in[127:120] ;
assign n4317 =  ( n4316 ) == ( bv_8_149_n384 )  ;
assign n4318 = state_in[127:120] ;
assign n4319 =  ( n4318 ) == ( bv_8_148_n388 )  ;
assign n4320 = state_in[127:120] ;
assign n4321 =  ( n4320 ) == ( bv_8_147_n392 )  ;
assign n4322 = state_in[127:120] ;
assign n4323 =  ( n4322 ) == ( bv_8_146_n337 )  ;
assign n4324 = state_in[127:120] ;
assign n4325 =  ( n4324 ) == ( bv_8_145_n397 )  ;
assign n4326 = state_in[127:120] ;
assign n4327 =  ( n4326 ) == ( bv_8_144_n173 )  ;
assign n4328 = state_in[127:120] ;
assign n4329 =  ( n4328 ) == ( bv_8_143_n403 )  ;
assign n4330 = state_in[127:120] ;
assign n4331 =  ( n4330 ) == ( bv_8_142_n406 )  ;
assign n4332 = state_in[127:120] ;
assign n4333 =  ( n4332 ) == ( bv_8_141_n410 )  ;
assign n4334 = state_in[127:120] ;
assign n4335 =  ( n4334 ) == ( bv_8_140_n376 )  ;
assign n4336 = state_in[127:120] ;
assign n4337 =  ( n4336 ) == ( bv_8_139_n297 )  ;
assign n4338 = state_in[127:120] ;
assign n4339 =  ( n4338 ) == ( bv_8_138_n418 )  ;
assign n4340 = state_in[127:120] ;
assign n4341 =  ( n4340 ) == ( bv_8_137_n421 )  ;
assign n4342 = state_in[127:120] ;
assign n4343 =  ( n4342 ) == ( bv_8_136_n425 )  ;
assign n4344 = state_in[127:120] ;
assign n4345 =  ( n4344 ) == ( bv_8_135_n81 )  ;
assign n4346 = state_in[127:120] ;
assign n4347 =  ( n4346 ) == ( bv_8_134_n431 )  ;
assign n4348 = state_in[127:120] ;
assign n4349 =  ( n4348 ) == ( bv_8_133_n434 )  ;
assign n4350 = state_in[127:120] ;
assign n4351 =  ( n4350 ) == ( bv_8_132_n41 )  ;
assign n4352 = state_in[127:120] ;
assign n4353 =  ( n4352 ) == ( bv_8_131_n440 )  ;
assign n4354 = state_in[127:120] ;
assign n4355 =  ( n4354 ) == ( bv_8_130_n33 )  ;
assign n4356 = state_in[127:120] ;
assign n4357 =  ( n4356 ) == ( bv_8_129_n446 )  ;
assign n4358 = state_in[127:120] ;
assign n4359 =  ( n4358 ) == ( bv_8_128_n450 )  ;
assign n4360 = state_in[127:120] ;
assign n4361 =  ( n4360 ) == ( bv_8_127_n453 )  ;
assign n4362 = state_in[127:120] ;
assign n4363 =  ( n4362 ) == ( bv_8_126_n456 )  ;
assign n4364 = state_in[127:120] ;
assign n4365 =  ( n4364 ) == ( bv_8_125_n459 )  ;
assign n4366 = state_in[127:120] ;
assign n4367 =  ( n4366 ) == ( bv_8_124_n184 )  ;
assign n4368 = state_in[127:120] ;
assign n4369 =  ( n4368 ) == ( bv_8_123_n17 )  ;
assign n4370 = state_in[127:120] ;
assign n4371 =  ( n4370 ) == ( bv_8_122_n416 )  ;
assign n4372 = state_in[127:120] ;
assign n4373 =  ( n4372 ) == ( bv_8_121_n470 )  ;
assign n4374 = state_in[127:120] ;
assign n4375 =  ( n4374 ) == ( bv_8_120_n474 )  ;
assign n4376 = state_in[127:120] ;
assign n4377 =  ( n4376 ) == ( bv_8_119_n472 )  ;
assign n4378 = state_in[127:120] ;
assign n4379 =  ( n4378 ) == ( bv_8_118_n480 )  ;
assign n4380 = state_in[127:120] ;
assign n4381 =  ( n4380 ) == ( bv_8_117_n484 )  ;
assign n4382 = state_in[127:120] ;
assign n4383 =  ( n4382 ) == ( bv_8_116_n345 )  ;
assign n4384 = state_in[127:120] ;
assign n4385 =  ( n4384 ) == ( bv_8_115_n222 )  ;
assign n4386 = state_in[127:120] ;
assign n4387 =  ( n4386 ) == ( bv_8_114_n494 )  ;
assign n4388 = state_in[127:120] ;
assign n4389 =  ( n4388 ) == ( bv_8_113_n180 )  ;
assign n4390 = state_in[127:120] ;
assign n4391 =  ( n4390 ) == ( bv_8_112_n482 )  ;
assign n4392 = state_in[127:120] ;
assign n4393 =  ( n4392 ) == ( bv_8_111_n244 )  ;
assign n4394 = state_in[127:120] ;
assign n4395 =  ( n4394 ) == ( bv_8_110_n294 )  ;
assign n4396 = state_in[127:120] ;
assign n4397 =  ( n4396 ) == ( bv_8_109_n9 )  ;
assign n4398 = state_in[127:120] ;
assign n4399 =  ( n4398 ) == ( bv_8_108_n510 )  ;
assign n4400 = state_in[127:120] ;
assign n4401 =  ( n4400 ) == ( bv_8_107_n370 )  ;
assign n4402 = state_in[127:120] ;
assign n4403 =  ( n4402 ) == ( bv_8_106_n155 )  ;
assign n4404 = state_in[127:120] ;
assign n4405 =  ( n4404 ) == ( bv_8_105_n148 )  ;
assign n4406 = state_in[127:120] ;
assign n4407 =  ( n4406 ) == ( bv_8_104_n520 )  ;
assign n4408 = state_in[127:120] ;
assign n4409 =  ( n4408 ) == ( bv_8_103_n523 )  ;
assign n4410 = state_in[127:120] ;
assign n4411 =  ( n4410 ) == ( bv_8_102_n527 )  ;
assign n4412 = state_in[127:120] ;
assign n4413 =  ( n4412 ) == ( bv_8_101_n49 )  ;
assign n4414 = state_in[127:120] ;
assign n4415 =  ( n4414 ) == ( bv_8_100_n348 )  ;
assign n4416 = state_in[127:120] ;
assign n4417 =  ( n4416 ) == ( bv_8_99_n476 )  ;
assign n4418 = state_in[127:120] ;
assign n4419 =  ( n4418 ) == ( bv_8_98_n536 )  ;
assign n4420 = state_in[127:120] ;
assign n4421 =  ( n4420 ) == ( bv_8_97_n198 )  ;
assign n4422 = state_in[127:120] ;
assign n4423 =  ( n4422 ) == ( bv_8_96_n542 )  ;
assign n4424 = state_in[127:120] ;
assign n4425 =  ( n4424 ) == ( bv_8_95_n545 )  ;
assign n4426 = state_in[127:120] ;
assign n4427 =  ( n4426 ) == ( bv_8_94_n548 )  ;
assign n4428 = state_in[127:120] ;
assign n4429 =  ( n4428 ) == ( bv_8_93_n498 )  ;
assign n4430 = state_in[127:120] ;
assign n4431 =  ( n4430 ) == ( bv_8_92_n234 )  ;
assign n4432 = state_in[127:120] ;
assign n4433 =  ( n4432 ) == ( bv_8_91_n555 )  ;
assign n4434 = state_in[127:120] ;
assign n4435 =  ( n4434 ) == ( bv_8_90_n25 )  ;
assign n4436 = state_in[127:120] ;
assign n4437 =  ( n4436 ) == ( bv_8_89_n61 )  ;
assign n4438 = state_in[127:120] ;
assign n4439 =  ( n4438 ) == ( bv_8_88_n562 )  ;
assign n4440 = state_in[127:120] ;
assign n4441 =  ( n4440 ) == ( bv_8_87_n226 )  ;
assign n4442 = state_in[127:120] ;
assign n4443 =  ( n4442 ) == ( bv_8_86_n567 )  ;
assign n4444 = state_in[127:120] ;
assign n4445 =  ( n4444 ) == ( bv_8_85_n423 )  ;
assign n4446 = state_in[127:120] ;
assign n4447 =  ( n4446 ) == ( bv_8_84_n386 )  ;
assign n4448 = state_in[127:120] ;
assign n4449 =  ( n4448 ) == ( bv_8_83_n575 )  ;
assign n4450 = state_in[127:120] ;
assign n4451 =  ( n4450 ) == ( bv_8_82_n578 )  ;
assign n4452 = state_in[127:120] ;
assign n4453 =  ( n4452 ) == ( bv_8_81_n582 )  ;
assign n4454 = state_in[127:120] ;
assign n4455 =  ( n4454 ) == ( bv_8_80_n73 )  ;
assign n4456 = state_in[127:120] ;
assign n4457 =  ( n4456 ) == ( bv_8_79_n538 )  ;
assign n4458 = state_in[127:120] ;
assign n4459 =  ( n4458 ) == ( bv_8_78_n590 )  ;
assign n4460 = state_in[127:120] ;
assign n4461 =  ( n4460 ) == ( bv_8_77_n593 )  ;
assign n4462 = state_in[127:120] ;
assign n4463 =  ( n4462 ) == ( bv_8_76_n596 )  ;
assign n4464 = state_in[127:120] ;
assign n4465 =  ( n4464 ) == ( bv_8_75_n503 )  ;
assign n4466 = state_in[127:120] ;
assign n4467 =  ( n4466 ) == ( bv_8_74_n237 )  ;
assign n4468 = state_in[127:120] ;
assign n4469 =  ( n4468 ) == ( bv_8_73_n275 )  ;
assign n4470 = state_in[127:120] ;
assign n4471 =  ( n4470 ) == ( bv_8_72_n330 )  ;
assign n4472 = state_in[127:120] ;
assign n4473 =  ( n4472 ) == ( bv_8_71_n252 )  ;
assign n4474 = state_in[127:120] ;
assign n4475 =  ( n4474 ) == ( bv_8_70_n609 )  ;
assign n4476 = state_in[127:120] ;
assign n4477 =  ( n4476 ) == ( bv_8_69_n612 )  ;
assign n4478 = state_in[127:120] ;
assign n4479 =  ( n4478 ) == ( bv_8_68_n390 )  ;
assign n4480 = state_in[127:120] ;
assign n4481 =  ( n4480 ) == ( bv_8_67_n318 )  ;
assign n4482 = state_in[127:120] ;
assign n4483 =  ( n4482 ) == ( bv_8_66_n466 )  ;
assign n4484 = state_in[127:120] ;
assign n4485 =  ( n4484 ) == ( bv_8_65_n623 )  ;
assign n4486 = state_in[127:120] ;
assign n4487 =  ( n4486 ) == ( bv_8_64_n573 )  ;
assign n4488 = state_in[127:120] ;
assign n4489 =  ( n4488 ) == ( bv_8_63_n489 )  ;
assign n4490 = state_in[127:120] ;
assign n4491 =  ( n4490 ) == ( bv_8_62_n205 )  ;
assign n4492 = state_in[127:120] ;
assign n4493 =  ( n4492 ) == ( bv_8_61_n634 )  ;
assign n4494 = state_in[127:120] ;
assign n4495 =  ( n4494 ) == ( bv_8_60_n93 )  ;
assign n4496 = state_in[127:120] ;
assign n4497 =  ( n4496 ) == ( bv_8_59_n382 )  ;
assign n4498 = state_in[127:120] ;
assign n4499 =  ( n4498 ) == ( bv_8_58_n136 )  ;
assign n4500 = state_in[127:120] ;
assign n4501 =  ( n4500 ) == ( bv_8_57_n312 )  ;
assign n4502 = state_in[127:120] ;
assign n4503 =  ( n4502 ) == ( bv_8_56_n230 )  ;
assign n4504 = state_in[127:120] ;
assign n4505 =  ( n4504 ) == ( bv_8_55_n650 )  ;
assign n4506 = state_in[127:120] ;
assign n4507 =  ( n4506 ) == ( bv_8_54_n616 )  ;
assign n4508 = state_in[127:120] ;
assign n4509 =  ( n4508 ) == ( bv_8_53_n436 )  ;
assign n4510 = state_in[127:120] ;
assign n4511 =  ( n4510 ) == ( bv_8_52_n619 )  ;
assign n4512 = state_in[127:120] ;
assign n4513 =  ( n4512 ) == ( bv_8_51_n101 )  ;
assign n4514 = state_in[127:120] ;
assign n4515 =  ( n4514 ) == ( bv_8_50_n408 )  ;
assign n4516 = state_in[127:120] ;
assign n4517 =  ( n4516 ) == ( bv_8_49_n309 )  ;
assign n4518 = state_in[127:120] ;
assign n4519 =  ( n4518 ) == ( bv_8_48_n660 )  ;
assign n4520 = state_in[127:120] ;
assign n4521 =  ( n4520 ) == ( bv_8_47_n652 )  ;
assign n4522 = state_in[127:120] ;
assign n4523 =  ( n4522 ) == ( bv_8_46_n429 )  ;
assign n4524 = state_in[127:120] ;
assign n4525 =  ( n4524 ) == ( bv_8_45_n97 )  ;
assign n4526 = state_in[127:120] ;
assign n4527 =  ( n4526 ) == ( bv_8_44_n5 )  ;
assign n4528 = state_in[127:120] ;
assign n4529 =  ( n4528 ) == ( bv_8_43_n121 )  ;
assign n4530 = state_in[127:120] ;
assign n4531 =  ( n4530 ) == ( bv_8_42_n672 )  ;
assign n4532 = state_in[127:120] ;
assign n4533 =  ( n4532 ) == ( bv_8_41_n29 )  ;
assign n4534 = state_in[127:120] ;
assign n4535 =  ( n4534 ) == ( bv_8_40_n366 )  ;
assign n4536 = state_in[127:120] ;
assign n4537 =  ( n4536 ) == ( bv_8_39_n132 )  ;
assign n4538 = state_in[127:120] ;
assign n4539 =  ( n4538 ) == ( bv_8_38_n444 )  ;
assign n4540 = state_in[127:120] ;
assign n4541 =  ( n4540 ) == ( bv_8_37_n506 )  ;
assign n4542 = state_in[127:120] ;
assign n4543 =  ( n4542 ) == ( bv_8_36_n645 )  ;
assign n4544 = state_in[127:120] ;
assign n4545 =  ( n4544 ) == ( bv_8_35_n696 )  ;
assign n4546 = state_in[127:120] ;
assign n4547 =  ( n4546 ) == ( bv_8_34_n117 )  ;
assign n4548 = state_in[127:120] ;
assign n4549 =  ( n4548 ) == ( bv_8_33_n486 )  ;
assign n4550 = state_in[127:120] ;
assign n4551 =  ( n4550 ) == ( bv_8_32_n463 )  ;
assign n4552 = state_in[127:120] ;
assign n4553 =  ( n4552 ) == ( bv_8_31_n705 )  ;
assign n4554 = state_in[127:120] ;
assign n4555 =  ( n4554 ) == ( bv_8_30_n21 )  ;
assign n4556 = state_in[127:120] ;
assign n4557 =  ( n4556 ) == ( bv_8_29_n625 )  ;
assign n4558 = state_in[127:120] ;
assign n4559 =  ( n4558 ) == ( bv_8_28_n162 )  ;
assign n4560 = state_in[127:120] ;
assign n4561 =  ( n4560 ) == ( bv_8_27_n642 )  ;
assign n4562 = state_in[127:120] ;
assign n4563 =  ( n4562 ) == ( bv_8_26_n53 )  ;
assign n4564 = state_in[127:120] ;
assign n4565 =  ( n4564 ) == ( bv_8_25_n399 )  ;
assign n4566 = state_in[127:120] ;
assign n4567 =  ( n4566 ) == ( bv_8_24_n448 )  ;
assign n4568 = state_in[127:120] ;
assign n4569 =  ( n4568 ) == ( bv_8_23_n144 )  ;
assign n4570 = state_in[127:120] ;
assign n4571 =  ( n4570 ) == ( bv_8_22_n357 )  ;
assign n4572 = state_in[127:120] ;
assign n4573 =  ( n4572 ) == ( bv_8_21_n89 )  ;
assign n4574 = state_in[127:120] ;
assign n4575 =  ( n4574 ) == ( bv_8_20_n341 )  ;
assign n4576 = state_in[127:120] ;
assign n4577 =  ( n4576 ) == ( bv_8_19_n588 )  ;
assign n4578 = state_in[127:120] ;
assign n4579 =  ( n4578 ) == ( bv_8_18_n628 )  ;
assign n4580 = state_in[127:120] ;
assign n4581 =  ( n4580 ) == ( bv_8_17_n525 )  ;
assign n4582 = state_in[127:120] ;
assign n4583 =  ( n4582 ) == ( bv_8_16_n248 )  ;
assign n4584 = state_in[127:120] ;
assign n4585 =  ( n4584 ) == ( bv_8_15_n190 )  ;
assign n4586 = state_in[127:120] ;
assign n4587 =  ( n4586 ) == ( bv_8_14_n648 )  ;
assign n4588 = state_in[127:120] ;
assign n4589 =  ( n4588 ) == ( bv_8_13_n194 )  ;
assign n4590 = state_in[127:120] ;
assign n4591 =  ( n4590 ) == ( bv_8_12_n333 )  ;
assign n4592 = state_in[127:120] ;
assign n4593 =  ( n4592 ) == ( bv_8_11_n379 )  ;
assign n4594 = state_in[127:120] ;
assign n4595 =  ( n4594 ) == ( bv_8_10_n655 )  ;
assign n4596 = state_in[127:120] ;
assign n4597 =  ( n4596 ) == ( bv_8_9_n57 )  ;
assign n4598 = state_in[127:120] ;
assign n4599 =  ( n4598 ) == ( bv_8_8_n669 )  ;
assign n4600 = state_in[127:120] ;
assign n4601 =  ( n4600 ) == ( bv_8_7_n105 )  ;
assign n4602 = state_in[127:120] ;
assign n4603 =  ( n4602 ) == ( bv_8_6_n169 )  ;
assign n4604 = state_in[127:120] ;
assign n4605 =  ( n4604 ) == ( bv_8_5_n492 )  ;
assign n4606 = state_in[127:120] ;
assign n4607 =  ( n4606 ) == ( bv_8_4_n516 )  ;
assign n4608 = state_in[127:120] ;
assign n4609 =  ( n4608 ) == ( bv_8_3_n65 )  ;
assign n4610 = state_in[127:120] ;
assign n4611 =  ( n4610 ) == ( bv_8_2_n751 )  ;
assign n4612 = state_in[127:120] ;
assign n4613 =  ( n4612 ) == ( bv_8_1_n287 )  ;
assign n4614 = state_in[127:120] ;
assign n4615 =  ( n4614 ) == ( bv_8_0_n580 )  ;
assign n4616 =  ( n4615 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n4617 =  ( n4613 ) ? ( bv_8_124_n184 ) : ( n4616 ) ;
assign n4618 =  ( n4611 ) ? ( bv_8_119_n472 ) : ( n4617 ) ;
assign n4619 =  ( n4609 ) ? ( bv_8_123_n17 ) : ( n4618 ) ;
assign n4620 =  ( n4607 ) ? ( bv_8_242_n55 ) : ( n4619 ) ;
assign n4621 =  ( n4605 ) ? ( bv_8_107_n370 ) : ( n4620 ) ;
assign n4622 =  ( n4603 ) ? ( bv_8_111_n244 ) : ( n4621 ) ;
assign n4623 =  ( n4601 ) ? ( bv_8_197_n224 ) : ( n4622 ) ;
assign n4624 =  ( n4599 ) ? ( bv_8_48_n660 ) : ( n4623 ) ;
assign n4625 =  ( n4597 ) ? ( bv_8_1_n287 ) : ( n4624 ) ;
assign n4626 =  ( n4595 ) ? ( bv_8_103_n523 ) : ( n4625 ) ;
assign n4627 =  ( n4593 ) ? ( bv_8_43_n121 ) : ( n4626 ) ;
assign n4628 =  ( n4591 ) ? ( bv_8_254_n7 ) : ( n4627 ) ;
assign n4629 =  ( n4589 ) ? ( bv_8_215_n45 ) : ( n4628 ) ;
assign n4630 =  ( n4587 ) ? ( bv_8_171_n314 ) : ( n4629 ) ;
assign n4631 =  ( n4585 ) ? ( bv_8_118_n480 ) : ( n4630 ) ;
assign n4632 =  ( n4583 ) ? ( bv_8_202_n207 ) : ( n4631 ) ;
assign n4633 =  ( n4581 ) ? ( bv_8_130_n33 ) : ( n4632 ) ;
assign n4634 =  ( n4579 ) ? ( bv_8_201_n85 ) : ( n4633 ) ;
assign n4635 =  ( n4577 ) ? ( bv_8_125_n459 ) : ( n4634 ) ;
assign n4636 =  ( n4575 ) ? ( bv_8_250_n23 ) : ( n4635 ) ;
assign n4637 =  ( n4573 ) ? ( bv_8_89_n61 ) : ( n4636 ) ;
assign n4638 =  ( n4571 ) ? ( bv_8_71_n252 ) : ( n4637 ) ;
assign n4639 =  ( n4569 ) ? ( bv_8_240_n63 ) : ( n4638 ) ;
assign n4640 =  ( n4567 ) ? ( bv_8_173_n307 ) : ( n4639 ) ;
assign n4641 =  ( n4565 ) ? ( bv_8_212_n171 ) : ( n4640 ) ;
assign n4642 =  ( n4563 ) ? ( bv_8_162_n343 ) : ( n4641 ) ;
assign n4643 =  ( n4561 ) ? ( bv_8_175_n302 ) : ( n4642 ) ;
assign n4644 =  ( n4559 ) ? ( bv_8_156_n279 ) : ( n4643 ) ;
assign n4645 =  ( n4557 ) ? ( bv_8_164_n335 ) : ( n4644 ) ;
assign n4646 =  ( n4555 ) ? ( bv_8_114_n494 ) : ( n4645 ) ;
assign n4647 =  ( n4553 ) ? ( bv_8_192_n242 ) : ( n4646 ) ;
assign n4648 =  ( n4551 ) ? ( bv_8_183_n273 ) : ( n4647 ) ;
assign n4649 =  ( n4549 ) ? ( bv_8_253_n11 ) : ( n4648 ) ;
assign n4650 =  ( n4547 ) ? ( bv_8_147_n392 ) : ( n4649 ) ;
assign n4651 =  ( n4545 ) ? ( bv_8_38_n444 ) : ( n4650 ) ;
assign n4652 =  ( n4543 ) ? ( bv_8_54_n616 ) : ( n4651 ) ;
assign n4653 =  ( n4541 ) ? ( bv_8_63_n489 ) : ( n4652 ) ;
assign n4654 =  ( n4539 ) ? ( bv_8_247_n35 ) : ( n4653 ) ;
assign n4655 =  ( n4537 ) ? ( bv_8_204_n177 ) : ( n4654 ) ;
assign n4656 =  ( n4535 ) ? ( bv_8_52_n619 ) : ( n4655 ) ;
assign n4657 =  ( n4533 ) ? ( bv_8_165_n69 ) : ( n4656 ) ;
assign n4658 =  ( n4531 ) ? ( bv_8_229_n107 ) : ( n4657 ) ;
assign n4659 =  ( n4529 ) ? ( bv_8_241_n59 ) : ( n4658 ) ;
assign n4660 =  ( n4527 ) ? ( bv_8_113_n180 ) : ( n4659 ) ;
assign n4661 =  ( n4525 ) ? ( bv_8_216_n157 ) : ( n4660 ) ;
assign n4662 =  ( n4523 ) ? ( bv_8_49_n309 ) : ( n4661 ) ;
assign n4663 =  ( n4521 ) ? ( bv_8_21_n89 ) : ( n4662 ) ;
assign n4664 =  ( n4519 ) ? ( bv_8_4_n516 ) : ( n4663 ) ;
assign n4665 =  ( n4517 ) ? ( bv_8_199_n216 ) : ( n4664 ) ;
assign n4666 =  ( n4515 ) ? ( bv_8_35_n696 ) : ( n4665 ) ;
assign n4667 =  ( n4513 ) ? ( bv_8_195_n232 ) : ( n4666 ) ;
assign n4668 =  ( n4511 ) ? ( bv_8_24_n448 ) : ( n4667 ) ;
assign n4669 =  ( n4509 ) ? ( bv_8_150_n201 ) : ( n4668 ) ;
assign n4670 =  ( n4507 ) ? ( bv_8_5_n492 ) : ( n4669 ) ;
assign n4671 =  ( n4505 ) ? ( bv_8_154_n368 ) : ( n4670 ) ;
assign n4672 =  ( n4503 ) ? ( bv_8_7_n105 ) : ( n4671 ) ;
assign n4673 =  ( n4501 ) ? ( bv_8_18_n628 ) : ( n4672 ) ;
assign n4674 =  ( n4499 ) ? ( bv_8_128_n450 ) : ( n4673 ) ;
assign n4675 =  ( n4497 ) ? ( bv_8_226_n119 ) : ( n4674 ) ;
assign n4676 =  ( n4495 ) ? ( bv_8_235_n83 ) : ( n4675 ) ;
assign n4677 =  ( n4493 ) ? ( bv_8_39_n132 ) : ( n4676 ) ;
assign n4678 =  ( n4491 ) ? ( bv_8_178_n292 ) : ( n4677 ) ;
assign n4679 =  ( n4489 ) ? ( bv_8_117_n484 ) : ( n4678 ) ;
assign n4680 =  ( n4487 ) ? ( bv_8_9_n57 ) : ( n4679 ) ;
assign n4681 =  ( n4485 ) ? ( bv_8_131_n440 ) : ( n4680 ) ;
assign n4682 =  ( n4483 ) ? ( bv_8_44_n5 ) : ( n4681 ) ;
assign n4683 =  ( n4481 ) ? ( bv_8_26_n53 ) : ( n4682 ) ;
assign n4684 =  ( n4479 ) ? ( bv_8_27_n642 ) : ( n4683 ) ;
assign n4685 =  ( n4477 ) ? ( bv_8_110_n294 ) : ( n4684 ) ;
assign n4686 =  ( n4475 ) ? ( bv_8_90_n25 ) : ( n4685 ) ;
assign n4687 =  ( n4473 ) ? ( bv_8_160_n350 ) : ( n4686 ) ;
assign n4688 =  ( n4471 ) ? ( bv_8_82_n578 ) : ( n4687 ) ;
assign n4689 =  ( n4469 ) ? ( bv_8_59_n382 ) : ( n4688 ) ;
assign n4690 =  ( n4467 ) ? ( bv_8_214_n164 ) : ( n4689 ) ;
assign n4691 =  ( n4465 ) ? ( bv_8_179_n289 ) : ( n4690 ) ;
assign n4692 =  ( n4463 ) ? ( bv_8_41_n29 ) : ( n4691 ) ;
assign n4693 =  ( n4461 ) ? ( bv_8_227_n115 ) : ( n4692 ) ;
assign n4694 =  ( n4459 ) ? ( bv_8_47_n652 ) : ( n4693 ) ;
assign n4695 =  ( n4457 ) ? ( bv_8_132_n41 ) : ( n4694 ) ;
assign n4696 =  ( n4455 ) ? ( bv_8_83_n575 ) : ( n4695 ) ;
assign n4697 =  ( n4453 ) ? ( bv_8_209_n182 ) : ( n4696 ) ;
assign n4698 =  ( n4451 ) ? ( bv_8_0_n580 ) : ( n4697 ) ;
assign n4699 =  ( n4449 ) ? ( bv_8_237_n75 ) : ( n4698 ) ;
assign n4700 =  ( n4447 ) ? ( bv_8_32_n463 ) : ( n4699 ) ;
assign n4701 =  ( n4445 ) ? ( bv_8_252_n15 ) : ( n4700 ) ;
assign n4702 =  ( n4443 ) ? ( bv_8_177_n283 ) : ( n4701 ) ;
assign n4703 =  ( n4441 ) ? ( bv_8_91_n555 ) : ( n4702 ) ;
assign n4704 =  ( n4439 ) ? ( bv_8_106_n155 ) : ( n4703 ) ;
assign n4705 =  ( n4437 ) ? ( bv_8_203_n203 ) : ( n4704 ) ;
assign n4706 =  ( n4435 ) ? ( bv_8_190_n250 ) : ( n4705 ) ;
assign n4707 =  ( n4433 ) ? ( bv_8_57_n312 ) : ( n4706 ) ;
assign n4708 =  ( n4431 ) ? ( bv_8_74_n237 ) : ( n4707 ) ;
assign n4709 =  ( n4429 ) ? ( bv_8_76_n596 ) : ( n4708 ) ;
assign n4710 =  ( n4427 ) ? ( bv_8_88_n562 ) : ( n4709 ) ;
assign n4711 =  ( n4425 ) ? ( bv_8_207_n188 ) : ( n4710 ) ;
assign n4712 =  ( n4423 ) ? ( bv_8_208_n37 ) : ( n4711 ) ;
assign n4713 =  ( n4421 ) ? ( bv_8_239_n67 ) : ( n4712 ) ;
assign n4714 =  ( n4419 ) ? ( bv_8_170_n77 ) : ( n4713 ) ;
assign n4715 =  ( n4417 ) ? ( bv_8_251_n19 ) : ( n4714 ) ;
assign n4716 =  ( n4415 ) ? ( bv_8_67_n318 ) : ( n4715 ) ;
assign n4717 =  ( n4413 ) ? ( bv_8_77_n593 ) : ( n4716 ) ;
assign n4718 =  ( n4411 ) ? ( bv_8_51_n101 ) : ( n4717 ) ;
assign n4719 =  ( n4409 ) ? ( bv_8_133_n434 ) : ( n4718 ) ;
assign n4720 =  ( n4407 ) ? ( bv_8_69_n612 ) : ( n4719 ) ;
assign n4721 =  ( n4405 ) ? ( bv_8_249_n27 ) : ( n4720 ) ;
assign n4722 =  ( n4403 ) ? ( bv_8_2_n751 ) : ( n4721 ) ;
assign n4723 =  ( n4401 ) ? ( bv_8_127_n453 ) : ( n4722 ) ;
assign n4724 =  ( n4399 ) ? ( bv_8_80_n73 ) : ( n4723 ) ;
assign n4725 =  ( n4397 ) ? ( bv_8_60_n93 ) : ( n4724 ) ;
assign n4726 =  ( n4395 ) ? ( bv_8_159_n323 ) : ( n4725 ) ;
assign n4727 =  ( n4393 ) ? ( bv_8_168_n13 ) : ( n4726 ) ;
assign n4728 =  ( n4391 ) ? ( bv_8_81_n582 ) : ( n4727 ) ;
assign n4729 =  ( n4389 ) ? ( bv_8_163_n339 ) : ( n4728 ) ;
assign n4730 =  ( n4387 ) ? ( bv_8_64_n573 ) : ( n4729 ) ;
assign n4731 =  ( n4385 ) ? ( bv_8_143_n403 ) : ( n4730 ) ;
assign n4732 =  ( n4383 ) ? ( bv_8_146_n337 ) : ( n4731 ) ;
assign n4733 =  ( n4381 ) ? ( bv_8_157_n359 ) : ( n4732 ) ;
assign n4734 =  ( n4379 ) ? ( bv_8_56_n230 ) : ( n4733 ) ;
assign n4735 =  ( n4377 ) ? ( bv_8_245_n43 ) : ( n4734 ) ;
assign n4736 =  ( n4375 ) ? ( bv_8_188_n257 ) : ( n4735 ) ;
assign n4737 =  ( n4373 ) ? ( bv_8_182_n277 ) : ( n4736 ) ;
assign n4738 =  ( n4371 ) ? ( bv_8_218_n150 ) : ( n4737 ) ;
assign n4739 =  ( n4369 ) ? ( bv_8_33_n486 ) : ( n4738 ) ;
assign n4740 =  ( n4367 ) ? ( bv_8_16_n248 ) : ( n4739 ) ;
assign n4741 =  ( n4365 ) ? ( bv_8_255_n3 ) : ( n4740 ) ;
assign n4742 =  ( n4363 ) ? ( bv_8_243_n51 ) : ( n4741 ) ;
assign n4743 =  ( n4361 ) ? ( bv_8_210_n113 ) : ( n4742 ) ;
assign n4744 =  ( n4359 ) ? ( bv_8_205_n196 ) : ( n4743 ) ;
assign n4745 =  ( n4357 ) ? ( bv_8_12_n333 ) : ( n4744 ) ;
assign n4746 =  ( n4355 ) ? ( bv_8_19_n588 ) : ( n4745 ) ;
assign n4747 =  ( n4353 ) ? ( bv_8_236_n79 ) : ( n4746 ) ;
assign n4748 =  ( n4351 ) ? ( bv_8_95_n545 ) : ( n4747 ) ;
assign n4749 =  ( n4349 ) ? ( bv_8_151_n218 ) : ( n4748 ) ;
assign n4750 =  ( n4347 ) ? ( bv_8_68_n390 ) : ( n4749 ) ;
assign n4751 =  ( n4345 ) ? ( bv_8_23_n144 ) : ( n4750 ) ;
assign n4752 =  ( n4343 ) ? ( bv_8_196_n228 ) : ( n4751 ) ;
assign n4753 =  ( n4341 ) ? ( bv_8_167_n325 ) : ( n4752 ) ;
assign n4754 =  ( n4339 ) ? ( bv_8_126_n456 ) : ( n4753 ) ;
assign n4755 =  ( n4337 ) ? ( bv_8_61_n634 ) : ( n4754 ) ;
assign n4756 =  ( n4335 ) ? ( bv_8_100_n348 ) : ( n4755 ) ;
assign n4757 =  ( n4333 ) ? ( bv_8_93_n498 ) : ( n4756 ) ;
assign n4758 =  ( n4331 ) ? ( bv_8_25_n399 ) : ( n4757 ) ;
assign n4759 =  ( n4329 ) ? ( bv_8_115_n222 ) : ( n4758 ) ;
assign n4760 =  ( n4327 ) ? ( bv_8_96_n542 ) : ( n4759 ) ;
assign n4761 =  ( n4325 ) ? ( bv_8_129_n446 ) : ( n4760 ) ;
assign n4762 =  ( n4323 ) ? ( bv_8_79_n538 ) : ( n4761 ) ;
assign n4763 =  ( n4321 ) ? ( bv_8_220_n142 ) : ( n4762 ) ;
assign n4764 =  ( n4319 ) ? ( bv_8_34_n117 ) : ( n4763 ) ;
assign n4765 =  ( n4317 ) ? ( bv_8_42_n672 ) : ( n4764 ) ;
assign n4766 =  ( n4315 ) ? ( bv_8_144_n173 ) : ( n4765 ) ;
assign n4767 =  ( n4313 ) ? ( bv_8_136_n425 ) : ( n4766 ) ;
assign n4768 =  ( n4311 ) ? ( bv_8_70_n609 ) : ( n4767 ) ;
assign n4769 =  ( n4309 ) ? ( bv_8_238_n71 ) : ( n4768 ) ;
assign n4770 =  ( n4307 ) ? ( bv_8_184_n270 ) : ( n4769 ) ;
assign n4771 =  ( n4305 ) ? ( bv_8_20_n341 ) : ( n4770 ) ;
assign n4772 =  ( n4303 ) ? ( bv_8_222_n134 ) : ( n4771 ) ;
assign n4773 =  ( n4301 ) ? ( bv_8_94_n548 ) : ( n4772 ) ;
assign n4774 =  ( n4299 ) ? ( bv_8_11_n379 ) : ( n4773 ) ;
assign n4775 =  ( n4297 ) ? ( bv_8_219_n146 ) : ( n4774 ) ;
assign n4776 =  ( n4295 ) ? ( bv_8_224_n126 ) : ( n4775 ) ;
assign n4777 =  ( n4293 ) ? ( bv_8_50_n408 ) : ( n4776 ) ;
assign n4778 =  ( n4291 ) ? ( bv_8_58_n136 ) : ( n4777 ) ;
assign n4779 =  ( n4289 ) ? ( bv_8_10_n655 ) : ( n4778 ) ;
assign n4780 =  ( n4287 ) ? ( bv_8_73_n275 ) : ( n4779 ) ;
assign n4781 =  ( n4285 ) ? ( bv_8_6_n169 ) : ( n4780 ) ;
assign n4782 =  ( n4283 ) ? ( bv_8_36_n645 ) : ( n4781 ) ;
assign n4783 =  ( n4281 ) ? ( bv_8_92_n234 ) : ( n4782 ) ;
assign n4784 =  ( n4279 ) ? ( bv_8_194_n159 ) : ( n4783 ) ;
assign n4785 =  ( n4277 ) ? ( bv_8_211_n175 ) : ( n4784 ) ;
assign n4786 =  ( n4275 ) ? ( bv_8_172_n268 ) : ( n4785 ) ;
assign n4787 =  ( n4273 ) ? ( bv_8_98_n536 ) : ( n4786 ) ;
assign n4788 =  ( n4271 ) ? ( bv_8_145_n397 ) : ( n4787 ) ;
assign n4789 =  ( n4269 ) ? ( bv_8_149_n384 ) : ( n4788 ) ;
assign n4790 =  ( n4267 ) ? ( bv_8_228_n111 ) : ( n4789 ) ;
assign n4791 =  ( n4265 ) ? ( bv_8_121_n470 ) : ( n4790 ) ;
assign n4792 =  ( n4263 ) ? ( bv_8_231_n99 ) : ( n4791 ) ;
assign n4793 =  ( n4261 ) ? ( bv_8_200_n213 ) : ( n4792 ) ;
assign n4794 =  ( n4259 ) ? ( bv_8_55_n650 ) : ( n4793 ) ;
assign n4795 =  ( n4257 ) ? ( bv_8_109_n9 ) : ( n4794 ) ;
assign n4796 =  ( n4255 ) ? ( bv_8_141_n410 ) : ( n4795 ) ;
assign n4797 =  ( n4253 ) ? ( bv_8_213_n167 ) : ( n4796 ) ;
assign n4798 =  ( n4251 ) ? ( bv_8_78_n590 ) : ( n4797 ) ;
assign n4799 =  ( n4249 ) ? ( bv_8_169_n109 ) : ( n4798 ) ;
assign n4800 =  ( n4247 ) ? ( bv_8_108_n510 ) : ( n4799 ) ;
assign n4801 =  ( n4245 ) ? ( bv_8_86_n567 ) : ( n4800 ) ;
assign n4802 =  ( n4243 ) ? ( bv_8_244_n47 ) : ( n4801 ) ;
assign n4803 =  ( n4241 ) ? ( bv_8_234_n87 ) : ( n4802 ) ;
assign n4804 =  ( n4239 ) ? ( bv_8_101_n49 ) : ( n4803 ) ;
assign n4805 =  ( n4237 ) ? ( bv_8_122_n416 ) : ( n4804 ) ;
assign n4806 =  ( n4235 ) ? ( bv_8_174_n152 ) : ( n4805 ) ;
assign n4807 =  ( n4233 ) ? ( bv_8_8_n669 ) : ( n4806 ) ;
assign n4808 =  ( n4231 ) ? ( bv_8_186_n263 ) : ( n4807 ) ;
assign n4809 =  ( n4229 ) ? ( bv_8_120_n474 ) : ( n4808 ) ;
assign n4810 =  ( n4227 ) ? ( bv_8_37_n506 ) : ( n4809 ) ;
assign n4811 =  ( n4225 ) ? ( bv_8_46_n429 ) : ( n4810 ) ;
assign n4812 =  ( n4223 ) ? ( bv_8_28_n162 ) : ( n4811 ) ;
assign n4813 =  ( n4221 ) ? ( bv_8_166_n328 ) : ( n4812 ) ;
assign n4814 =  ( n4219 ) ? ( bv_8_180_n285 ) : ( n4813 ) ;
assign n4815 =  ( n4217 ) ? ( bv_8_198_n220 ) : ( n4814 ) ;
assign n4816 =  ( n4215 ) ? ( bv_8_232_n95 ) : ( n4815 ) ;
assign n4817 =  ( n4213 ) ? ( bv_8_221_n138 ) : ( n4816 ) ;
assign n4818 =  ( n4211 ) ? ( bv_8_116_n345 ) : ( n4817 ) ;
assign n4819 =  ( n4209 ) ? ( bv_8_31_n705 ) : ( n4818 ) ;
assign n4820 =  ( n4207 ) ? ( bv_8_75_n503 ) : ( n4819 ) ;
assign n4821 =  ( n4205 ) ? ( bv_8_189_n254 ) : ( n4820 ) ;
assign n4822 =  ( n4203 ) ? ( bv_8_139_n297 ) : ( n4821 ) ;
assign n4823 =  ( n4201 ) ? ( bv_8_138_n418 ) : ( n4822 ) ;
assign n4824 =  ( n4199 ) ? ( bv_8_112_n482 ) : ( n4823 ) ;
assign n4825 =  ( n4197 ) ? ( bv_8_62_n205 ) : ( n4824 ) ;
assign n4826 =  ( n4195 ) ? ( bv_8_181_n281 ) : ( n4825 ) ;
assign n4827 =  ( n4193 ) ? ( bv_8_102_n527 ) : ( n4826 ) ;
assign n4828 =  ( n4191 ) ? ( bv_8_72_n330 ) : ( n4827 ) ;
assign n4829 =  ( n4189 ) ? ( bv_8_3_n65 ) : ( n4828 ) ;
assign n4830 =  ( n4187 ) ? ( bv_8_246_n39 ) : ( n4829 ) ;
assign n4831 =  ( n4185 ) ? ( bv_8_14_n648 ) : ( n4830 ) ;
assign n4832 =  ( n4183 ) ? ( bv_8_97_n198 ) : ( n4831 ) ;
assign n4833 =  ( n4181 ) ? ( bv_8_53_n436 ) : ( n4832 ) ;
assign n4834 =  ( n4179 ) ? ( bv_8_87_n226 ) : ( n4833 ) ;
assign n4835 =  ( n4177 ) ? ( bv_8_185_n266 ) : ( n4834 ) ;
assign n4836 =  ( n4175 ) ? ( bv_8_134_n431 ) : ( n4835 ) ;
assign n4837 =  ( n4173 ) ? ( bv_8_193_n239 ) : ( n4836 ) ;
assign n4838 =  ( n4171 ) ? ( bv_8_29_n625 ) : ( n4837 ) ;
assign n4839 =  ( n4169 ) ? ( bv_8_158_n355 ) : ( n4838 ) ;
assign n4840 =  ( n4167 ) ? ( bv_8_225_n123 ) : ( n4839 ) ;
assign n4841 =  ( n4165 ) ? ( bv_8_248_n31 ) : ( n4840 ) ;
assign n4842 =  ( n4163 ) ? ( bv_8_152_n374 ) : ( n4841 ) ;
assign n4843 =  ( n4161 ) ? ( bv_8_17_n525 ) : ( n4842 ) ;
assign n4844 =  ( n4159 ) ? ( bv_8_105_n148 ) : ( n4843 ) ;
assign n4845 =  ( n4157 ) ? ( bv_8_217_n128 ) : ( n4844 ) ;
assign n4846 =  ( n4155 ) ? ( bv_8_142_n406 ) : ( n4845 ) ;
assign n4847 =  ( n4153 ) ? ( bv_8_148_n388 ) : ( n4846 ) ;
assign n4848 =  ( n4151 ) ? ( bv_8_155_n364 ) : ( n4847 ) ;
assign n4849 =  ( n4149 ) ? ( bv_8_30_n21 ) : ( n4848 ) ;
assign n4850 =  ( n4147 ) ? ( bv_8_135_n81 ) : ( n4849 ) ;
assign n4851 =  ( n4145 ) ? ( bv_8_233_n91 ) : ( n4850 ) ;
assign n4852 =  ( n4143 ) ? ( bv_8_206_n192 ) : ( n4851 ) ;
assign n4853 =  ( n4141 ) ? ( bv_8_85_n423 ) : ( n4852 ) ;
assign n4854 =  ( n4139 ) ? ( bv_8_40_n366 ) : ( n4853 ) ;
assign n4855 =  ( n4137 ) ? ( bv_8_223_n130 ) : ( n4854 ) ;
assign n4856 =  ( n4135 ) ? ( bv_8_140_n376 ) : ( n4855 ) ;
assign n4857 =  ( n4133 ) ? ( bv_8_161_n211 ) : ( n4856 ) ;
assign n4858 =  ( n4131 ) ? ( bv_8_137_n421 ) : ( n4857 ) ;
assign n4859 =  ( n4129 ) ? ( bv_8_13_n194 ) : ( n4858 ) ;
assign n4860 =  ( n4127 ) ? ( bv_8_191_n246 ) : ( n4859 ) ;
assign n4861 =  ( n4125 ) ? ( bv_8_230_n103 ) : ( n4860 ) ;
assign n4862 =  ( n4123 ) ? ( bv_8_66_n466 ) : ( n4861 ) ;
assign n4863 =  ( n4121 ) ? ( bv_8_104_n520 ) : ( n4862 ) ;
assign n4864 =  ( n4119 ) ? ( bv_8_65_n623 ) : ( n4863 ) ;
assign n4865 =  ( n4117 ) ? ( bv_8_153_n140 ) : ( n4864 ) ;
assign n4866 =  ( n4115 ) ? ( bv_8_45_n97 ) : ( n4865 ) ;
assign n4867 =  ( n4113 ) ? ( bv_8_15_n190 ) : ( n4866 ) ;
assign n4868 =  ( n4111 ) ? ( bv_8_176_n299 ) : ( n4867 ) ;
assign n4869 =  ( n4109 ) ? ( bv_8_84_n386 ) : ( n4868 ) ;
assign n4870 =  ( n4107 ) ? ( bv_8_187_n260 ) : ( n4869 ) ;
assign n4871 =  ( n4105 ) ? ( bv_8_22_n357 ) : ( n4870 ) ;
assign n4872 =  ( n4871 ) ^ ( n2562 )  ;
assign n4873 =  ( n4872 ) ^ ( n3331 )  ;
assign n4874 = state_in[47:40] ;
assign n4875 =  ( n4874 ) == ( bv_8_255_n3 )  ;
assign n4876 = state_in[47:40] ;
assign n4877 =  ( n4876 ) == ( bv_8_254_n7 )  ;
assign n4878 = state_in[47:40] ;
assign n4879 =  ( n4878 ) == ( bv_8_253_n11 )  ;
assign n4880 = state_in[47:40] ;
assign n4881 =  ( n4880 ) == ( bv_8_252_n15 )  ;
assign n4882 = state_in[47:40] ;
assign n4883 =  ( n4882 ) == ( bv_8_251_n19 )  ;
assign n4884 = state_in[47:40] ;
assign n4885 =  ( n4884 ) == ( bv_8_250_n23 )  ;
assign n4886 = state_in[47:40] ;
assign n4887 =  ( n4886 ) == ( bv_8_249_n27 )  ;
assign n4888 = state_in[47:40] ;
assign n4889 =  ( n4888 ) == ( bv_8_248_n31 )  ;
assign n4890 = state_in[47:40] ;
assign n4891 =  ( n4890 ) == ( bv_8_247_n35 )  ;
assign n4892 = state_in[47:40] ;
assign n4893 =  ( n4892 ) == ( bv_8_246_n39 )  ;
assign n4894 = state_in[47:40] ;
assign n4895 =  ( n4894 ) == ( bv_8_245_n43 )  ;
assign n4896 = state_in[47:40] ;
assign n4897 =  ( n4896 ) == ( bv_8_244_n47 )  ;
assign n4898 = state_in[47:40] ;
assign n4899 =  ( n4898 ) == ( bv_8_243_n51 )  ;
assign n4900 = state_in[47:40] ;
assign n4901 =  ( n4900 ) == ( bv_8_242_n55 )  ;
assign n4902 = state_in[47:40] ;
assign n4903 =  ( n4902 ) == ( bv_8_241_n59 )  ;
assign n4904 = state_in[47:40] ;
assign n4905 =  ( n4904 ) == ( bv_8_240_n63 )  ;
assign n4906 = state_in[47:40] ;
assign n4907 =  ( n4906 ) == ( bv_8_239_n67 )  ;
assign n4908 = state_in[47:40] ;
assign n4909 =  ( n4908 ) == ( bv_8_238_n71 )  ;
assign n4910 = state_in[47:40] ;
assign n4911 =  ( n4910 ) == ( bv_8_237_n75 )  ;
assign n4912 = state_in[47:40] ;
assign n4913 =  ( n4912 ) == ( bv_8_236_n79 )  ;
assign n4914 = state_in[47:40] ;
assign n4915 =  ( n4914 ) == ( bv_8_235_n83 )  ;
assign n4916 = state_in[47:40] ;
assign n4917 =  ( n4916 ) == ( bv_8_234_n87 )  ;
assign n4918 = state_in[47:40] ;
assign n4919 =  ( n4918 ) == ( bv_8_233_n91 )  ;
assign n4920 = state_in[47:40] ;
assign n4921 =  ( n4920 ) == ( bv_8_232_n95 )  ;
assign n4922 = state_in[47:40] ;
assign n4923 =  ( n4922 ) == ( bv_8_231_n99 )  ;
assign n4924 = state_in[47:40] ;
assign n4925 =  ( n4924 ) == ( bv_8_230_n103 )  ;
assign n4926 = state_in[47:40] ;
assign n4927 =  ( n4926 ) == ( bv_8_229_n107 )  ;
assign n4928 = state_in[47:40] ;
assign n4929 =  ( n4928 ) == ( bv_8_228_n111 )  ;
assign n4930 = state_in[47:40] ;
assign n4931 =  ( n4930 ) == ( bv_8_227_n115 )  ;
assign n4932 = state_in[47:40] ;
assign n4933 =  ( n4932 ) == ( bv_8_226_n119 )  ;
assign n4934 = state_in[47:40] ;
assign n4935 =  ( n4934 ) == ( bv_8_225_n123 )  ;
assign n4936 = state_in[47:40] ;
assign n4937 =  ( n4936 ) == ( bv_8_224_n126 )  ;
assign n4938 = state_in[47:40] ;
assign n4939 =  ( n4938 ) == ( bv_8_223_n130 )  ;
assign n4940 = state_in[47:40] ;
assign n4941 =  ( n4940 ) == ( bv_8_222_n134 )  ;
assign n4942 = state_in[47:40] ;
assign n4943 =  ( n4942 ) == ( bv_8_221_n138 )  ;
assign n4944 = state_in[47:40] ;
assign n4945 =  ( n4944 ) == ( bv_8_220_n142 )  ;
assign n4946 = state_in[47:40] ;
assign n4947 =  ( n4946 ) == ( bv_8_219_n146 )  ;
assign n4948 = state_in[47:40] ;
assign n4949 =  ( n4948 ) == ( bv_8_218_n150 )  ;
assign n4950 = state_in[47:40] ;
assign n4951 =  ( n4950 ) == ( bv_8_217_n128 )  ;
assign n4952 = state_in[47:40] ;
assign n4953 =  ( n4952 ) == ( bv_8_216_n157 )  ;
assign n4954 = state_in[47:40] ;
assign n4955 =  ( n4954 ) == ( bv_8_215_n45 )  ;
assign n4956 = state_in[47:40] ;
assign n4957 =  ( n4956 ) == ( bv_8_214_n164 )  ;
assign n4958 = state_in[47:40] ;
assign n4959 =  ( n4958 ) == ( bv_8_213_n167 )  ;
assign n4960 = state_in[47:40] ;
assign n4961 =  ( n4960 ) == ( bv_8_212_n171 )  ;
assign n4962 = state_in[47:40] ;
assign n4963 =  ( n4962 ) == ( bv_8_211_n175 )  ;
assign n4964 = state_in[47:40] ;
assign n4965 =  ( n4964 ) == ( bv_8_210_n113 )  ;
assign n4966 = state_in[47:40] ;
assign n4967 =  ( n4966 ) == ( bv_8_209_n182 )  ;
assign n4968 = state_in[47:40] ;
assign n4969 =  ( n4968 ) == ( bv_8_208_n37 )  ;
assign n4970 = state_in[47:40] ;
assign n4971 =  ( n4970 ) == ( bv_8_207_n188 )  ;
assign n4972 = state_in[47:40] ;
assign n4973 =  ( n4972 ) == ( bv_8_206_n192 )  ;
assign n4974 = state_in[47:40] ;
assign n4975 =  ( n4974 ) == ( bv_8_205_n196 )  ;
assign n4976 = state_in[47:40] ;
assign n4977 =  ( n4976 ) == ( bv_8_204_n177 )  ;
assign n4978 = state_in[47:40] ;
assign n4979 =  ( n4978 ) == ( bv_8_203_n203 )  ;
assign n4980 = state_in[47:40] ;
assign n4981 =  ( n4980 ) == ( bv_8_202_n207 )  ;
assign n4982 = state_in[47:40] ;
assign n4983 =  ( n4982 ) == ( bv_8_201_n85 )  ;
assign n4984 = state_in[47:40] ;
assign n4985 =  ( n4984 ) == ( bv_8_200_n213 )  ;
assign n4986 = state_in[47:40] ;
assign n4987 =  ( n4986 ) == ( bv_8_199_n216 )  ;
assign n4988 = state_in[47:40] ;
assign n4989 =  ( n4988 ) == ( bv_8_198_n220 )  ;
assign n4990 = state_in[47:40] ;
assign n4991 =  ( n4990 ) == ( bv_8_197_n224 )  ;
assign n4992 = state_in[47:40] ;
assign n4993 =  ( n4992 ) == ( bv_8_196_n228 )  ;
assign n4994 = state_in[47:40] ;
assign n4995 =  ( n4994 ) == ( bv_8_195_n232 )  ;
assign n4996 = state_in[47:40] ;
assign n4997 =  ( n4996 ) == ( bv_8_194_n159 )  ;
assign n4998 = state_in[47:40] ;
assign n4999 =  ( n4998 ) == ( bv_8_193_n239 )  ;
assign n5000 = state_in[47:40] ;
assign n5001 =  ( n5000 ) == ( bv_8_192_n242 )  ;
assign n5002 = state_in[47:40] ;
assign n5003 =  ( n5002 ) == ( bv_8_191_n246 )  ;
assign n5004 = state_in[47:40] ;
assign n5005 =  ( n5004 ) == ( bv_8_190_n250 )  ;
assign n5006 = state_in[47:40] ;
assign n5007 =  ( n5006 ) == ( bv_8_189_n254 )  ;
assign n5008 = state_in[47:40] ;
assign n5009 =  ( n5008 ) == ( bv_8_188_n257 )  ;
assign n5010 = state_in[47:40] ;
assign n5011 =  ( n5010 ) == ( bv_8_187_n260 )  ;
assign n5012 = state_in[47:40] ;
assign n5013 =  ( n5012 ) == ( bv_8_186_n263 )  ;
assign n5014 = state_in[47:40] ;
assign n5015 =  ( n5014 ) == ( bv_8_185_n266 )  ;
assign n5016 = state_in[47:40] ;
assign n5017 =  ( n5016 ) == ( bv_8_184_n270 )  ;
assign n5018 = state_in[47:40] ;
assign n5019 =  ( n5018 ) == ( bv_8_183_n273 )  ;
assign n5020 = state_in[47:40] ;
assign n5021 =  ( n5020 ) == ( bv_8_182_n277 )  ;
assign n5022 = state_in[47:40] ;
assign n5023 =  ( n5022 ) == ( bv_8_181_n281 )  ;
assign n5024 = state_in[47:40] ;
assign n5025 =  ( n5024 ) == ( bv_8_180_n285 )  ;
assign n5026 = state_in[47:40] ;
assign n5027 =  ( n5026 ) == ( bv_8_179_n289 )  ;
assign n5028 = state_in[47:40] ;
assign n5029 =  ( n5028 ) == ( bv_8_178_n292 )  ;
assign n5030 = state_in[47:40] ;
assign n5031 =  ( n5030 ) == ( bv_8_177_n283 )  ;
assign n5032 = state_in[47:40] ;
assign n5033 =  ( n5032 ) == ( bv_8_176_n299 )  ;
assign n5034 = state_in[47:40] ;
assign n5035 =  ( n5034 ) == ( bv_8_175_n302 )  ;
assign n5036 = state_in[47:40] ;
assign n5037 =  ( n5036 ) == ( bv_8_174_n152 )  ;
assign n5038 = state_in[47:40] ;
assign n5039 =  ( n5038 ) == ( bv_8_173_n307 )  ;
assign n5040 = state_in[47:40] ;
assign n5041 =  ( n5040 ) == ( bv_8_172_n268 )  ;
assign n5042 = state_in[47:40] ;
assign n5043 =  ( n5042 ) == ( bv_8_171_n314 )  ;
assign n5044 = state_in[47:40] ;
assign n5045 =  ( n5044 ) == ( bv_8_170_n77 )  ;
assign n5046 = state_in[47:40] ;
assign n5047 =  ( n5046 ) == ( bv_8_169_n109 )  ;
assign n5048 = state_in[47:40] ;
assign n5049 =  ( n5048 ) == ( bv_8_168_n13 )  ;
assign n5050 = state_in[47:40] ;
assign n5051 =  ( n5050 ) == ( bv_8_167_n325 )  ;
assign n5052 = state_in[47:40] ;
assign n5053 =  ( n5052 ) == ( bv_8_166_n328 )  ;
assign n5054 = state_in[47:40] ;
assign n5055 =  ( n5054 ) == ( bv_8_165_n69 )  ;
assign n5056 = state_in[47:40] ;
assign n5057 =  ( n5056 ) == ( bv_8_164_n335 )  ;
assign n5058 = state_in[47:40] ;
assign n5059 =  ( n5058 ) == ( bv_8_163_n339 )  ;
assign n5060 = state_in[47:40] ;
assign n5061 =  ( n5060 ) == ( bv_8_162_n343 )  ;
assign n5062 = state_in[47:40] ;
assign n5063 =  ( n5062 ) == ( bv_8_161_n211 )  ;
assign n5064 = state_in[47:40] ;
assign n5065 =  ( n5064 ) == ( bv_8_160_n350 )  ;
assign n5066 = state_in[47:40] ;
assign n5067 =  ( n5066 ) == ( bv_8_159_n323 )  ;
assign n5068 = state_in[47:40] ;
assign n5069 =  ( n5068 ) == ( bv_8_158_n355 )  ;
assign n5070 = state_in[47:40] ;
assign n5071 =  ( n5070 ) == ( bv_8_157_n359 )  ;
assign n5072 = state_in[47:40] ;
assign n5073 =  ( n5072 ) == ( bv_8_156_n279 )  ;
assign n5074 = state_in[47:40] ;
assign n5075 =  ( n5074 ) == ( bv_8_155_n364 )  ;
assign n5076 = state_in[47:40] ;
assign n5077 =  ( n5076 ) == ( bv_8_154_n368 )  ;
assign n5078 = state_in[47:40] ;
assign n5079 =  ( n5078 ) == ( bv_8_153_n140 )  ;
assign n5080 = state_in[47:40] ;
assign n5081 =  ( n5080 ) == ( bv_8_152_n374 )  ;
assign n5082 = state_in[47:40] ;
assign n5083 =  ( n5082 ) == ( bv_8_151_n218 )  ;
assign n5084 = state_in[47:40] ;
assign n5085 =  ( n5084 ) == ( bv_8_150_n201 )  ;
assign n5086 = state_in[47:40] ;
assign n5087 =  ( n5086 ) == ( bv_8_149_n384 )  ;
assign n5088 = state_in[47:40] ;
assign n5089 =  ( n5088 ) == ( bv_8_148_n388 )  ;
assign n5090 = state_in[47:40] ;
assign n5091 =  ( n5090 ) == ( bv_8_147_n392 )  ;
assign n5092 = state_in[47:40] ;
assign n5093 =  ( n5092 ) == ( bv_8_146_n337 )  ;
assign n5094 = state_in[47:40] ;
assign n5095 =  ( n5094 ) == ( bv_8_145_n397 )  ;
assign n5096 = state_in[47:40] ;
assign n5097 =  ( n5096 ) == ( bv_8_144_n173 )  ;
assign n5098 = state_in[47:40] ;
assign n5099 =  ( n5098 ) == ( bv_8_143_n403 )  ;
assign n5100 = state_in[47:40] ;
assign n5101 =  ( n5100 ) == ( bv_8_142_n406 )  ;
assign n5102 = state_in[47:40] ;
assign n5103 =  ( n5102 ) == ( bv_8_141_n410 )  ;
assign n5104 = state_in[47:40] ;
assign n5105 =  ( n5104 ) == ( bv_8_140_n376 )  ;
assign n5106 = state_in[47:40] ;
assign n5107 =  ( n5106 ) == ( bv_8_139_n297 )  ;
assign n5108 = state_in[47:40] ;
assign n5109 =  ( n5108 ) == ( bv_8_138_n418 )  ;
assign n5110 = state_in[47:40] ;
assign n5111 =  ( n5110 ) == ( bv_8_137_n421 )  ;
assign n5112 = state_in[47:40] ;
assign n5113 =  ( n5112 ) == ( bv_8_136_n425 )  ;
assign n5114 = state_in[47:40] ;
assign n5115 =  ( n5114 ) == ( bv_8_135_n81 )  ;
assign n5116 = state_in[47:40] ;
assign n5117 =  ( n5116 ) == ( bv_8_134_n431 )  ;
assign n5118 = state_in[47:40] ;
assign n5119 =  ( n5118 ) == ( bv_8_133_n434 )  ;
assign n5120 = state_in[47:40] ;
assign n5121 =  ( n5120 ) == ( bv_8_132_n41 )  ;
assign n5122 = state_in[47:40] ;
assign n5123 =  ( n5122 ) == ( bv_8_131_n440 )  ;
assign n5124 = state_in[47:40] ;
assign n5125 =  ( n5124 ) == ( bv_8_130_n33 )  ;
assign n5126 = state_in[47:40] ;
assign n5127 =  ( n5126 ) == ( bv_8_129_n446 )  ;
assign n5128 = state_in[47:40] ;
assign n5129 =  ( n5128 ) == ( bv_8_128_n450 )  ;
assign n5130 = state_in[47:40] ;
assign n5131 =  ( n5130 ) == ( bv_8_127_n453 )  ;
assign n5132 = state_in[47:40] ;
assign n5133 =  ( n5132 ) == ( bv_8_126_n456 )  ;
assign n5134 = state_in[47:40] ;
assign n5135 =  ( n5134 ) == ( bv_8_125_n459 )  ;
assign n5136 = state_in[47:40] ;
assign n5137 =  ( n5136 ) == ( bv_8_124_n184 )  ;
assign n5138 = state_in[47:40] ;
assign n5139 =  ( n5138 ) == ( bv_8_123_n17 )  ;
assign n5140 = state_in[47:40] ;
assign n5141 =  ( n5140 ) == ( bv_8_122_n416 )  ;
assign n5142 = state_in[47:40] ;
assign n5143 =  ( n5142 ) == ( bv_8_121_n470 )  ;
assign n5144 = state_in[47:40] ;
assign n5145 =  ( n5144 ) == ( bv_8_120_n474 )  ;
assign n5146 = state_in[47:40] ;
assign n5147 =  ( n5146 ) == ( bv_8_119_n472 )  ;
assign n5148 = state_in[47:40] ;
assign n5149 =  ( n5148 ) == ( bv_8_118_n480 )  ;
assign n5150 = state_in[47:40] ;
assign n5151 =  ( n5150 ) == ( bv_8_117_n484 )  ;
assign n5152 = state_in[47:40] ;
assign n5153 =  ( n5152 ) == ( bv_8_116_n345 )  ;
assign n5154 = state_in[47:40] ;
assign n5155 =  ( n5154 ) == ( bv_8_115_n222 )  ;
assign n5156 = state_in[47:40] ;
assign n5157 =  ( n5156 ) == ( bv_8_114_n494 )  ;
assign n5158 = state_in[47:40] ;
assign n5159 =  ( n5158 ) == ( bv_8_113_n180 )  ;
assign n5160 = state_in[47:40] ;
assign n5161 =  ( n5160 ) == ( bv_8_112_n482 )  ;
assign n5162 = state_in[47:40] ;
assign n5163 =  ( n5162 ) == ( bv_8_111_n244 )  ;
assign n5164 = state_in[47:40] ;
assign n5165 =  ( n5164 ) == ( bv_8_110_n294 )  ;
assign n5166 = state_in[47:40] ;
assign n5167 =  ( n5166 ) == ( bv_8_109_n9 )  ;
assign n5168 = state_in[47:40] ;
assign n5169 =  ( n5168 ) == ( bv_8_108_n510 )  ;
assign n5170 = state_in[47:40] ;
assign n5171 =  ( n5170 ) == ( bv_8_107_n370 )  ;
assign n5172 = state_in[47:40] ;
assign n5173 =  ( n5172 ) == ( bv_8_106_n155 )  ;
assign n5174 = state_in[47:40] ;
assign n5175 =  ( n5174 ) == ( bv_8_105_n148 )  ;
assign n5176 = state_in[47:40] ;
assign n5177 =  ( n5176 ) == ( bv_8_104_n520 )  ;
assign n5178 = state_in[47:40] ;
assign n5179 =  ( n5178 ) == ( bv_8_103_n523 )  ;
assign n5180 = state_in[47:40] ;
assign n5181 =  ( n5180 ) == ( bv_8_102_n527 )  ;
assign n5182 = state_in[47:40] ;
assign n5183 =  ( n5182 ) == ( bv_8_101_n49 )  ;
assign n5184 = state_in[47:40] ;
assign n5185 =  ( n5184 ) == ( bv_8_100_n348 )  ;
assign n5186 = state_in[47:40] ;
assign n5187 =  ( n5186 ) == ( bv_8_99_n476 )  ;
assign n5188 = state_in[47:40] ;
assign n5189 =  ( n5188 ) == ( bv_8_98_n536 )  ;
assign n5190 = state_in[47:40] ;
assign n5191 =  ( n5190 ) == ( bv_8_97_n198 )  ;
assign n5192 = state_in[47:40] ;
assign n5193 =  ( n5192 ) == ( bv_8_96_n542 )  ;
assign n5194 = state_in[47:40] ;
assign n5195 =  ( n5194 ) == ( bv_8_95_n545 )  ;
assign n5196 = state_in[47:40] ;
assign n5197 =  ( n5196 ) == ( bv_8_94_n548 )  ;
assign n5198 = state_in[47:40] ;
assign n5199 =  ( n5198 ) == ( bv_8_93_n498 )  ;
assign n5200 = state_in[47:40] ;
assign n5201 =  ( n5200 ) == ( bv_8_92_n234 )  ;
assign n5202 = state_in[47:40] ;
assign n5203 =  ( n5202 ) == ( bv_8_91_n555 )  ;
assign n5204 = state_in[47:40] ;
assign n5205 =  ( n5204 ) == ( bv_8_90_n25 )  ;
assign n5206 = state_in[47:40] ;
assign n5207 =  ( n5206 ) == ( bv_8_89_n61 )  ;
assign n5208 = state_in[47:40] ;
assign n5209 =  ( n5208 ) == ( bv_8_88_n562 )  ;
assign n5210 = state_in[47:40] ;
assign n5211 =  ( n5210 ) == ( bv_8_87_n226 )  ;
assign n5212 = state_in[47:40] ;
assign n5213 =  ( n5212 ) == ( bv_8_86_n567 )  ;
assign n5214 = state_in[47:40] ;
assign n5215 =  ( n5214 ) == ( bv_8_85_n423 )  ;
assign n5216 = state_in[47:40] ;
assign n5217 =  ( n5216 ) == ( bv_8_84_n386 )  ;
assign n5218 = state_in[47:40] ;
assign n5219 =  ( n5218 ) == ( bv_8_83_n575 )  ;
assign n5220 = state_in[47:40] ;
assign n5221 =  ( n5220 ) == ( bv_8_82_n578 )  ;
assign n5222 = state_in[47:40] ;
assign n5223 =  ( n5222 ) == ( bv_8_81_n582 )  ;
assign n5224 = state_in[47:40] ;
assign n5225 =  ( n5224 ) == ( bv_8_80_n73 )  ;
assign n5226 = state_in[47:40] ;
assign n5227 =  ( n5226 ) == ( bv_8_79_n538 )  ;
assign n5228 = state_in[47:40] ;
assign n5229 =  ( n5228 ) == ( bv_8_78_n590 )  ;
assign n5230 = state_in[47:40] ;
assign n5231 =  ( n5230 ) == ( bv_8_77_n593 )  ;
assign n5232 = state_in[47:40] ;
assign n5233 =  ( n5232 ) == ( bv_8_76_n596 )  ;
assign n5234 = state_in[47:40] ;
assign n5235 =  ( n5234 ) == ( bv_8_75_n503 )  ;
assign n5236 = state_in[47:40] ;
assign n5237 =  ( n5236 ) == ( bv_8_74_n237 )  ;
assign n5238 = state_in[47:40] ;
assign n5239 =  ( n5238 ) == ( bv_8_73_n275 )  ;
assign n5240 = state_in[47:40] ;
assign n5241 =  ( n5240 ) == ( bv_8_72_n330 )  ;
assign n5242 = state_in[47:40] ;
assign n5243 =  ( n5242 ) == ( bv_8_71_n252 )  ;
assign n5244 = state_in[47:40] ;
assign n5245 =  ( n5244 ) == ( bv_8_70_n609 )  ;
assign n5246 = state_in[47:40] ;
assign n5247 =  ( n5246 ) == ( bv_8_69_n612 )  ;
assign n5248 = state_in[47:40] ;
assign n5249 =  ( n5248 ) == ( bv_8_68_n390 )  ;
assign n5250 = state_in[47:40] ;
assign n5251 =  ( n5250 ) == ( bv_8_67_n318 )  ;
assign n5252 = state_in[47:40] ;
assign n5253 =  ( n5252 ) == ( bv_8_66_n466 )  ;
assign n5254 = state_in[47:40] ;
assign n5255 =  ( n5254 ) == ( bv_8_65_n623 )  ;
assign n5256 = state_in[47:40] ;
assign n5257 =  ( n5256 ) == ( bv_8_64_n573 )  ;
assign n5258 = state_in[47:40] ;
assign n5259 =  ( n5258 ) == ( bv_8_63_n489 )  ;
assign n5260 = state_in[47:40] ;
assign n5261 =  ( n5260 ) == ( bv_8_62_n205 )  ;
assign n5262 = state_in[47:40] ;
assign n5263 =  ( n5262 ) == ( bv_8_61_n634 )  ;
assign n5264 = state_in[47:40] ;
assign n5265 =  ( n5264 ) == ( bv_8_60_n93 )  ;
assign n5266 = state_in[47:40] ;
assign n5267 =  ( n5266 ) == ( bv_8_59_n382 )  ;
assign n5268 = state_in[47:40] ;
assign n5269 =  ( n5268 ) == ( bv_8_58_n136 )  ;
assign n5270 = state_in[47:40] ;
assign n5271 =  ( n5270 ) == ( bv_8_57_n312 )  ;
assign n5272 = state_in[47:40] ;
assign n5273 =  ( n5272 ) == ( bv_8_56_n230 )  ;
assign n5274 = state_in[47:40] ;
assign n5275 =  ( n5274 ) == ( bv_8_55_n650 )  ;
assign n5276 = state_in[47:40] ;
assign n5277 =  ( n5276 ) == ( bv_8_54_n616 )  ;
assign n5278 = state_in[47:40] ;
assign n5279 =  ( n5278 ) == ( bv_8_53_n436 )  ;
assign n5280 = state_in[47:40] ;
assign n5281 =  ( n5280 ) == ( bv_8_52_n619 )  ;
assign n5282 = state_in[47:40] ;
assign n5283 =  ( n5282 ) == ( bv_8_51_n101 )  ;
assign n5284 = state_in[47:40] ;
assign n5285 =  ( n5284 ) == ( bv_8_50_n408 )  ;
assign n5286 = state_in[47:40] ;
assign n5287 =  ( n5286 ) == ( bv_8_49_n309 )  ;
assign n5288 = state_in[47:40] ;
assign n5289 =  ( n5288 ) == ( bv_8_48_n660 )  ;
assign n5290 = state_in[47:40] ;
assign n5291 =  ( n5290 ) == ( bv_8_47_n652 )  ;
assign n5292 = state_in[47:40] ;
assign n5293 =  ( n5292 ) == ( bv_8_46_n429 )  ;
assign n5294 = state_in[47:40] ;
assign n5295 =  ( n5294 ) == ( bv_8_45_n97 )  ;
assign n5296 = state_in[47:40] ;
assign n5297 =  ( n5296 ) == ( bv_8_44_n5 )  ;
assign n5298 = state_in[47:40] ;
assign n5299 =  ( n5298 ) == ( bv_8_43_n121 )  ;
assign n5300 = state_in[47:40] ;
assign n5301 =  ( n5300 ) == ( bv_8_42_n672 )  ;
assign n5302 = state_in[47:40] ;
assign n5303 =  ( n5302 ) == ( bv_8_41_n29 )  ;
assign n5304 = state_in[47:40] ;
assign n5305 =  ( n5304 ) == ( bv_8_40_n366 )  ;
assign n5306 = state_in[47:40] ;
assign n5307 =  ( n5306 ) == ( bv_8_39_n132 )  ;
assign n5308 = state_in[47:40] ;
assign n5309 =  ( n5308 ) == ( bv_8_38_n444 )  ;
assign n5310 = state_in[47:40] ;
assign n5311 =  ( n5310 ) == ( bv_8_37_n506 )  ;
assign n5312 = state_in[47:40] ;
assign n5313 =  ( n5312 ) == ( bv_8_36_n645 )  ;
assign n5314 = state_in[47:40] ;
assign n5315 =  ( n5314 ) == ( bv_8_35_n696 )  ;
assign n5316 = state_in[47:40] ;
assign n5317 =  ( n5316 ) == ( bv_8_34_n117 )  ;
assign n5318 = state_in[47:40] ;
assign n5319 =  ( n5318 ) == ( bv_8_33_n486 )  ;
assign n5320 = state_in[47:40] ;
assign n5321 =  ( n5320 ) == ( bv_8_32_n463 )  ;
assign n5322 = state_in[47:40] ;
assign n5323 =  ( n5322 ) == ( bv_8_31_n705 )  ;
assign n5324 = state_in[47:40] ;
assign n5325 =  ( n5324 ) == ( bv_8_30_n21 )  ;
assign n5326 = state_in[47:40] ;
assign n5327 =  ( n5326 ) == ( bv_8_29_n625 )  ;
assign n5328 = state_in[47:40] ;
assign n5329 =  ( n5328 ) == ( bv_8_28_n162 )  ;
assign n5330 = state_in[47:40] ;
assign n5331 =  ( n5330 ) == ( bv_8_27_n642 )  ;
assign n5332 = state_in[47:40] ;
assign n5333 =  ( n5332 ) == ( bv_8_26_n53 )  ;
assign n5334 = state_in[47:40] ;
assign n5335 =  ( n5334 ) == ( bv_8_25_n399 )  ;
assign n5336 = state_in[47:40] ;
assign n5337 =  ( n5336 ) == ( bv_8_24_n448 )  ;
assign n5338 = state_in[47:40] ;
assign n5339 =  ( n5338 ) == ( bv_8_23_n144 )  ;
assign n5340 = state_in[47:40] ;
assign n5341 =  ( n5340 ) == ( bv_8_22_n357 )  ;
assign n5342 = state_in[47:40] ;
assign n5343 =  ( n5342 ) == ( bv_8_21_n89 )  ;
assign n5344 = state_in[47:40] ;
assign n5345 =  ( n5344 ) == ( bv_8_20_n341 )  ;
assign n5346 = state_in[47:40] ;
assign n5347 =  ( n5346 ) == ( bv_8_19_n588 )  ;
assign n5348 = state_in[47:40] ;
assign n5349 =  ( n5348 ) == ( bv_8_18_n628 )  ;
assign n5350 = state_in[47:40] ;
assign n5351 =  ( n5350 ) == ( bv_8_17_n525 )  ;
assign n5352 = state_in[47:40] ;
assign n5353 =  ( n5352 ) == ( bv_8_16_n248 )  ;
assign n5354 = state_in[47:40] ;
assign n5355 =  ( n5354 ) == ( bv_8_15_n190 )  ;
assign n5356 = state_in[47:40] ;
assign n5357 =  ( n5356 ) == ( bv_8_14_n648 )  ;
assign n5358 = state_in[47:40] ;
assign n5359 =  ( n5358 ) == ( bv_8_13_n194 )  ;
assign n5360 = state_in[47:40] ;
assign n5361 =  ( n5360 ) == ( bv_8_12_n333 )  ;
assign n5362 = state_in[47:40] ;
assign n5363 =  ( n5362 ) == ( bv_8_11_n379 )  ;
assign n5364 = state_in[47:40] ;
assign n5365 =  ( n5364 ) == ( bv_8_10_n655 )  ;
assign n5366 = state_in[47:40] ;
assign n5367 =  ( n5366 ) == ( bv_8_9_n57 )  ;
assign n5368 = state_in[47:40] ;
assign n5369 =  ( n5368 ) == ( bv_8_8_n669 )  ;
assign n5370 = state_in[47:40] ;
assign n5371 =  ( n5370 ) == ( bv_8_7_n105 )  ;
assign n5372 = state_in[47:40] ;
assign n5373 =  ( n5372 ) == ( bv_8_6_n169 )  ;
assign n5374 = state_in[47:40] ;
assign n5375 =  ( n5374 ) == ( bv_8_5_n492 )  ;
assign n5376 = state_in[47:40] ;
assign n5377 =  ( n5376 ) == ( bv_8_4_n516 )  ;
assign n5378 = state_in[47:40] ;
assign n5379 =  ( n5378 ) == ( bv_8_3_n65 )  ;
assign n5380 = state_in[47:40] ;
assign n5381 =  ( n5380 ) == ( bv_8_2_n751 )  ;
assign n5382 = state_in[47:40] ;
assign n5383 =  ( n5382 ) == ( bv_8_1_n287 )  ;
assign n5384 = state_in[47:40] ;
assign n5385 =  ( n5384 ) == ( bv_8_0_n580 )  ;
assign n5386 =  ( n5385 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n5387 =  ( n5383 ) ? ( bv_8_248_n31 ) : ( n5386 ) ;
assign n5388 =  ( n5381 ) ? ( bv_8_238_n71 ) : ( n5387 ) ;
assign n5389 =  ( n5379 ) ? ( bv_8_246_n39 ) : ( n5388 ) ;
assign n5390 =  ( n5377 ) ? ( bv_8_255_n3 ) : ( n5389 ) ;
assign n5391 =  ( n5375 ) ? ( bv_8_214_n164 ) : ( n5390 ) ;
assign n5392 =  ( n5373 ) ? ( bv_8_222_n134 ) : ( n5391 ) ;
assign n5393 =  ( n5371 ) ? ( bv_8_145_n397 ) : ( n5392 ) ;
assign n5394 =  ( n5369 ) ? ( bv_8_96_n542 ) : ( n5393 ) ;
assign n5395 =  ( n5367 ) ? ( bv_8_2_n751 ) : ( n5394 ) ;
assign n5396 =  ( n5365 ) ? ( bv_8_206_n192 ) : ( n5395 ) ;
assign n5397 =  ( n5363 ) ? ( bv_8_86_n567 ) : ( n5396 ) ;
assign n5398 =  ( n5361 ) ? ( bv_8_231_n99 ) : ( n5397 ) ;
assign n5399 =  ( n5359 ) ? ( bv_8_181_n281 ) : ( n5398 ) ;
assign n5400 =  ( n5357 ) ? ( bv_8_77_n593 ) : ( n5399 ) ;
assign n5401 =  ( n5355 ) ? ( bv_8_236_n79 ) : ( n5400 ) ;
assign n5402 =  ( n5353 ) ? ( bv_8_143_n403 ) : ( n5401 ) ;
assign n5403 =  ( n5351 ) ? ( bv_8_31_n705 ) : ( n5402 ) ;
assign n5404 =  ( n5349 ) ? ( bv_8_137_n421 ) : ( n5403 ) ;
assign n5405 =  ( n5347 ) ? ( bv_8_250_n23 ) : ( n5404 ) ;
assign n5406 =  ( n5345 ) ? ( bv_8_239_n67 ) : ( n5405 ) ;
assign n5407 =  ( n5343 ) ? ( bv_8_178_n292 ) : ( n5406 ) ;
assign n5408 =  ( n5341 ) ? ( bv_8_142_n406 ) : ( n5407 ) ;
assign n5409 =  ( n5339 ) ? ( bv_8_251_n19 ) : ( n5408 ) ;
assign n5410 =  ( n5337 ) ? ( bv_8_65_n623 ) : ( n5409 ) ;
assign n5411 =  ( n5335 ) ? ( bv_8_179_n289 ) : ( n5410 ) ;
assign n5412 =  ( n5333 ) ? ( bv_8_95_n545 ) : ( n5411 ) ;
assign n5413 =  ( n5331 ) ? ( bv_8_69_n612 ) : ( n5412 ) ;
assign n5414 =  ( n5329 ) ? ( bv_8_35_n696 ) : ( n5413 ) ;
assign n5415 =  ( n5327 ) ? ( bv_8_83_n575 ) : ( n5414 ) ;
assign n5416 =  ( n5325 ) ? ( bv_8_228_n111 ) : ( n5415 ) ;
assign n5417 =  ( n5323 ) ? ( bv_8_155_n364 ) : ( n5416 ) ;
assign n5418 =  ( n5321 ) ? ( bv_8_117_n484 ) : ( n5417 ) ;
assign n5419 =  ( n5319 ) ? ( bv_8_225_n123 ) : ( n5418 ) ;
assign n5420 =  ( n5317 ) ? ( bv_8_61_n634 ) : ( n5419 ) ;
assign n5421 =  ( n5315 ) ? ( bv_8_76_n596 ) : ( n5420 ) ;
assign n5422 =  ( n5313 ) ? ( bv_8_108_n510 ) : ( n5421 ) ;
assign n5423 =  ( n5311 ) ? ( bv_8_126_n456 ) : ( n5422 ) ;
assign n5424 =  ( n5309 ) ? ( bv_8_245_n43 ) : ( n5423 ) ;
assign n5425 =  ( n5307 ) ? ( bv_8_131_n440 ) : ( n5424 ) ;
assign n5426 =  ( n5305 ) ? ( bv_8_104_n520 ) : ( n5425 ) ;
assign n5427 =  ( n5303 ) ? ( bv_8_81_n582 ) : ( n5426 ) ;
assign n5428 =  ( n5301 ) ? ( bv_8_209_n182 ) : ( n5427 ) ;
assign n5429 =  ( n5299 ) ? ( bv_8_249_n27 ) : ( n5428 ) ;
assign n5430 =  ( n5297 ) ? ( bv_8_226_n119 ) : ( n5429 ) ;
assign n5431 =  ( n5295 ) ? ( bv_8_171_n314 ) : ( n5430 ) ;
assign n5432 =  ( n5293 ) ? ( bv_8_98_n536 ) : ( n5431 ) ;
assign n5433 =  ( n5291 ) ? ( bv_8_42_n672 ) : ( n5432 ) ;
assign n5434 =  ( n5289 ) ? ( bv_8_8_n669 ) : ( n5433 ) ;
assign n5435 =  ( n5287 ) ? ( bv_8_149_n384 ) : ( n5434 ) ;
assign n5436 =  ( n5285 ) ? ( bv_8_70_n609 ) : ( n5435 ) ;
assign n5437 =  ( n5283 ) ? ( bv_8_157_n359 ) : ( n5436 ) ;
assign n5438 =  ( n5281 ) ? ( bv_8_48_n660 ) : ( n5437 ) ;
assign n5439 =  ( n5279 ) ? ( bv_8_55_n650 ) : ( n5438 ) ;
assign n5440 =  ( n5277 ) ? ( bv_8_10_n655 ) : ( n5439 ) ;
assign n5441 =  ( n5275 ) ? ( bv_8_47_n652 ) : ( n5440 ) ;
assign n5442 =  ( n5273 ) ? ( bv_8_14_n648 ) : ( n5441 ) ;
assign n5443 =  ( n5271 ) ? ( bv_8_36_n645 ) : ( n5442 ) ;
assign n5444 =  ( n5269 ) ? ( bv_8_27_n642 ) : ( n5443 ) ;
assign n5445 =  ( n5267 ) ? ( bv_8_223_n130 ) : ( n5444 ) ;
assign n5446 =  ( n5265 ) ? ( bv_8_205_n196 ) : ( n5445 ) ;
assign n5447 =  ( n5263 ) ? ( bv_8_78_n590 ) : ( n5446 ) ;
assign n5448 =  ( n5261 ) ? ( bv_8_127_n453 ) : ( n5447 ) ;
assign n5449 =  ( n5259 ) ? ( bv_8_234_n87 ) : ( n5448 ) ;
assign n5450 =  ( n5257 ) ? ( bv_8_18_n628 ) : ( n5449 ) ;
assign n5451 =  ( n5255 ) ? ( bv_8_29_n625 ) : ( n5450 ) ;
assign n5452 =  ( n5253 ) ? ( bv_8_88_n562 ) : ( n5451 ) ;
assign n5453 =  ( n5251 ) ? ( bv_8_52_n619 ) : ( n5452 ) ;
assign n5454 =  ( n5249 ) ? ( bv_8_54_n616 ) : ( n5453 ) ;
assign n5455 =  ( n5247 ) ? ( bv_8_220_n142 ) : ( n5454 ) ;
assign n5456 =  ( n5245 ) ? ( bv_8_180_n285 ) : ( n5455 ) ;
assign n5457 =  ( n5243 ) ? ( bv_8_91_n555 ) : ( n5456 ) ;
assign n5458 =  ( n5241 ) ? ( bv_8_164_n335 ) : ( n5457 ) ;
assign n5459 =  ( n5239 ) ? ( bv_8_118_n480 ) : ( n5458 ) ;
assign n5460 =  ( n5237 ) ? ( bv_8_183_n273 ) : ( n5459 ) ;
assign n5461 =  ( n5235 ) ? ( bv_8_125_n459 ) : ( n5460 ) ;
assign n5462 =  ( n5233 ) ? ( bv_8_82_n578 ) : ( n5461 ) ;
assign n5463 =  ( n5231 ) ? ( bv_8_221_n138 ) : ( n5462 ) ;
assign n5464 =  ( n5229 ) ? ( bv_8_94_n548 ) : ( n5463 ) ;
assign n5465 =  ( n5227 ) ? ( bv_8_19_n588 ) : ( n5464 ) ;
assign n5466 =  ( n5225 ) ? ( bv_8_166_n328 ) : ( n5465 ) ;
assign n5467 =  ( n5223 ) ? ( bv_8_185_n266 ) : ( n5466 ) ;
assign n5468 =  ( n5221 ) ? ( bv_8_0_n580 ) : ( n5467 ) ;
assign n5469 =  ( n5219 ) ? ( bv_8_193_n239 ) : ( n5468 ) ;
assign n5470 =  ( n5217 ) ? ( bv_8_64_n573 ) : ( n5469 ) ;
assign n5471 =  ( n5215 ) ? ( bv_8_227_n115 ) : ( n5470 ) ;
assign n5472 =  ( n5213 ) ? ( bv_8_121_n470 ) : ( n5471 ) ;
assign n5473 =  ( n5211 ) ? ( bv_8_182_n277 ) : ( n5472 ) ;
assign n5474 =  ( n5209 ) ? ( bv_8_212_n171 ) : ( n5473 ) ;
assign n5475 =  ( n5207 ) ? ( bv_8_141_n410 ) : ( n5474 ) ;
assign n5476 =  ( n5205 ) ? ( bv_8_103_n523 ) : ( n5475 ) ;
assign n5477 =  ( n5203 ) ? ( bv_8_114_n494 ) : ( n5476 ) ;
assign n5478 =  ( n5201 ) ? ( bv_8_148_n388 ) : ( n5477 ) ;
assign n5479 =  ( n5199 ) ? ( bv_8_152_n374 ) : ( n5478 ) ;
assign n5480 =  ( n5197 ) ? ( bv_8_176_n299 ) : ( n5479 ) ;
assign n5481 =  ( n5195 ) ? ( bv_8_133_n434 ) : ( n5480 ) ;
assign n5482 =  ( n5193 ) ? ( bv_8_187_n260 ) : ( n5481 ) ;
assign n5483 =  ( n5191 ) ? ( bv_8_197_n224 ) : ( n5482 ) ;
assign n5484 =  ( n5189 ) ? ( bv_8_79_n538 ) : ( n5483 ) ;
assign n5485 =  ( n5187 ) ? ( bv_8_237_n75 ) : ( n5484 ) ;
assign n5486 =  ( n5185 ) ? ( bv_8_134_n431 ) : ( n5485 ) ;
assign n5487 =  ( n5183 ) ? ( bv_8_154_n368 ) : ( n5486 ) ;
assign n5488 =  ( n5181 ) ? ( bv_8_102_n527 ) : ( n5487 ) ;
assign n5489 =  ( n5179 ) ? ( bv_8_17_n525 ) : ( n5488 ) ;
assign n5490 =  ( n5177 ) ? ( bv_8_138_n418 ) : ( n5489 ) ;
assign n5491 =  ( n5175 ) ? ( bv_8_233_n91 ) : ( n5490 ) ;
assign n5492 =  ( n5173 ) ? ( bv_8_4_n516 ) : ( n5491 ) ;
assign n5493 =  ( n5171 ) ? ( bv_8_254_n7 ) : ( n5492 ) ;
assign n5494 =  ( n5169 ) ? ( bv_8_160_n350 ) : ( n5493 ) ;
assign n5495 =  ( n5167 ) ? ( bv_8_120_n474 ) : ( n5494 ) ;
assign n5496 =  ( n5165 ) ? ( bv_8_37_n506 ) : ( n5495 ) ;
assign n5497 =  ( n5163 ) ? ( bv_8_75_n503 ) : ( n5496 ) ;
assign n5498 =  ( n5161 ) ? ( bv_8_162_n343 ) : ( n5497 ) ;
assign n5499 =  ( n5159 ) ? ( bv_8_93_n498 ) : ( n5498 ) ;
assign n5500 =  ( n5157 ) ? ( bv_8_128_n450 ) : ( n5499 ) ;
assign n5501 =  ( n5155 ) ? ( bv_8_5_n492 ) : ( n5500 ) ;
assign n5502 =  ( n5153 ) ? ( bv_8_63_n489 ) : ( n5501 ) ;
assign n5503 =  ( n5151 ) ? ( bv_8_33_n486 ) : ( n5502 ) ;
assign n5504 =  ( n5149 ) ? ( bv_8_112_n482 ) : ( n5503 ) ;
assign n5505 =  ( n5147 ) ? ( bv_8_241_n59 ) : ( n5504 ) ;
assign n5506 =  ( n5145 ) ? ( bv_8_99_n476 ) : ( n5505 ) ;
assign n5507 =  ( n5143 ) ? ( bv_8_119_n472 ) : ( n5506 ) ;
assign n5508 =  ( n5141 ) ? ( bv_8_175_n302 ) : ( n5507 ) ;
assign n5509 =  ( n5139 ) ? ( bv_8_66_n466 ) : ( n5508 ) ;
assign n5510 =  ( n5137 ) ? ( bv_8_32_n463 ) : ( n5509 ) ;
assign n5511 =  ( n5135 ) ? ( bv_8_229_n107 ) : ( n5510 ) ;
assign n5512 =  ( n5133 ) ? ( bv_8_253_n11 ) : ( n5511 ) ;
assign n5513 =  ( n5131 ) ? ( bv_8_191_n246 ) : ( n5512 ) ;
assign n5514 =  ( n5129 ) ? ( bv_8_129_n446 ) : ( n5513 ) ;
assign n5515 =  ( n5127 ) ? ( bv_8_24_n448 ) : ( n5514 ) ;
assign n5516 =  ( n5125 ) ? ( bv_8_38_n444 ) : ( n5515 ) ;
assign n5517 =  ( n5123 ) ? ( bv_8_195_n232 ) : ( n5516 ) ;
assign n5518 =  ( n5121 ) ? ( bv_8_190_n250 ) : ( n5517 ) ;
assign n5519 =  ( n5119 ) ? ( bv_8_53_n436 ) : ( n5518 ) ;
assign n5520 =  ( n5117 ) ? ( bv_8_136_n425 ) : ( n5519 ) ;
assign n5521 =  ( n5115 ) ? ( bv_8_46_n429 ) : ( n5520 ) ;
assign n5522 =  ( n5113 ) ? ( bv_8_147_n392 ) : ( n5521 ) ;
assign n5523 =  ( n5111 ) ? ( bv_8_85_n423 ) : ( n5522 ) ;
assign n5524 =  ( n5109 ) ? ( bv_8_252_n15 ) : ( n5523 ) ;
assign n5525 =  ( n5107 ) ? ( bv_8_122_n416 ) : ( n5524 ) ;
assign n5526 =  ( n5105 ) ? ( bv_8_200_n213 ) : ( n5525 ) ;
assign n5527 =  ( n5103 ) ? ( bv_8_186_n263 ) : ( n5526 ) ;
assign n5528 =  ( n5101 ) ? ( bv_8_50_n408 ) : ( n5527 ) ;
assign n5529 =  ( n5099 ) ? ( bv_8_230_n103 ) : ( n5528 ) ;
assign n5530 =  ( n5097 ) ? ( bv_8_192_n242 ) : ( n5529 ) ;
assign n5531 =  ( n5095 ) ? ( bv_8_25_n399 ) : ( n5530 ) ;
assign n5532 =  ( n5093 ) ? ( bv_8_158_n355 ) : ( n5531 ) ;
assign n5533 =  ( n5091 ) ? ( bv_8_163_n339 ) : ( n5532 ) ;
assign n5534 =  ( n5089 ) ? ( bv_8_68_n390 ) : ( n5533 ) ;
assign n5535 =  ( n5087 ) ? ( bv_8_84_n386 ) : ( n5534 ) ;
assign n5536 =  ( n5085 ) ? ( bv_8_59_n382 ) : ( n5535 ) ;
assign n5537 =  ( n5083 ) ? ( bv_8_11_n379 ) : ( n5536 ) ;
assign n5538 =  ( n5081 ) ? ( bv_8_140_n376 ) : ( n5537 ) ;
assign n5539 =  ( n5079 ) ? ( bv_8_199_n216 ) : ( n5538 ) ;
assign n5540 =  ( n5077 ) ? ( bv_8_107_n370 ) : ( n5539 ) ;
assign n5541 =  ( n5075 ) ? ( bv_8_40_n366 ) : ( n5540 ) ;
assign n5542 =  ( n5073 ) ? ( bv_8_167_n325 ) : ( n5541 ) ;
assign n5543 =  ( n5071 ) ? ( bv_8_188_n257 ) : ( n5542 ) ;
assign n5544 =  ( n5069 ) ? ( bv_8_22_n357 ) : ( n5543 ) ;
assign n5545 =  ( n5067 ) ? ( bv_8_173_n307 ) : ( n5544 ) ;
assign n5546 =  ( n5065 ) ? ( bv_8_219_n146 ) : ( n5545 ) ;
assign n5547 =  ( n5063 ) ? ( bv_8_100_n348 ) : ( n5546 ) ;
assign n5548 =  ( n5061 ) ? ( bv_8_116_n345 ) : ( n5547 ) ;
assign n5549 =  ( n5059 ) ? ( bv_8_20_n341 ) : ( n5548 ) ;
assign n5550 =  ( n5057 ) ? ( bv_8_146_n337 ) : ( n5549 ) ;
assign n5551 =  ( n5055 ) ? ( bv_8_12_n333 ) : ( n5550 ) ;
assign n5552 =  ( n5053 ) ? ( bv_8_72_n330 ) : ( n5551 ) ;
assign n5553 =  ( n5051 ) ? ( bv_8_184_n270 ) : ( n5552 ) ;
assign n5554 =  ( n5049 ) ? ( bv_8_159_n323 ) : ( n5553 ) ;
assign n5555 =  ( n5047 ) ? ( bv_8_189_n254 ) : ( n5554 ) ;
assign n5556 =  ( n5045 ) ? ( bv_8_67_n318 ) : ( n5555 ) ;
assign n5557 =  ( n5043 ) ? ( bv_8_196_n228 ) : ( n5556 ) ;
assign n5558 =  ( n5041 ) ? ( bv_8_57_n312 ) : ( n5557 ) ;
assign n5559 =  ( n5039 ) ? ( bv_8_49_n309 ) : ( n5558 ) ;
assign n5560 =  ( n5037 ) ? ( bv_8_211_n175 ) : ( n5559 ) ;
assign n5561 =  ( n5035 ) ? ( bv_8_242_n55 ) : ( n5560 ) ;
assign n5562 =  ( n5033 ) ? ( bv_8_213_n167 ) : ( n5561 ) ;
assign n5563 =  ( n5031 ) ? ( bv_8_139_n297 ) : ( n5562 ) ;
assign n5564 =  ( n5029 ) ? ( bv_8_110_n294 ) : ( n5563 ) ;
assign n5565 =  ( n5027 ) ? ( bv_8_218_n150 ) : ( n5564 ) ;
assign n5566 =  ( n5025 ) ? ( bv_8_1_n287 ) : ( n5565 ) ;
assign n5567 =  ( n5023 ) ? ( bv_8_177_n283 ) : ( n5566 ) ;
assign n5568 =  ( n5021 ) ? ( bv_8_156_n279 ) : ( n5567 ) ;
assign n5569 =  ( n5019 ) ? ( bv_8_73_n275 ) : ( n5568 ) ;
assign n5570 =  ( n5017 ) ? ( bv_8_216_n157 ) : ( n5569 ) ;
assign n5571 =  ( n5015 ) ? ( bv_8_172_n268 ) : ( n5570 ) ;
assign n5572 =  ( n5013 ) ? ( bv_8_243_n51 ) : ( n5571 ) ;
assign n5573 =  ( n5011 ) ? ( bv_8_207_n188 ) : ( n5572 ) ;
assign n5574 =  ( n5009 ) ? ( bv_8_202_n207 ) : ( n5573 ) ;
assign n5575 =  ( n5007 ) ? ( bv_8_244_n47 ) : ( n5574 ) ;
assign n5576 =  ( n5005 ) ? ( bv_8_71_n252 ) : ( n5575 ) ;
assign n5577 =  ( n5003 ) ? ( bv_8_16_n248 ) : ( n5576 ) ;
assign n5578 =  ( n5001 ) ? ( bv_8_111_n244 ) : ( n5577 ) ;
assign n5579 =  ( n4999 ) ? ( bv_8_240_n63 ) : ( n5578 ) ;
assign n5580 =  ( n4997 ) ? ( bv_8_74_n237 ) : ( n5579 ) ;
assign n5581 =  ( n4995 ) ? ( bv_8_92_n234 ) : ( n5580 ) ;
assign n5582 =  ( n4993 ) ? ( bv_8_56_n230 ) : ( n5581 ) ;
assign n5583 =  ( n4991 ) ? ( bv_8_87_n226 ) : ( n5582 ) ;
assign n5584 =  ( n4989 ) ? ( bv_8_115_n222 ) : ( n5583 ) ;
assign n5585 =  ( n4987 ) ? ( bv_8_151_n218 ) : ( n5584 ) ;
assign n5586 =  ( n4985 ) ? ( bv_8_203_n203 ) : ( n5585 ) ;
assign n5587 =  ( n4983 ) ? ( bv_8_161_n211 ) : ( n5586 ) ;
assign n5588 =  ( n4981 ) ? ( bv_8_232_n95 ) : ( n5587 ) ;
assign n5589 =  ( n4979 ) ? ( bv_8_62_n205 ) : ( n5588 ) ;
assign n5590 =  ( n4977 ) ? ( bv_8_150_n201 ) : ( n5589 ) ;
assign n5591 =  ( n4975 ) ? ( bv_8_97_n198 ) : ( n5590 ) ;
assign n5592 =  ( n4973 ) ? ( bv_8_13_n194 ) : ( n5591 ) ;
assign n5593 =  ( n4971 ) ? ( bv_8_15_n190 ) : ( n5592 ) ;
assign n5594 =  ( n4969 ) ? ( bv_8_224_n126 ) : ( n5593 ) ;
assign n5595 =  ( n4967 ) ? ( bv_8_124_n184 ) : ( n5594 ) ;
assign n5596 =  ( n4965 ) ? ( bv_8_113_n180 ) : ( n5595 ) ;
assign n5597 =  ( n4963 ) ? ( bv_8_204_n177 ) : ( n5596 ) ;
assign n5598 =  ( n4961 ) ? ( bv_8_144_n173 ) : ( n5597 ) ;
assign n5599 =  ( n4959 ) ? ( bv_8_6_n169 ) : ( n5598 ) ;
assign n5600 =  ( n4957 ) ? ( bv_8_247_n35 ) : ( n5599 ) ;
assign n5601 =  ( n4955 ) ? ( bv_8_28_n162 ) : ( n5600 ) ;
assign n5602 =  ( n4953 ) ? ( bv_8_194_n159 ) : ( n5601 ) ;
assign n5603 =  ( n4951 ) ? ( bv_8_106_n155 ) : ( n5602 ) ;
assign n5604 =  ( n4949 ) ? ( bv_8_174_n152 ) : ( n5603 ) ;
assign n5605 =  ( n4947 ) ? ( bv_8_105_n148 ) : ( n5604 ) ;
assign n5606 =  ( n4945 ) ? ( bv_8_23_n144 ) : ( n5605 ) ;
assign n5607 =  ( n4943 ) ? ( bv_8_153_n140 ) : ( n5606 ) ;
assign n5608 =  ( n4941 ) ? ( bv_8_58_n136 ) : ( n5607 ) ;
assign n5609 =  ( n4939 ) ? ( bv_8_39_n132 ) : ( n5608 ) ;
assign n5610 =  ( n4937 ) ? ( bv_8_217_n128 ) : ( n5609 ) ;
assign n5611 =  ( n4935 ) ? ( bv_8_235_n83 ) : ( n5610 ) ;
assign n5612 =  ( n4933 ) ? ( bv_8_43_n121 ) : ( n5611 ) ;
assign n5613 =  ( n4931 ) ? ( bv_8_34_n117 ) : ( n5612 ) ;
assign n5614 =  ( n4929 ) ? ( bv_8_210_n113 ) : ( n5613 ) ;
assign n5615 =  ( n4927 ) ? ( bv_8_169_n109 ) : ( n5614 ) ;
assign n5616 =  ( n4925 ) ? ( bv_8_7_n105 ) : ( n5615 ) ;
assign n5617 =  ( n4923 ) ? ( bv_8_51_n101 ) : ( n5616 ) ;
assign n5618 =  ( n4921 ) ? ( bv_8_45_n97 ) : ( n5617 ) ;
assign n5619 =  ( n4919 ) ? ( bv_8_60_n93 ) : ( n5618 ) ;
assign n5620 =  ( n4917 ) ? ( bv_8_21_n89 ) : ( n5619 ) ;
assign n5621 =  ( n4915 ) ? ( bv_8_201_n85 ) : ( n5620 ) ;
assign n5622 =  ( n4913 ) ? ( bv_8_135_n81 ) : ( n5621 ) ;
assign n5623 =  ( n4911 ) ? ( bv_8_170_n77 ) : ( n5622 ) ;
assign n5624 =  ( n4909 ) ? ( bv_8_80_n73 ) : ( n5623 ) ;
assign n5625 =  ( n4907 ) ? ( bv_8_165_n69 ) : ( n5624 ) ;
assign n5626 =  ( n4905 ) ? ( bv_8_3_n65 ) : ( n5625 ) ;
assign n5627 =  ( n4903 ) ? ( bv_8_89_n61 ) : ( n5626 ) ;
assign n5628 =  ( n4901 ) ? ( bv_8_9_n57 ) : ( n5627 ) ;
assign n5629 =  ( n4899 ) ? ( bv_8_26_n53 ) : ( n5628 ) ;
assign n5630 =  ( n4897 ) ? ( bv_8_101_n49 ) : ( n5629 ) ;
assign n5631 =  ( n4895 ) ? ( bv_8_215_n45 ) : ( n5630 ) ;
assign n5632 =  ( n4893 ) ? ( bv_8_132_n41 ) : ( n5631 ) ;
assign n5633 =  ( n4891 ) ? ( bv_8_208_n37 ) : ( n5632 ) ;
assign n5634 =  ( n4889 ) ? ( bv_8_130_n33 ) : ( n5633 ) ;
assign n5635 =  ( n4887 ) ? ( bv_8_41_n29 ) : ( n5634 ) ;
assign n5636 =  ( n4885 ) ? ( bv_8_90_n25 ) : ( n5635 ) ;
assign n5637 =  ( n4883 ) ? ( bv_8_30_n21 ) : ( n5636 ) ;
assign n5638 =  ( n4881 ) ? ( bv_8_123_n17 ) : ( n5637 ) ;
assign n5639 =  ( n4879 ) ? ( bv_8_168_n13 ) : ( n5638 ) ;
assign n5640 =  ( n4877 ) ? ( bv_8_109_n9 ) : ( n5639 ) ;
assign n5641 =  ( n4875 ) ? ( bv_8_44_n5 ) : ( n5640 ) ;
assign n5642 =  ( n4873 ) ^ ( n5641 )  ;
assign n5643 =  ( n5642 ) ^ ( n4100 )  ;
assign n5644 = key[119:112] ;
assign n5645 =  ( n5643 ) ^ ( n5644 )  ;
assign n5646 =  { ( n4103 ) , ( n5645 ) }  ;
assign n5647 =  ( n4871 ) ^ ( n1793 )  ;
assign n5648 =  ( n5647 ) ^ ( n5641 )  ;
assign n5649 =  ( n5648 ) ^ ( n4100 )  ;
assign n5650 = state_in[7:0] ;
assign n5651 =  ( n5650 ) == ( bv_8_255_n3 )  ;
assign n5652 = state_in[7:0] ;
assign n5653 =  ( n5652 ) == ( bv_8_254_n7 )  ;
assign n5654 = state_in[7:0] ;
assign n5655 =  ( n5654 ) == ( bv_8_253_n11 )  ;
assign n5656 = state_in[7:0] ;
assign n5657 =  ( n5656 ) == ( bv_8_252_n15 )  ;
assign n5658 = state_in[7:0] ;
assign n5659 =  ( n5658 ) == ( bv_8_251_n19 )  ;
assign n5660 = state_in[7:0] ;
assign n5661 =  ( n5660 ) == ( bv_8_250_n23 )  ;
assign n5662 = state_in[7:0] ;
assign n5663 =  ( n5662 ) == ( bv_8_249_n27 )  ;
assign n5664 = state_in[7:0] ;
assign n5665 =  ( n5664 ) == ( bv_8_248_n31 )  ;
assign n5666 = state_in[7:0] ;
assign n5667 =  ( n5666 ) == ( bv_8_247_n35 )  ;
assign n5668 = state_in[7:0] ;
assign n5669 =  ( n5668 ) == ( bv_8_246_n39 )  ;
assign n5670 = state_in[7:0] ;
assign n5671 =  ( n5670 ) == ( bv_8_245_n43 )  ;
assign n5672 = state_in[7:0] ;
assign n5673 =  ( n5672 ) == ( bv_8_244_n47 )  ;
assign n5674 = state_in[7:0] ;
assign n5675 =  ( n5674 ) == ( bv_8_243_n51 )  ;
assign n5676 = state_in[7:0] ;
assign n5677 =  ( n5676 ) == ( bv_8_242_n55 )  ;
assign n5678 = state_in[7:0] ;
assign n5679 =  ( n5678 ) == ( bv_8_241_n59 )  ;
assign n5680 = state_in[7:0] ;
assign n5681 =  ( n5680 ) == ( bv_8_240_n63 )  ;
assign n5682 = state_in[7:0] ;
assign n5683 =  ( n5682 ) == ( bv_8_239_n67 )  ;
assign n5684 = state_in[7:0] ;
assign n5685 =  ( n5684 ) == ( bv_8_238_n71 )  ;
assign n5686 = state_in[7:0] ;
assign n5687 =  ( n5686 ) == ( bv_8_237_n75 )  ;
assign n5688 = state_in[7:0] ;
assign n5689 =  ( n5688 ) == ( bv_8_236_n79 )  ;
assign n5690 = state_in[7:0] ;
assign n5691 =  ( n5690 ) == ( bv_8_235_n83 )  ;
assign n5692 = state_in[7:0] ;
assign n5693 =  ( n5692 ) == ( bv_8_234_n87 )  ;
assign n5694 = state_in[7:0] ;
assign n5695 =  ( n5694 ) == ( bv_8_233_n91 )  ;
assign n5696 = state_in[7:0] ;
assign n5697 =  ( n5696 ) == ( bv_8_232_n95 )  ;
assign n5698 = state_in[7:0] ;
assign n5699 =  ( n5698 ) == ( bv_8_231_n99 )  ;
assign n5700 = state_in[7:0] ;
assign n5701 =  ( n5700 ) == ( bv_8_230_n103 )  ;
assign n5702 = state_in[7:0] ;
assign n5703 =  ( n5702 ) == ( bv_8_229_n107 )  ;
assign n5704 = state_in[7:0] ;
assign n5705 =  ( n5704 ) == ( bv_8_228_n111 )  ;
assign n5706 = state_in[7:0] ;
assign n5707 =  ( n5706 ) == ( bv_8_227_n115 )  ;
assign n5708 = state_in[7:0] ;
assign n5709 =  ( n5708 ) == ( bv_8_226_n119 )  ;
assign n5710 = state_in[7:0] ;
assign n5711 =  ( n5710 ) == ( bv_8_225_n123 )  ;
assign n5712 = state_in[7:0] ;
assign n5713 =  ( n5712 ) == ( bv_8_224_n126 )  ;
assign n5714 = state_in[7:0] ;
assign n5715 =  ( n5714 ) == ( bv_8_223_n130 )  ;
assign n5716 = state_in[7:0] ;
assign n5717 =  ( n5716 ) == ( bv_8_222_n134 )  ;
assign n5718 = state_in[7:0] ;
assign n5719 =  ( n5718 ) == ( bv_8_221_n138 )  ;
assign n5720 = state_in[7:0] ;
assign n5721 =  ( n5720 ) == ( bv_8_220_n142 )  ;
assign n5722 = state_in[7:0] ;
assign n5723 =  ( n5722 ) == ( bv_8_219_n146 )  ;
assign n5724 = state_in[7:0] ;
assign n5725 =  ( n5724 ) == ( bv_8_218_n150 )  ;
assign n5726 = state_in[7:0] ;
assign n5727 =  ( n5726 ) == ( bv_8_217_n128 )  ;
assign n5728 = state_in[7:0] ;
assign n5729 =  ( n5728 ) == ( bv_8_216_n157 )  ;
assign n5730 = state_in[7:0] ;
assign n5731 =  ( n5730 ) == ( bv_8_215_n45 )  ;
assign n5732 = state_in[7:0] ;
assign n5733 =  ( n5732 ) == ( bv_8_214_n164 )  ;
assign n5734 = state_in[7:0] ;
assign n5735 =  ( n5734 ) == ( bv_8_213_n167 )  ;
assign n5736 = state_in[7:0] ;
assign n5737 =  ( n5736 ) == ( bv_8_212_n171 )  ;
assign n5738 = state_in[7:0] ;
assign n5739 =  ( n5738 ) == ( bv_8_211_n175 )  ;
assign n5740 = state_in[7:0] ;
assign n5741 =  ( n5740 ) == ( bv_8_210_n113 )  ;
assign n5742 = state_in[7:0] ;
assign n5743 =  ( n5742 ) == ( bv_8_209_n182 )  ;
assign n5744 = state_in[7:0] ;
assign n5745 =  ( n5744 ) == ( bv_8_208_n37 )  ;
assign n5746 = state_in[7:0] ;
assign n5747 =  ( n5746 ) == ( bv_8_207_n188 )  ;
assign n5748 = state_in[7:0] ;
assign n5749 =  ( n5748 ) == ( bv_8_206_n192 )  ;
assign n5750 = state_in[7:0] ;
assign n5751 =  ( n5750 ) == ( bv_8_205_n196 )  ;
assign n5752 = state_in[7:0] ;
assign n5753 =  ( n5752 ) == ( bv_8_204_n177 )  ;
assign n5754 = state_in[7:0] ;
assign n5755 =  ( n5754 ) == ( bv_8_203_n203 )  ;
assign n5756 = state_in[7:0] ;
assign n5757 =  ( n5756 ) == ( bv_8_202_n207 )  ;
assign n5758 = state_in[7:0] ;
assign n5759 =  ( n5758 ) == ( bv_8_201_n85 )  ;
assign n5760 = state_in[7:0] ;
assign n5761 =  ( n5760 ) == ( bv_8_200_n213 )  ;
assign n5762 = state_in[7:0] ;
assign n5763 =  ( n5762 ) == ( bv_8_199_n216 )  ;
assign n5764 = state_in[7:0] ;
assign n5765 =  ( n5764 ) == ( bv_8_198_n220 )  ;
assign n5766 = state_in[7:0] ;
assign n5767 =  ( n5766 ) == ( bv_8_197_n224 )  ;
assign n5768 = state_in[7:0] ;
assign n5769 =  ( n5768 ) == ( bv_8_196_n228 )  ;
assign n5770 = state_in[7:0] ;
assign n5771 =  ( n5770 ) == ( bv_8_195_n232 )  ;
assign n5772 = state_in[7:0] ;
assign n5773 =  ( n5772 ) == ( bv_8_194_n159 )  ;
assign n5774 = state_in[7:0] ;
assign n5775 =  ( n5774 ) == ( bv_8_193_n239 )  ;
assign n5776 = state_in[7:0] ;
assign n5777 =  ( n5776 ) == ( bv_8_192_n242 )  ;
assign n5778 = state_in[7:0] ;
assign n5779 =  ( n5778 ) == ( bv_8_191_n246 )  ;
assign n5780 = state_in[7:0] ;
assign n5781 =  ( n5780 ) == ( bv_8_190_n250 )  ;
assign n5782 = state_in[7:0] ;
assign n5783 =  ( n5782 ) == ( bv_8_189_n254 )  ;
assign n5784 = state_in[7:0] ;
assign n5785 =  ( n5784 ) == ( bv_8_188_n257 )  ;
assign n5786 = state_in[7:0] ;
assign n5787 =  ( n5786 ) == ( bv_8_187_n260 )  ;
assign n5788 = state_in[7:0] ;
assign n5789 =  ( n5788 ) == ( bv_8_186_n263 )  ;
assign n5790 = state_in[7:0] ;
assign n5791 =  ( n5790 ) == ( bv_8_185_n266 )  ;
assign n5792 = state_in[7:0] ;
assign n5793 =  ( n5792 ) == ( bv_8_184_n270 )  ;
assign n5794 = state_in[7:0] ;
assign n5795 =  ( n5794 ) == ( bv_8_183_n273 )  ;
assign n5796 = state_in[7:0] ;
assign n5797 =  ( n5796 ) == ( bv_8_182_n277 )  ;
assign n5798 = state_in[7:0] ;
assign n5799 =  ( n5798 ) == ( bv_8_181_n281 )  ;
assign n5800 = state_in[7:0] ;
assign n5801 =  ( n5800 ) == ( bv_8_180_n285 )  ;
assign n5802 = state_in[7:0] ;
assign n5803 =  ( n5802 ) == ( bv_8_179_n289 )  ;
assign n5804 = state_in[7:0] ;
assign n5805 =  ( n5804 ) == ( bv_8_178_n292 )  ;
assign n5806 = state_in[7:0] ;
assign n5807 =  ( n5806 ) == ( bv_8_177_n283 )  ;
assign n5808 = state_in[7:0] ;
assign n5809 =  ( n5808 ) == ( bv_8_176_n299 )  ;
assign n5810 = state_in[7:0] ;
assign n5811 =  ( n5810 ) == ( bv_8_175_n302 )  ;
assign n5812 = state_in[7:0] ;
assign n5813 =  ( n5812 ) == ( bv_8_174_n152 )  ;
assign n5814 = state_in[7:0] ;
assign n5815 =  ( n5814 ) == ( bv_8_173_n307 )  ;
assign n5816 = state_in[7:0] ;
assign n5817 =  ( n5816 ) == ( bv_8_172_n268 )  ;
assign n5818 = state_in[7:0] ;
assign n5819 =  ( n5818 ) == ( bv_8_171_n314 )  ;
assign n5820 = state_in[7:0] ;
assign n5821 =  ( n5820 ) == ( bv_8_170_n77 )  ;
assign n5822 = state_in[7:0] ;
assign n5823 =  ( n5822 ) == ( bv_8_169_n109 )  ;
assign n5824 = state_in[7:0] ;
assign n5825 =  ( n5824 ) == ( bv_8_168_n13 )  ;
assign n5826 = state_in[7:0] ;
assign n5827 =  ( n5826 ) == ( bv_8_167_n325 )  ;
assign n5828 = state_in[7:0] ;
assign n5829 =  ( n5828 ) == ( bv_8_166_n328 )  ;
assign n5830 = state_in[7:0] ;
assign n5831 =  ( n5830 ) == ( bv_8_165_n69 )  ;
assign n5832 = state_in[7:0] ;
assign n5833 =  ( n5832 ) == ( bv_8_164_n335 )  ;
assign n5834 = state_in[7:0] ;
assign n5835 =  ( n5834 ) == ( bv_8_163_n339 )  ;
assign n5836 = state_in[7:0] ;
assign n5837 =  ( n5836 ) == ( bv_8_162_n343 )  ;
assign n5838 = state_in[7:0] ;
assign n5839 =  ( n5838 ) == ( bv_8_161_n211 )  ;
assign n5840 = state_in[7:0] ;
assign n5841 =  ( n5840 ) == ( bv_8_160_n350 )  ;
assign n5842 = state_in[7:0] ;
assign n5843 =  ( n5842 ) == ( bv_8_159_n323 )  ;
assign n5844 = state_in[7:0] ;
assign n5845 =  ( n5844 ) == ( bv_8_158_n355 )  ;
assign n5846 = state_in[7:0] ;
assign n5847 =  ( n5846 ) == ( bv_8_157_n359 )  ;
assign n5848 = state_in[7:0] ;
assign n5849 =  ( n5848 ) == ( bv_8_156_n279 )  ;
assign n5850 = state_in[7:0] ;
assign n5851 =  ( n5850 ) == ( bv_8_155_n364 )  ;
assign n5852 = state_in[7:0] ;
assign n5853 =  ( n5852 ) == ( bv_8_154_n368 )  ;
assign n5854 = state_in[7:0] ;
assign n5855 =  ( n5854 ) == ( bv_8_153_n140 )  ;
assign n5856 = state_in[7:0] ;
assign n5857 =  ( n5856 ) == ( bv_8_152_n374 )  ;
assign n5858 = state_in[7:0] ;
assign n5859 =  ( n5858 ) == ( bv_8_151_n218 )  ;
assign n5860 = state_in[7:0] ;
assign n5861 =  ( n5860 ) == ( bv_8_150_n201 )  ;
assign n5862 = state_in[7:0] ;
assign n5863 =  ( n5862 ) == ( bv_8_149_n384 )  ;
assign n5864 = state_in[7:0] ;
assign n5865 =  ( n5864 ) == ( bv_8_148_n388 )  ;
assign n5866 = state_in[7:0] ;
assign n5867 =  ( n5866 ) == ( bv_8_147_n392 )  ;
assign n5868 = state_in[7:0] ;
assign n5869 =  ( n5868 ) == ( bv_8_146_n337 )  ;
assign n5870 = state_in[7:0] ;
assign n5871 =  ( n5870 ) == ( bv_8_145_n397 )  ;
assign n5872 = state_in[7:0] ;
assign n5873 =  ( n5872 ) == ( bv_8_144_n173 )  ;
assign n5874 = state_in[7:0] ;
assign n5875 =  ( n5874 ) == ( bv_8_143_n403 )  ;
assign n5876 = state_in[7:0] ;
assign n5877 =  ( n5876 ) == ( bv_8_142_n406 )  ;
assign n5878 = state_in[7:0] ;
assign n5879 =  ( n5878 ) == ( bv_8_141_n410 )  ;
assign n5880 = state_in[7:0] ;
assign n5881 =  ( n5880 ) == ( bv_8_140_n376 )  ;
assign n5882 = state_in[7:0] ;
assign n5883 =  ( n5882 ) == ( bv_8_139_n297 )  ;
assign n5884 = state_in[7:0] ;
assign n5885 =  ( n5884 ) == ( bv_8_138_n418 )  ;
assign n5886 = state_in[7:0] ;
assign n5887 =  ( n5886 ) == ( bv_8_137_n421 )  ;
assign n5888 = state_in[7:0] ;
assign n5889 =  ( n5888 ) == ( bv_8_136_n425 )  ;
assign n5890 = state_in[7:0] ;
assign n5891 =  ( n5890 ) == ( bv_8_135_n81 )  ;
assign n5892 = state_in[7:0] ;
assign n5893 =  ( n5892 ) == ( bv_8_134_n431 )  ;
assign n5894 = state_in[7:0] ;
assign n5895 =  ( n5894 ) == ( bv_8_133_n434 )  ;
assign n5896 = state_in[7:0] ;
assign n5897 =  ( n5896 ) == ( bv_8_132_n41 )  ;
assign n5898 = state_in[7:0] ;
assign n5899 =  ( n5898 ) == ( bv_8_131_n440 )  ;
assign n5900 = state_in[7:0] ;
assign n5901 =  ( n5900 ) == ( bv_8_130_n33 )  ;
assign n5902 = state_in[7:0] ;
assign n5903 =  ( n5902 ) == ( bv_8_129_n446 )  ;
assign n5904 = state_in[7:0] ;
assign n5905 =  ( n5904 ) == ( bv_8_128_n450 )  ;
assign n5906 = state_in[7:0] ;
assign n5907 =  ( n5906 ) == ( bv_8_127_n453 )  ;
assign n5908 = state_in[7:0] ;
assign n5909 =  ( n5908 ) == ( bv_8_126_n456 )  ;
assign n5910 = state_in[7:0] ;
assign n5911 =  ( n5910 ) == ( bv_8_125_n459 )  ;
assign n5912 = state_in[7:0] ;
assign n5913 =  ( n5912 ) == ( bv_8_124_n184 )  ;
assign n5914 = state_in[7:0] ;
assign n5915 =  ( n5914 ) == ( bv_8_123_n17 )  ;
assign n5916 = state_in[7:0] ;
assign n5917 =  ( n5916 ) == ( bv_8_122_n416 )  ;
assign n5918 = state_in[7:0] ;
assign n5919 =  ( n5918 ) == ( bv_8_121_n470 )  ;
assign n5920 = state_in[7:0] ;
assign n5921 =  ( n5920 ) == ( bv_8_120_n474 )  ;
assign n5922 = state_in[7:0] ;
assign n5923 =  ( n5922 ) == ( bv_8_119_n472 )  ;
assign n5924 = state_in[7:0] ;
assign n5925 =  ( n5924 ) == ( bv_8_118_n480 )  ;
assign n5926 = state_in[7:0] ;
assign n5927 =  ( n5926 ) == ( bv_8_117_n484 )  ;
assign n5928 = state_in[7:0] ;
assign n5929 =  ( n5928 ) == ( bv_8_116_n345 )  ;
assign n5930 = state_in[7:0] ;
assign n5931 =  ( n5930 ) == ( bv_8_115_n222 )  ;
assign n5932 = state_in[7:0] ;
assign n5933 =  ( n5932 ) == ( bv_8_114_n494 )  ;
assign n5934 = state_in[7:0] ;
assign n5935 =  ( n5934 ) == ( bv_8_113_n180 )  ;
assign n5936 = state_in[7:0] ;
assign n5937 =  ( n5936 ) == ( bv_8_112_n482 )  ;
assign n5938 = state_in[7:0] ;
assign n5939 =  ( n5938 ) == ( bv_8_111_n244 )  ;
assign n5940 = state_in[7:0] ;
assign n5941 =  ( n5940 ) == ( bv_8_110_n294 )  ;
assign n5942 = state_in[7:0] ;
assign n5943 =  ( n5942 ) == ( bv_8_109_n9 )  ;
assign n5944 = state_in[7:0] ;
assign n5945 =  ( n5944 ) == ( bv_8_108_n510 )  ;
assign n5946 = state_in[7:0] ;
assign n5947 =  ( n5946 ) == ( bv_8_107_n370 )  ;
assign n5948 = state_in[7:0] ;
assign n5949 =  ( n5948 ) == ( bv_8_106_n155 )  ;
assign n5950 = state_in[7:0] ;
assign n5951 =  ( n5950 ) == ( bv_8_105_n148 )  ;
assign n5952 = state_in[7:0] ;
assign n5953 =  ( n5952 ) == ( bv_8_104_n520 )  ;
assign n5954 = state_in[7:0] ;
assign n5955 =  ( n5954 ) == ( bv_8_103_n523 )  ;
assign n5956 = state_in[7:0] ;
assign n5957 =  ( n5956 ) == ( bv_8_102_n527 )  ;
assign n5958 = state_in[7:0] ;
assign n5959 =  ( n5958 ) == ( bv_8_101_n49 )  ;
assign n5960 = state_in[7:0] ;
assign n5961 =  ( n5960 ) == ( bv_8_100_n348 )  ;
assign n5962 = state_in[7:0] ;
assign n5963 =  ( n5962 ) == ( bv_8_99_n476 )  ;
assign n5964 = state_in[7:0] ;
assign n5965 =  ( n5964 ) == ( bv_8_98_n536 )  ;
assign n5966 = state_in[7:0] ;
assign n5967 =  ( n5966 ) == ( bv_8_97_n198 )  ;
assign n5968 = state_in[7:0] ;
assign n5969 =  ( n5968 ) == ( bv_8_96_n542 )  ;
assign n5970 = state_in[7:0] ;
assign n5971 =  ( n5970 ) == ( bv_8_95_n545 )  ;
assign n5972 = state_in[7:0] ;
assign n5973 =  ( n5972 ) == ( bv_8_94_n548 )  ;
assign n5974 = state_in[7:0] ;
assign n5975 =  ( n5974 ) == ( bv_8_93_n498 )  ;
assign n5976 = state_in[7:0] ;
assign n5977 =  ( n5976 ) == ( bv_8_92_n234 )  ;
assign n5978 = state_in[7:0] ;
assign n5979 =  ( n5978 ) == ( bv_8_91_n555 )  ;
assign n5980 = state_in[7:0] ;
assign n5981 =  ( n5980 ) == ( bv_8_90_n25 )  ;
assign n5982 = state_in[7:0] ;
assign n5983 =  ( n5982 ) == ( bv_8_89_n61 )  ;
assign n5984 = state_in[7:0] ;
assign n5985 =  ( n5984 ) == ( bv_8_88_n562 )  ;
assign n5986 = state_in[7:0] ;
assign n5987 =  ( n5986 ) == ( bv_8_87_n226 )  ;
assign n5988 = state_in[7:0] ;
assign n5989 =  ( n5988 ) == ( bv_8_86_n567 )  ;
assign n5990 = state_in[7:0] ;
assign n5991 =  ( n5990 ) == ( bv_8_85_n423 )  ;
assign n5992 = state_in[7:0] ;
assign n5993 =  ( n5992 ) == ( bv_8_84_n386 )  ;
assign n5994 = state_in[7:0] ;
assign n5995 =  ( n5994 ) == ( bv_8_83_n575 )  ;
assign n5996 = state_in[7:0] ;
assign n5997 =  ( n5996 ) == ( bv_8_82_n578 )  ;
assign n5998 = state_in[7:0] ;
assign n5999 =  ( n5998 ) == ( bv_8_81_n582 )  ;
assign n6000 = state_in[7:0] ;
assign n6001 =  ( n6000 ) == ( bv_8_80_n73 )  ;
assign n6002 = state_in[7:0] ;
assign n6003 =  ( n6002 ) == ( bv_8_79_n538 )  ;
assign n6004 = state_in[7:0] ;
assign n6005 =  ( n6004 ) == ( bv_8_78_n590 )  ;
assign n6006 = state_in[7:0] ;
assign n6007 =  ( n6006 ) == ( bv_8_77_n593 )  ;
assign n6008 = state_in[7:0] ;
assign n6009 =  ( n6008 ) == ( bv_8_76_n596 )  ;
assign n6010 = state_in[7:0] ;
assign n6011 =  ( n6010 ) == ( bv_8_75_n503 )  ;
assign n6012 = state_in[7:0] ;
assign n6013 =  ( n6012 ) == ( bv_8_74_n237 )  ;
assign n6014 = state_in[7:0] ;
assign n6015 =  ( n6014 ) == ( bv_8_73_n275 )  ;
assign n6016 = state_in[7:0] ;
assign n6017 =  ( n6016 ) == ( bv_8_72_n330 )  ;
assign n6018 = state_in[7:0] ;
assign n6019 =  ( n6018 ) == ( bv_8_71_n252 )  ;
assign n6020 = state_in[7:0] ;
assign n6021 =  ( n6020 ) == ( bv_8_70_n609 )  ;
assign n6022 = state_in[7:0] ;
assign n6023 =  ( n6022 ) == ( bv_8_69_n612 )  ;
assign n6024 = state_in[7:0] ;
assign n6025 =  ( n6024 ) == ( bv_8_68_n390 )  ;
assign n6026 = state_in[7:0] ;
assign n6027 =  ( n6026 ) == ( bv_8_67_n318 )  ;
assign n6028 = state_in[7:0] ;
assign n6029 =  ( n6028 ) == ( bv_8_66_n466 )  ;
assign n6030 = state_in[7:0] ;
assign n6031 =  ( n6030 ) == ( bv_8_65_n623 )  ;
assign n6032 = state_in[7:0] ;
assign n6033 =  ( n6032 ) == ( bv_8_64_n573 )  ;
assign n6034 = state_in[7:0] ;
assign n6035 =  ( n6034 ) == ( bv_8_63_n489 )  ;
assign n6036 = state_in[7:0] ;
assign n6037 =  ( n6036 ) == ( bv_8_62_n205 )  ;
assign n6038 = state_in[7:0] ;
assign n6039 =  ( n6038 ) == ( bv_8_61_n634 )  ;
assign n6040 = state_in[7:0] ;
assign n6041 =  ( n6040 ) == ( bv_8_60_n93 )  ;
assign n6042 = state_in[7:0] ;
assign n6043 =  ( n6042 ) == ( bv_8_59_n382 )  ;
assign n6044 = state_in[7:0] ;
assign n6045 =  ( n6044 ) == ( bv_8_58_n136 )  ;
assign n6046 = state_in[7:0] ;
assign n6047 =  ( n6046 ) == ( bv_8_57_n312 )  ;
assign n6048 = state_in[7:0] ;
assign n6049 =  ( n6048 ) == ( bv_8_56_n230 )  ;
assign n6050 = state_in[7:0] ;
assign n6051 =  ( n6050 ) == ( bv_8_55_n650 )  ;
assign n6052 = state_in[7:0] ;
assign n6053 =  ( n6052 ) == ( bv_8_54_n616 )  ;
assign n6054 = state_in[7:0] ;
assign n6055 =  ( n6054 ) == ( bv_8_53_n436 )  ;
assign n6056 = state_in[7:0] ;
assign n6057 =  ( n6056 ) == ( bv_8_52_n619 )  ;
assign n6058 = state_in[7:0] ;
assign n6059 =  ( n6058 ) == ( bv_8_51_n101 )  ;
assign n6060 = state_in[7:0] ;
assign n6061 =  ( n6060 ) == ( bv_8_50_n408 )  ;
assign n6062 = state_in[7:0] ;
assign n6063 =  ( n6062 ) == ( bv_8_49_n309 )  ;
assign n6064 = state_in[7:0] ;
assign n6065 =  ( n6064 ) == ( bv_8_48_n660 )  ;
assign n6066 = state_in[7:0] ;
assign n6067 =  ( n6066 ) == ( bv_8_47_n652 )  ;
assign n6068 = state_in[7:0] ;
assign n6069 =  ( n6068 ) == ( bv_8_46_n429 )  ;
assign n6070 = state_in[7:0] ;
assign n6071 =  ( n6070 ) == ( bv_8_45_n97 )  ;
assign n6072 = state_in[7:0] ;
assign n6073 =  ( n6072 ) == ( bv_8_44_n5 )  ;
assign n6074 = state_in[7:0] ;
assign n6075 =  ( n6074 ) == ( bv_8_43_n121 )  ;
assign n6076 = state_in[7:0] ;
assign n6077 =  ( n6076 ) == ( bv_8_42_n672 )  ;
assign n6078 = state_in[7:0] ;
assign n6079 =  ( n6078 ) == ( bv_8_41_n29 )  ;
assign n6080 = state_in[7:0] ;
assign n6081 =  ( n6080 ) == ( bv_8_40_n366 )  ;
assign n6082 = state_in[7:0] ;
assign n6083 =  ( n6082 ) == ( bv_8_39_n132 )  ;
assign n6084 = state_in[7:0] ;
assign n6085 =  ( n6084 ) == ( bv_8_38_n444 )  ;
assign n6086 = state_in[7:0] ;
assign n6087 =  ( n6086 ) == ( bv_8_37_n506 )  ;
assign n6088 = state_in[7:0] ;
assign n6089 =  ( n6088 ) == ( bv_8_36_n645 )  ;
assign n6090 = state_in[7:0] ;
assign n6091 =  ( n6090 ) == ( bv_8_35_n696 )  ;
assign n6092 = state_in[7:0] ;
assign n6093 =  ( n6092 ) == ( bv_8_34_n117 )  ;
assign n6094 = state_in[7:0] ;
assign n6095 =  ( n6094 ) == ( bv_8_33_n486 )  ;
assign n6096 = state_in[7:0] ;
assign n6097 =  ( n6096 ) == ( bv_8_32_n463 )  ;
assign n6098 = state_in[7:0] ;
assign n6099 =  ( n6098 ) == ( bv_8_31_n705 )  ;
assign n6100 = state_in[7:0] ;
assign n6101 =  ( n6100 ) == ( bv_8_30_n21 )  ;
assign n6102 = state_in[7:0] ;
assign n6103 =  ( n6102 ) == ( bv_8_29_n625 )  ;
assign n6104 = state_in[7:0] ;
assign n6105 =  ( n6104 ) == ( bv_8_28_n162 )  ;
assign n6106 = state_in[7:0] ;
assign n6107 =  ( n6106 ) == ( bv_8_27_n642 )  ;
assign n6108 = state_in[7:0] ;
assign n6109 =  ( n6108 ) == ( bv_8_26_n53 )  ;
assign n6110 = state_in[7:0] ;
assign n6111 =  ( n6110 ) == ( bv_8_25_n399 )  ;
assign n6112 = state_in[7:0] ;
assign n6113 =  ( n6112 ) == ( bv_8_24_n448 )  ;
assign n6114 = state_in[7:0] ;
assign n6115 =  ( n6114 ) == ( bv_8_23_n144 )  ;
assign n6116 = state_in[7:0] ;
assign n6117 =  ( n6116 ) == ( bv_8_22_n357 )  ;
assign n6118 = state_in[7:0] ;
assign n6119 =  ( n6118 ) == ( bv_8_21_n89 )  ;
assign n6120 = state_in[7:0] ;
assign n6121 =  ( n6120 ) == ( bv_8_20_n341 )  ;
assign n6122 = state_in[7:0] ;
assign n6123 =  ( n6122 ) == ( bv_8_19_n588 )  ;
assign n6124 = state_in[7:0] ;
assign n6125 =  ( n6124 ) == ( bv_8_18_n628 )  ;
assign n6126 = state_in[7:0] ;
assign n6127 =  ( n6126 ) == ( bv_8_17_n525 )  ;
assign n6128 = state_in[7:0] ;
assign n6129 =  ( n6128 ) == ( bv_8_16_n248 )  ;
assign n6130 = state_in[7:0] ;
assign n6131 =  ( n6130 ) == ( bv_8_15_n190 )  ;
assign n6132 = state_in[7:0] ;
assign n6133 =  ( n6132 ) == ( bv_8_14_n648 )  ;
assign n6134 = state_in[7:0] ;
assign n6135 =  ( n6134 ) == ( bv_8_13_n194 )  ;
assign n6136 = state_in[7:0] ;
assign n6137 =  ( n6136 ) == ( bv_8_12_n333 )  ;
assign n6138 = state_in[7:0] ;
assign n6139 =  ( n6138 ) == ( bv_8_11_n379 )  ;
assign n6140 = state_in[7:0] ;
assign n6141 =  ( n6140 ) == ( bv_8_10_n655 )  ;
assign n6142 = state_in[7:0] ;
assign n6143 =  ( n6142 ) == ( bv_8_9_n57 )  ;
assign n6144 = state_in[7:0] ;
assign n6145 =  ( n6144 ) == ( bv_8_8_n669 )  ;
assign n6146 = state_in[7:0] ;
assign n6147 =  ( n6146 ) == ( bv_8_7_n105 )  ;
assign n6148 = state_in[7:0] ;
assign n6149 =  ( n6148 ) == ( bv_8_6_n169 )  ;
assign n6150 = state_in[7:0] ;
assign n6151 =  ( n6150 ) == ( bv_8_5_n492 )  ;
assign n6152 = state_in[7:0] ;
assign n6153 =  ( n6152 ) == ( bv_8_4_n516 )  ;
assign n6154 = state_in[7:0] ;
assign n6155 =  ( n6154 ) == ( bv_8_3_n65 )  ;
assign n6156 = state_in[7:0] ;
assign n6157 =  ( n6156 ) == ( bv_8_2_n751 )  ;
assign n6158 = state_in[7:0] ;
assign n6159 =  ( n6158 ) == ( bv_8_1_n287 )  ;
assign n6160 = state_in[7:0] ;
assign n6161 =  ( n6160 ) == ( bv_8_0_n580 )  ;
assign n6162 =  ( n6161 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n6163 =  ( n6159 ) ? ( bv_8_248_n31 ) : ( n6162 ) ;
assign n6164 =  ( n6157 ) ? ( bv_8_238_n71 ) : ( n6163 ) ;
assign n6165 =  ( n6155 ) ? ( bv_8_246_n39 ) : ( n6164 ) ;
assign n6166 =  ( n6153 ) ? ( bv_8_255_n3 ) : ( n6165 ) ;
assign n6167 =  ( n6151 ) ? ( bv_8_214_n164 ) : ( n6166 ) ;
assign n6168 =  ( n6149 ) ? ( bv_8_222_n134 ) : ( n6167 ) ;
assign n6169 =  ( n6147 ) ? ( bv_8_145_n397 ) : ( n6168 ) ;
assign n6170 =  ( n6145 ) ? ( bv_8_96_n542 ) : ( n6169 ) ;
assign n6171 =  ( n6143 ) ? ( bv_8_2_n751 ) : ( n6170 ) ;
assign n6172 =  ( n6141 ) ? ( bv_8_206_n192 ) : ( n6171 ) ;
assign n6173 =  ( n6139 ) ? ( bv_8_86_n567 ) : ( n6172 ) ;
assign n6174 =  ( n6137 ) ? ( bv_8_231_n99 ) : ( n6173 ) ;
assign n6175 =  ( n6135 ) ? ( bv_8_181_n281 ) : ( n6174 ) ;
assign n6176 =  ( n6133 ) ? ( bv_8_77_n593 ) : ( n6175 ) ;
assign n6177 =  ( n6131 ) ? ( bv_8_236_n79 ) : ( n6176 ) ;
assign n6178 =  ( n6129 ) ? ( bv_8_143_n403 ) : ( n6177 ) ;
assign n6179 =  ( n6127 ) ? ( bv_8_31_n705 ) : ( n6178 ) ;
assign n6180 =  ( n6125 ) ? ( bv_8_137_n421 ) : ( n6179 ) ;
assign n6181 =  ( n6123 ) ? ( bv_8_250_n23 ) : ( n6180 ) ;
assign n6182 =  ( n6121 ) ? ( bv_8_239_n67 ) : ( n6181 ) ;
assign n6183 =  ( n6119 ) ? ( bv_8_178_n292 ) : ( n6182 ) ;
assign n6184 =  ( n6117 ) ? ( bv_8_142_n406 ) : ( n6183 ) ;
assign n6185 =  ( n6115 ) ? ( bv_8_251_n19 ) : ( n6184 ) ;
assign n6186 =  ( n6113 ) ? ( bv_8_65_n623 ) : ( n6185 ) ;
assign n6187 =  ( n6111 ) ? ( bv_8_179_n289 ) : ( n6186 ) ;
assign n6188 =  ( n6109 ) ? ( bv_8_95_n545 ) : ( n6187 ) ;
assign n6189 =  ( n6107 ) ? ( bv_8_69_n612 ) : ( n6188 ) ;
assign n6190 =  ( n6105 ) ? ( bv_8_35_n696 ) : ( n6189 ) ;
assign n6191 =  ( n6103 ) ? ( bv_8_83_n575 ) : ( n6190 ) ;
assign n6192 =  ( n6101 ) ? ( bv_8_228_n111 ) : ( n6191 ) ;
assign n6193 =  ( n6099 ) ? ( bv_8_155_n364 ) : ( n6192 ) ;
assign n6194 =  ( n6097 ) ? ( bv_8_117_n484 ) : ( n6193 ) ;
assign n6195 =  ( n6095 ) ? ( bv_8_225_n123 ) : ( n6194 ) ;
assign n6196 =  ( n6093 ) ? ( bv_8_61_n634 ) : ( n6195 ) ;
assign n6197 =  ( n6091 ) ? ( bv_8_76_n596 ) : ( n6196 ) ;
assign n6198 =  ( n6089 ) ? ( bv_8_108_n510 ) : ( n6197 ) ;
assign n6199 =  ( n6087 ) ? ( bv_8_126_n456 ) : ( n6198 ) ;
assign n6200 =  ( n6085 ) ? ( bv_8_245_n43 ) : ( n6199 ) ;
assign n6201 =  ( n6083 ) ? ( bv_8_131_n440 ) : ( n6200 ) ;
assign n6202 =  ( n6081 ) ? ( bv_8_104_n520 ) : ( n6201 ) ;
assign n6203 =  ( n6079 ) ? ( bv_8_81_n582 ) : ( n6202 ) ;
assign n6204 =  ( n6077 ) ? ( bv_8_209_n182 ) : ( n6203 ) ;
assign n6205 =  ( n6075 ) ? ( bv_8_249_n27 ) : ( n6204 ) ;
assign n6206 =  ( n6073 ) ? ( bv_8_226_n119 ) : ( n6205 ) ;
assign n6207 =  ( n6071 ) ? ( bv_8_171_n314 ) : ( n6206 ) ;
assign n6208 =  ( n6069 ) ? ( bv_8_98_n536 ) : ( n6207 ) ;
assign n6209 =  ( n6067 ) ? ( bv_8_42_n672 ) : ( n6208 ) ;
assign n6210 =  ( n6065 ) ? ( bv_8_8_n669 ) : ( n6209 ) ;
assign n6211 =  ( n6063 ) ? ( bv_8_149_n384 ) : ( n6210 ) ;
assign n6212 =  ( n6061 ) ? ( bv_8_70_n609 ) : ( n6211 ) ;
assign n6213 =  ( n6059 ) ? ( bv_8_157_n359 ) : ( n6212 ) ;
assign n6214 =  ( n6057 ) ? ( bv_8_48_n660 ) : ( n6213 ) ;
assign n6215 =  ( n6055 ) ? ( bv_8_55_n650 ) : ( n6214 ) ;
assign n6216 =  ( n6053 ) ? ( bv_8_10_n655 ) : ( n6215 ) ;
assign n6217 =  ( n6051 ) ? ( bv_8_47_n652 ) : ( n6216 ) ;
assign n6218 =  ( n6049 ) ? ( bv_8_14_n648 ) : ( n6217 ) ;
assign n6219 =  ( n6047 ) ? ( bv_8_36_n645 ) : ( n6218 ) ;
assign n6220 =  ( n6045 ) ? ( bv_8_27_n642 ) : ( n6219 ) ;
assign n6221 =  ( n6043 ) ? ( bv_8_223_n130 ) : ( n6220 ) ;
assign n6222 =  ( n6041 ) ? ( bv_8_205_n196 ) : ( n6221 ) ;
assign n6223 =  ( n6039 ) ? ( bv_8_78_n590 ) : ( n6222 ) ;
assign n6224 =  ( n6037 ) ? ( bv_8_127_n453 ) : ( n6223 ) ;
assign n6225 =  ( n6035 ) ? ( bv_8_234_n87 ) : ( n6224 ) ;
assign n6226 =  ( n6033 ) ? ( bv_8_18_n628 ) : ( n6225 ) ;
assign n6227 =  ( n6031 ) ? ( bv_8_29_n625 ) : ( n6226 ) ;
assign n6228 =  ( n6029 ) ? ( bv_8_88_n562 ) : ( n6227 ) ;
assign n6229 =  ( n6027 ) ? ( bv_8_52_n619 ) : ( n6228 ) ;
assign n6230 =  ( n6025 ) ? ( bv_8_54_n616 ) : ( n6229 ) ;
assign n6231 =  ( n6023 ) ? ( bv_8_220_n142 ) : ( n6230 ) ;
assign n6232 =  ( n6021 ) ? ( bv_8_180_n285 ) : ( n6231 ) ;
assign n6233 =  ( n6019 ) ? ( bv_8_91_n555 ) : ( n6232 ) ;
assign n6234 =  ( n6017 ) ? ( bv_8_164_n335 ) : ( n6233 ) ;
assign n6235 =  ( n6015 ) ? ( bv_8_118_n480 ) : ( n6234 ) ;
assign n6236 =  ( n6013 ) ? ( bv_8_183_n273 ) : ( n6235 ) ;
assign n6237 =  ( n6011 ) ? ( bv_8_125_n459 ) : ( n6236 ) ;
assign n6238 =  ( n6009 ) ? ( bv_8_82_n578 ) : ( n6237 ) ;
assign n6239 =  ( n6007 ) ? ( bv_8_221_n138 ) : ( n6238 ) ;
assign n6240 =  ( n6005 ) ? ( bv_8_94_n548 ) : ( n6239 ) ;
assign n6241 =  ( n6003 ) ? ( bv_8_19_n588 ) : ( n6240 ) ;
assign n6242 =  ( n6001 ) ? ( bv_8_166_n328 ) : ( n6241 ) ;
assign n6243 =  ( n5999 ) ? ( bv_8_185_n266 ) : ( n6242 ) ;
assign n6244 =  ( n5997 ) ? ( bv_8_0_n580 ) : ( n6243 ) ;
assign n6245 =  ( n5995 ) ? ( bv_8_193_n239 ) : ( n6244 ) ;
assign n6246 =  ( n5993 ) ? ( bv_8_64_n573 ) : ( n6245 ) ;
assign n6247 =  ( n5991 ) ? ( bv_8_227_n115 ) : ( n6246 ) ;
assign n6248 =  ( n5989 ) ? ( bv_8_121_n470 ) : ( n6247 ) ;
assign n6249 =  ( n5987 ) ? ( bv_8_182_n277 ) : ( n6248 ) ;
assign n6250 =  ( n5985 ) ? ( bv_8_212_n171 ) : ( n6249 ) ;
assign n6251 =  ( n5983 ) ? ( bv_8_141_n410 ) : ( n6250 ) ;
assign n6252 =  ( n5981 ) ? ( bv_8_103_n523 ) : ( n6251 ) ;
assign n6253 =  ( n5979 ) ? ( bv_8_114_n494 ) : ( n6252 ) ;
assign n6254 =  ( n5977 ) ? ( bv_8_148_n388 ) : ( n6253 ) ;
assign n6255 =  ( n5975 ) ? ( bv_8_152_n374 ) : ( n6254 ) ;
assign n6256 =  ( n5973 ) ? ( bv_8_176_n299 ) : ( n6255 ) ;
assign n6257 =  ( n5971 ) ? ( bv_8_133_n434 ) : ( n6256 ) ;
assign n6258 =  ( n5969 ) ? ( bv_8_187_n260 ) : ( n6257 ) ;
assign n6259 =  ( n5967 ) ? ( bv_8_197_n224 ) : ( n6258 ) ;
assign n6260 =  ( n5965 ) ? ( bv_8_79_n538 ) : ( n6259 ) ;
assign n6261 =  ( n5963 ) ? ( bv_8_237_n75 ) : ( n6260 ) ;
assign n6262 =  ( n5961 ) ? ( bv_8_134_n431 ) : ( n6261 ) ;
assign n6263 =  ( n5959 ) ? ( bv_8_154_n368 ) : ( n6262 ) ;
assign n6264 =  ( n5957 ) ? ( bv_8_102_n527 ) : ( n6263 ) ;
assign n6265 =  ( n5955 ) ? ( bv_8_17_n525 ) : ( n6264 ) ;
assign n6266 =  ( n5953 ) ? ( bv_8_138_n418 ) : ( n6265 ) ;
assign n6267 =  ( n5951 ) ? ( bv_8_233_n91 ) : ( n6266 ) ;
assign n6268 =  ( n5949 ) ? ( bv_8_4_n516 ) : ( n6267 ) ;
assign n6269 =  ( n5947 ) ? ( bv_8_254_n7 ) : ( n6268 ) ;
assign n6270 =  ( n5945 ) ? ( bv_8_160_n350 ) : ( n6269 ) ;
assign n6271 =  ( n5943 ) ? ( bv_8_120_n474 ) : ( n6270 ) ;
assign n6272 =  ( n5941 ) ? ( bv_8_37_n506 ) : ( n6271 ) ;
assign n6273 =  ( n5939 ) ? ( bv_8_75_n503 ) : ( n6272 ) ;
assign n6274 =  ( n5937 ) ? ( bv_8_162_n343 ) : ( n6273 ) ;
assign n6275 =  ( n5935 ) ? ( bv_8_93_n498 ) : ( n6274 ) ;
assign n6276 =  ( n5933 ) ? ( bv_8_128_n450 ) : ( n6275 ) ;
assign n6277 =  ( n5931 ) ? ( bv_8_5_n492 ) : ( n6276 ) ;
assign n6278 =  ( n5929 ) ? ( bv_8_63_n489 ) : ( n6277 ) ;
assign n6279 =  ( n5927 ) ? ( bv_8_33_n486 ) : ( n6278 ) ;
assign n6280 =  ( n5925 ) ? ( bv_8_112_n482 ) : ( n6279 ) ;
assign n6281 =  ( n5923 ) ? ( bv_8_241_n59 ) : ( n6280 ) ;
assign n6282 =  ( n5921 ) ? ( bv_8_99_n476 ) : ( n6281 ) ;
assign n6283 =  ( n5919 ) ? ( bv_8_119_n472 ) : ( n6282 ) ;
assign n6284 =  ( n5917 ) ? ( bv_8_175_n302 ) : ( n6283 ) ;
assign n6285 =  ( n5915 ) ? ( bv_8_66_n466 ) : ( n6284 ) ;
assign n6286 =  ( n5913 ) ? ( bv_8_32_n463 ) : ( n6285 ) ;
assign n6287 =  ( n5911 ) ? ( bv_8_229_n107 ) : ( n6286 ) ;
assign n6288 =  ( n5909 ) ? ( bv_8_253_n11 ) : ( n6287 ) ;
assign n6289 =  ( n5907 ) ? ( bv_8_191_n246 ) : ( n6288 ) ;
assign n6290 =  ( n5905 ) ? ( bv_8_129_n446 ) : ( n6289 ) ;
assign n6291 =  ( n5903 ) ? ( bv_8_24_n448 ) : ( n6290 ) ;
assign n6292 =  ( n5901 ) ? ( bv_8_38_n444 ) : ( n6291 ) ;
assign n6293 =  ( n5899 ) ? ( bv_8_195_n232 ) : ( n6292 ) ;
assign n6294 =  ( n5897 ) ? ( bv_8_190_n250 ) : ( n6293 ) ;
assign n6295 =  ( n5895 ) ? ( bv_8_53_n436 ) : ( n6294 ) ;
assign n6296 =  ( n5893 ) ? ( bv_8_136_n425 ) : ( n6295 ) ;
assign n6297 =  ( n5891 ) ? ( bv_8_46_n429 ) : ( n6296 ) ;
assign n6298 =  ( n5889 ) ? ( bv_8_147_n392 ) : ( n6297 ) ;
assign n6299 =  ( n5887 ) ? ( bv_8_85_n423 ) : ( n6298 ) ;
assign n6300 =  ( n5885 ) ? ( bv_8_252_n15 ) : ( n6299 ) ;
assign n6301 =  ( n5883 ) ? ( bv_8_122_n416 ) : ( n6300 ) ;
assign n6302 =  ( n5881 ) ? ( bv_8_200_n213 ) : ( n6301 ) ;
assign n6303 =  ( n5879 ) ? ( bv_8_186_n263 ) : ( n6302 ) ;
assign n6304 =  ( n5877 ) ? ( bv_8_50_n408 ) : ( n6303 ) ;
assign n6305 =  ( n5875 ) ? ( bv_8_230_n103 ) : ( n6304 ) ;
assign n6306 =  ( n5873 ) ? ( bv_8_192_n242 ) : ( n6305 ) ;
assign n6307 =  ( n5871 ) ? ( bv_8_25_n399 ) : ( n6306 ) ;
assign n6308 =  ( n5869 ) ? ( bv_8_158_n355 ) : ( n6307 ) ;
assign n6309 =  ( n5867 ) ? ( bv_8_163_n339 ) : ( n6308 ) ;
assign n6310 =  ( n5865 ) ? ( bv_8_68_n390 ) : ( n6309 ) ;
assign n6311 =  ( n5863 ) ? ( bv_8_84_n386 ) : ( n6310 ) ;
assign n6312 =  ( n5861 ) ? ( bv_8_59_n382 ) : ( n6311 ) ;
assign n6313 =  ( n5859 ) ? ( bv_8_11_n379 ) : ( n6312 ) ;
assign n6314 =  ( n5857 ) ? ( bv_8_140_n376 ) : ( n6313 ) ;
assign n6315 =  ( n5855 ) ? ( bv_8_199_n216 ) : ( n6314 ) ;
assign n6316 =  ( n5853 ) ? ( bv_8_107_n370 ) : ( n6315 ) ;
assign n6317 =  ( n5851 ) ? ( bv_8_40_n366 ) : ( n6316 ) ;
assign n6318 =  ( n5849 ) ? ( bv_8_167_n325 ) : ( n6317 ) ;
assign n6319 =  ( n5847 ) ? ( bv_8_188_n257 ) : ( n6318 ) ;
assign n6320 =  ( n5845 ) ? ( bv_8_22_n357 ) : ( n6319 ) ;
assign n6321 =  ( n5843 ) ? ( bv_8_173_n307 ) : ( n6320 ) ;
assign n6322 =  ( n5841 ) ? ( bv_8_219_n146 ) : ( n6321 ) ;
assign n6323 =  ( n5839 ) ? ( bv_8_100_n348 ) : ( n6322 ) ;
assign n6324 =  ( n5837 ) ? ( bv_8_116_n345 ) : ( n6323 ) ;
assign n6325 =  ( n5835 ) ? ( bv_8_20_n341 ) : ( n6324 ) ;
assign n6326 =  ( n5833 ) ? ( bv_8_146_n337 ) : ( n6325 ) ;
assign n6327 =  ( n5831 ) ? ( bv_8_12_n333 ) : ( n6326 ) ;
assign n6328 =  ( n5829 ) ? ( bv_8_72_n330 ) : ( n6327 ) ;
assign n6329 =  ( n5827 ) ? ( bv_8_184_n270 ) : ( n6328 ) ;
assign n6330 =  ( n5825 ) ? ( bv_8_159_n323 ) : ( n6329 ) ;
assign n6331 =  ( n5823 ) ? ( bv_8_189_n254 ) : ( n6330 ) ;
assign n6332 =  ( n5821 ) ? ( bv_8_67_n318 ) : ( n6331 ) ;
assign n6333 =  ( n5819 ) ? ( bv_8_196_n228 ) : ( n6332 ) ;
assign n6334 =  ( n5817 ) ? ( bv_8_57_n312 ) : ( n6333 ) ;
assign n6335 =  ( n5815 ) ? ( bv_8_49_n309 ) : ( n6334 ) ;
assign n6336 =  ( n5813 ) ? ( bv_8_211_n175 ) : ( n6335 ) ;
assign n6337 =  ( n5811 ) ? ( bv_8_242_n55 ) : ( n6336 ) ;
assign n6338 =  ( n5809 ) ? ( bv_8_213_n167 ) : ( n6337 ) ;
assign n6339 =  ( n5807 ) ? ( bv_8_139_n297 ) : ( n6338 ) ;
assign n6340 =  ( n5805 ) ? ( bv_8_110_n294 ) : ( n6339 ) ;
assign n6341 =  ( n5803 ) ? ( bv_8_218_n150 ) : ( n6340 ) ;
assign n6342 =  ( n5801 ) ? ( bv_8_1_n287 ) : ( n6341 ) ;
assign n6343 =  ( n5799 ) ? ( bv_8_177_n283 ) : ( n6342 ) ;
assign n6344 =  ( n5797 ) ? ( bv_8_156_n279 ) : ( n6343 ) ;
assign n6345 =  ( n5795 ) ? ( bv_8_73_n275 ) : ( n6344 ) ;
assign n6346 =  ( n5793 ) ? ( bv_8_216_n157 ) : ( n6345 ) ;
assign n6347 =  ( n5791 ) ? ( bv_8_172_n268 ) : ( n6346 ) ;
assign n6348 =  ( n5789 ) ? ( bv_8_243_n51 ) : ( n6347 ) ;
assign n6349 =  ( n5787 ) ? ( bv_8_207_n188 ) : ( n6348 ) ;
assign n6350 =  ( n5785 ) ? ( bv_8_202_n207 ) : ( n6349 ) ;
assign n6351 =  ( n5783 ) ? ( bv_8_244_n47 ) : ( n6350 ) ;
assign n6352 =  ( n5781 ) ? ( bv_8_71_n252 ) : ( n6351 ) ;
assign n6353 =  ( n5779 ) ? ( bv_8_16_n248 ) : ( n6352 ) ;
assign n6354 =  ( n5777 ) ? ( bv_8_111_n244 ) : ( n6353 ) ;
assign n6355 =  ( n5775 ) ? ( bv_8_240_n63 ) : ( n6354 ) ;
assign n6356 =  ( n5773 ) ? ( bv_8_74_n237 ) : ( n6355 ) ;
assign n6357 =  ( n5771 ) ? ( bv_8_92_n234 ) : ( n6356 ) ;
assign n6358 =  ( n5769 ) ? ( bv_8_56_n230 ) : ( n6357 ) ;
assign n6359 =  ( n5767 ) ? ( bv_8_87_n226 ) : ( n6358 ) ;
assign n6360 =  ( n5765 ) ? ( bv_8_115_n222 ) : ( n6359 ) ;
assign n6361 =  ( n5763 ) ? ( bv_8_151_n218 ) : ( n6360 ) ;
assign n6362 =  ( n5761 ) ? ( bv_8_203_n203 ) : ( n6361 ) ;
assign n6363 =  ( n5759 ) ? ( bv_8_161_n211 ) : ( n6362 ) ;
assign n6364 =  ( n5757 ) ? ( bv_8_232_n95 ) : ( n6363 ) ;
assign n6365 =  ( n5755 ) ? ( bv_8_62_n205 ) : ( n6364 ) ;
assign n6366 =  ( n5753 ) ? ( bv_8_150_n201 ) : ( n6365 ) ;
assign n6367 =  ( n5751 ) ? ( bv_8_97_n198 ) : ( n6366 ) ;
assign n6368 =  ( n5749 ) ? ( bv_8_13_n194 ) : ( n6367 ) ;
assign n6369 =  ( n5747 ) ? ( bv_8_15_n190 ) : ( n6368 ) ;
assign n6370 =  ( n5745 ) ? ( bv_8_224_n126 ) : ( n6369 ) ;
assign n6371 =  ( n5743 ) ? ( bv_8_124_n184 ) : ( n6370 ) ;
assign n6372 =  ( n5741 ) ? ( bv_8_113_n180 ) : ( n6371 ) ;
assign n6373 =  ( n5739 ) ? ( bv_8_204_n177 ) : ( n6372 ) ;
assign n6374 =  ( n5737 ) ? ( bv_8_144_n173 ) : ( n6373 ) ;
assign n6375 =  ( n5735 ) ? ( bv_8_6_n169 ) : ( n6374 ) ;
assign n6376 =  ( n5733 ) ? ( bv_8_247_n35 ) : ( n6375 ) ;
assign n6377 =  ( n5731 ) ? ( bv_8_28_n162 ) : ( n6376 ) ;
assign n6378 =  ( n5729 ) ? ( bv_8_194_n159 ) : ( n6377 ) ;
assign n6379 =  ( n5727 ) ? ( bv_8_106_n155 ) : ( n6378 ) ;
assign n6380 =  ( n5725 ) ? ( bv_8_174_n152 ) : ( n6379 ) ;
assign n6381 =  ( n5723 ) ? ( bv_8_105_n148 ) : ( n6380 ) ;
assign n6382 =  ( n5721 ) ? ( bv_8_23_n144 ) : ( n6381 ) ;
assign n6383 =  ( n5719 ) ? ( bv_8_153_n140 ) : ( n6382 ) ;
assign n6384 =  ( n5717 ) ? ( bv_8_58_n136 ) : ( n6383 ) ;
assign n6385 =  ( n5715 ) ? ( bv_8_39_n132 ) : ( n6384 ) ;
assign n6386 =  ( n5713 ) ? ( bv_8_217_n128 ) : ( n6385 ) ;
assign n6387 =  ( n5711 ) ? ( bv_8_235_n83 ) : ( n6386 ) ;
assign n6388 =  ( n5709 ) ? ( bv_8_43_n121 ) : ( n6387 ) ;
assign n6389 =  ( n5707 ) ? ( bv_8_34_n117 ) : ( n6388 ) ;
assign n6390 =  ( n5705 ) ? ( bv_8_210_n113 ) : ( n6389 ) ;
assign n6391 =  ( n5703 ) ? ( bv_8_169_n109 ) : ( n6390 ) ;
assign n6392 =  ( n5701 ) ? ( bv_8_7_n105 ) : ( n6391 ) ;
assign n6393 =  ( n5699 ) ? ( bv_8_51_n101 ) : ( n6392 ) ;
assign n6394 =  ( n5697 ) ? ( bv_8_45_n97 ) : ( n6393 ) ;
assign n6395 =  ( n5695 ) ? ( bv_8_60_n93 ) : ( n6394 ) ;
assign n6396 =  ( n5693 ) ? ( bv_8_21_n89 ) : ( n6395 ) ;
assign n6397 =  ( n5691 ) ? ( bv_8_201_n85 ) : ( n6396 ) ;
assign n6398 =  ( n5689 ) ? ( bv_8_135_n81 ) : ( n6397 ) ;
assign n6399 =  ( n5687 ) ? ( bv_8_170_n77 ) : ( n6398 ) ;
assign n6400 =  ( n5685 ) ? ( bv_8_80_n73 ) : ( n6399 ) ;
assign n6401 =  ( n5683 ) ? ( bv_8_165_n69 ) : ( n6400 ) ;
assign n6402 =  ( n5681 ) ? ( bv_8_3_n65 ) : ( n6401 ) ;
assign n6403 =  ( n5679 ) ? ( bv_8_89_n61 ) : ( n6402 ) ;
assign n6404 =  ( n5677 ) ? ( bv_8_9_n57 ) : ( n6403 ) ;
assign n6405 =  ( n5675 ) ? ( bv_8_26_n53 ) : ( n6404 ) ;
assign n6406 =  ( n5673 ) ? ( bv_8_101_n49 ) : ( n6405 ) ;
assign n6407 =  ( n5671 ) ? ( bv_8_215_n45 ) : ( n6406 ) ;
assign n6408 =  ( n5669 ) ? ( bv_8_132_n41 ) : ( n6407 ) ;
assign n6409 =  ( n5667 ) ? ( bv_8_208_n37 ) : ( n6408 ) ;
assign n6410 =  ( n5665 ) ? ( bv_8_130_n33 ) : ( n6409 ) ;
assign n6411 =  ( n5663 ) ? ( bv_8_41_n29 ) : ( n6410 ) ;
assign n6412 =  ( n5661 ) ? ( bv_8_90_n25 ) : ( n6411 ) ;
assign n6413 =  ( n5659 ) ? ( bv_8_30_n21 ) : ( n6412 ) ;
assign n6414 =  ( n5657 ) ? ( bv_8_123_n17 ) : ( n6413 ) ;
assign n6415 =  ( n5655 ) ? ( bv_8_168_n13 ) : ( n6414 ) ;
assign n6416 =  ( n5653 ) ? ( bv_8_109_n9 ) : ( n6415 ) ;
assign n6417 =  ( n5651 ) ? ( bv_8_44_n5 ) : ( n6416 ) ;
assign n6418 =  ( n5649 ) ^ ( n6417 )  ;
assign n6419 = key[111:104] ;
assign n6420 =  ( n6418 ) ^ ( n6419 )  ;
assign n6421 =  { ( n5646 ) , ( n6420 ) }  ;
assign n6422 =  ( n4871 ) ^ ( n1025 )  ;
assign n6423 =  ( n6422 ) ^ ( n1793 )  ;
assign n6424 =  ( n6423 ) ^ ( n3331 )  ;
assign n6425 =  ( n6424 ) ^ ( n6417 )  ;
assign n6426 = key[103:96] ;
assign n6427 =  ( n6425 ) ^ ( n6426 )  ;
assign n6428 =  { ( n6421 ) , ( n6427 ) }  ;
assign n6429 = state_in[103:96] ;
assign n6430 =  ( n6429 ) == ( bv_8_255_n3 )  ;
assign n6431 = state_in[103:96] ;
assign n6432 =  ( n6431 ) == ( bv_8_254_n7 )  ;
assign n6433 = state_in[103:96] ;
assign n6434 =  ( n6433 ) == ( bv_8_253_n11 )  ;
assign n6435 = state_in[103:96] ;
assign n6436 =  ( n6435 ) == ( bv_8_252_n15 )  ;
assign n6437 = state_in[103:96] ;
assign n6438 =  ( n6437 ) == ( bv_8_251_n19 )  ;
assign n6439 = state_in[103:96] ;
assign n6440 =  ( n6439 ) == ( bv_8_250_n23 )  ;
assign n6441 = state_in[103:96] ;
assign n6442 =  ( n6441 ) == ( bv_8_249_n27 )  ;
assign n6443 = state_in[103:96] ;
assign n6444 =  ( n6443 ) == ( bv_8_248_n31 )  ;
assign n6445 = state_in[103:96] ;
assign n6446 =  ( n6445 ) == ( bv_8_247_n35 )  ;
assign n6447 = state_in[103:96] ;
assign n6448 =  ( n6447 ) == ( bv_8_246_n39 )  ;
assign n6449 = state_in[103:96] ;
assign n6450 =  ( n6449 ) == ( bv_8_245_n43 )  ;
assign n6451 = state_in[103:96] ;
assign n6452 =  ( n6451 ) == ( bv_8_244_n47 )  ;
assign n6453 = state_in[103:96] ;
assign n6454 =  ( n6453 ) == ( bv_8_243_n51 )  ;
assign n6455 = state_in[103:96] ;
assign n6456 =  ( n6455 ) == ( bv_8_242_n55 )  ;
assign n6457 = state_in[103:96] ;
assign n6458 =  ( n6457 ) == ( bv_8_241_n59 )  ;
assign n6459 = state_in[103:96] ;
assign n6460 =  ( n6459 ) == ( bv_8_240_n63 )  ;
assign n6461 = state_in[103:96] ;
assign n6462 =  ( n6461 ) == ( bv_8_239_n67 )  ;
assign n6463 = state_in[103:96] ;
assign n6464 =  ( n6463 ) == ( bv_8_238_n71 )  ;
assign n6465 = state_in[103:96] ;
assign n6466 =  ( n6465 ) == ( bv_8_237_n75 )  ;
assign n6467 = state_in[103:96] ;
assign n6468 =  ( n6467 ) == ( bv_8_236_n79 )  ;
assign n6469 = state_in[103:96] ;
assign n6470 =  ( n6469 ) == ( bv_8_235_n83 )  ;
assign n6471 = state_in[103:96] ;
assign n6472 =  ( n6471 ) == ( bv_8_234_n87 )  ;
assign n6473 = state_in[103:96] ;
assign n6474 =  ( n6473 ) == ( bv_8_233_n91 )  ;
assign n6475 = state_in[103:96] ;
assign n6476 =  ( n6475 ) == ( bv_8_232_n95 )  ;
assign n6477 = state_in[103:96] ;
assign n6478 =  ( n6477 ) == ( bv_8_231_n99 )  ;
assign n6479 = state_in[103:96] ;
assign n6480 =  ( n6479 ) == ( bv_8_230_n103 )  ;
assign n6481 = state_in[103:96] ;
assign n6482 =  ( n6481 ) == ( bv_8_229_n107 )  ;
assign n6483 = state_in[103:96] ;
assign n6484 =  ( n6483 ) == ( bv_8_228_n111 )  ;
assign n6485 = state_in[103:96] ;
assign n6486 =  ( n6485 ) == ( bv_8_227_n115 )  ;
assign n6487 = state_in[103:96] ;
assign n6488 =  ( n6487 ) == ( bv_8_226_n119 )  ;
assign n6489 = state_in[103:96] ;
assign n6490 =  ( n6489 ) == ( bv_8_225_n123 )  ;
assign n6491 = state_in[103:96] ;
assign n6492 =  ( n6491 ) == ( bv_8_224_n126 )  ;
assign n6493 = state_in[103:96] ;
assign n6494 =  ( n6493 ) == ( bv_8_223_n130 )  ;
assign n6495 = state_in[103:96] ;
assign n6496 =  ( n6495 ) == ( bv_8_222_n134 )  ;
assign n6497 = state_in[103:96] ;
assign n6498 =  ( n6497 ) == ( bv_8_221_n138 )  ;
assign n6499 = state_in[103:96] ;
assign n6500 =  ( n6499 ) == ( bv_8_220_n142 )  ;
assign n6501 = state_in[103:96] ;
assign n6502 =  ( n6501 ) == ( bv_8_219_n146 )  ;
assign n6503 = state_in[103:96] ;
assign n6504 =  ( n6503 ) == ( bv_8_218_n150 )  ;
assign n6505 = state_in[103:96] ;
assign n6506 =  ( n6505 ) == ( bv_8_217_n128 )  ;
assign n6507 = state_in[103:96] ;
assign n6508 =  ( n6507 ) == ( bv_8_216_n157 )  ;
assign n6509 = state_in[103:96] ;
assign n6510 =  ( n6509 ) == ( bv_8_215_n45 )  ;
assign n6511 = state_in[103:96] ;
assign n6512 =  ( n6511 ) == ( bv_8_214_n164 )  ;
assign n6513 = state_in[103:96] ;
assign n6514 =  ( n6513 ) == ( bv_8_213_n167 )  ;
assign n6515 = state_in[103:96] ;
assign n6516 =  ( n6515 ) == ( bv_8_212_n171 )  ;
assign n6517 = state_in[103:96] ;
assign n6518 =  ( n6517 ) == ( bv_8_211_n175 )  ;
assign n6519 = state_in[103:96] ;
assign n6520 =  ( n6519 ) == ( bv_8_210_n113 )  ;
assign n6521 = state_in[103:96] ;
assign n6522 =  ( n6521 ) == ( bv_8_209_n182 )  ;
assign n6523 = state_in[103:96] ;
assign n6524 =  ( n6523 ) == ( bv_8_208_n37 )  ;
assign n6525 = state_in[103:96] ;
assign n6526 =  ( n6525 ) == ( bv_8_207_n188 )  ;
assign n6527 = state_in[103:96] ;
assign n6528 =  ( n6527 ) == ( bv_8_206_n192 )  ;
assign n6529 = state_in[103:96] ;
assign n6530 =  ( n6529 ) == ( bv_8_205_n196 )  ;
assign n6531 = state_in[103:96] ;
assign n6532 =  ( n6531 ) == ( bv_8_204_n177 )  ;
assign n6533 = state_in[103:96] ;
assign n6534 =  ( n6533 ) == ( bv_8_203_n203 )  ;
assign n6535 = state_in[103:96] ;
assign n6536 =  ( n6535 ) == ( bv_8_202_n207 )  ;
assign n6537 = state_in[103:96] ;
assign n6538 =  ( n6537 ) == ( bv_8_201_n85 )  ;
assign n6539 = state_in[103:96] ;
assign n6540 =  ( n6539 ) == ( bv_8_200_n213 )  ;
assign n6541 = state_in[103:96] ;
assign n6542 =  ( n6541 ) == ( bv_8_199_n216 )  ;
assign n6543 = state_in[103:96] ;
assign n6544 =  ( n6543 ) == ( bv_8_198_n220 )  ;
assign n6545 = state_in[103:96] ;
assign n6546 =  ( n6545 ) == ( bv_8_197_n224 )  ;
assign n6547 = state_in[103:96] ;
assign n6548 =  ( n6547 ) == ( bv_8_196_n228 )  ;
assign n6549 = state_in[103:96] ;
assign n6550 =  ( n6549 ) == ( bv_8_195_n232 )  ;
assign n6551 = state_in[103:96] ;
assign n6552 =  ( n6551 ) == ( bv_8_194_n159 )  ;
assign n6553 = state_in[103:96] ;
assign n6554 =  ( n6553 ) == ( bv_8_193_n239 )  ;
assign n6555 = state_in[103:96] ;
assign n6556 =  ( n6555 ) == ( bv_8_192_n242 )  ;
assign n6557 = state_in[103:96] ;
assign n6558 =  ( n6557 ) == ( bv_8_191_n246 )  ;
assign n6559 = state_in[103:96] ;
assign n6560 =  ( n6559 ) == ( bv_8_190_n250 )  ;
assign n6561 = state_in[103:96] ;
assign n6562 =  ( n6561 ) == ( bv_8_189_n254 )  ;
assign n6563 = state_in[103:96] ;
assign n6564 =  ( n6563 ) == ( bv_8_188_n257 )  ;
assign n6565 = state_in[103:96] ;
assign n6566 =  ( n6565 ) == ( bv_8_187_n260 )  ;
assign n6567 = state_in[103:96] ;
assign n6568 =  ( n6567 ) == ( bv_8_186_n263 )  ;
assign n6569 = state_in[103:96] ;
assign n6570 =  ( n6569 ) == ( bv_8_185_n266 )  ;
assign n6571 = state_in[103:96] ;
assign n6572 =  ( n6571 ) == ( bv_8_184_n270 )  ;
assign n6573 = state_in[103:96] ;
assign n6574 =  ( n6573 ) == ( bv_8_183_n273 )  ;
assign n6575 = state_in[103:96] ;
assign n6576 =  ( n6575 ) == ( bv_8_182_n277 )  ;
assign n6577 = state_in[103:96] ;
assign n6578 =  ( n6577 ) == ( bv_8_181_n281 )  ;
assign n6579 = state_in[103:96] ;
assign n6580 =  ( n6579 ) == ( bv_8_180_n285 )  ;
assign n6581 = state_in[103:96] ;
assign n6582 =  ( n6581 ) == ( bv_8_179_n289 )  ;
assign n6583 = state_in[103:96] ;
assign n6584 =  ( n6583 ) == ( bv_8_178_n292 )  ;
assign n6585 = state_in[103:96] ;
assign n6586 =  ( n6585 ) == ( bv_8_177_n283 )  ;
assign n6587 = state_in[103:96] ;
assign n6588 =  ( n6587 ) == ( bv_8_176_n299 )  ;
assign n6589 = state_in[103:96] ;
assign n6590 =  ( n6589 ) == ( bv_8_175_n302 )  ;
assign n6591 = state_in[103:96] ;
assign n6592 =  ( n6591 ) == ( bv_8_174_n152 )  ;
assign n6593 = state_in[103:96] ;
assign n6594 =  ( n6593 ) == ( bv_8_173_n307 )  ;
assign n6595 = state_in[103:96] ;
assign n6596 =  ( n6595 ) == ( bv_8_172_n268 )  ;
assign n6597 = state_in[103:96] ;
assign n6598 =  ( n6597 ) == ( bv_8_171_n314 )  ;
assign n6599 = state_in[103:96] ;
assign n6600 =  ( n6599 ) == ( bv_8_170_n77 )  ;
assign n6601 = state_in[103:96] ;
assign n6602 =  ( n6601 ) == ( bv_8_169_n109 )  ;
assign n6603 = state_in[103:96] ;
assign n6604 =  ( n6603 ) == ( bv_8_168_n13 )  ;
assign n6605 = state_in[103:96] ;
assign n6606 =  ( n6605 ) == ( bv_8_167_n325 )  ;
assign n6607 = state_in[103:96] ;
assign n6608 =  ( n6607 ) == ( bv_8_166_n328 )  ;
assign n6609 = state_in[103:96] ;
assign n6610 =  ( n6609 ) == ( bv_8_165_n69 )  ;
assign n6611 = state_in[103:96] ;
assign n6612 =  ( n6611 ) == ( bv_8_164_n335 )  ;
assign n6613 = state_in[103:96] ;
assign n6614 =  ( n6613 ) == ( bv_8_163_n339 )  ;
assign n6615 = state_in[103:96] ;
assign n6616 =  ( n6615 ) == ( bv_8_162_n343 )  ;
assign n6617 = state_in[103:96] ;
assign n6618 =  ( n6617 ) == ( bv_8_161_n211 )  ;
assign n6619 = state_in[103:96] ;
assign n6620 =  ( n6619 ) == ( bv_8_160_n350 )  ;
assign n6621 = state_in[103:96] ;
assign n6622 =  ( n6621 ) == ( bv_8_159_n323 )  ;
assign n6623 = state_in[103:96] ;
assign n6624 =  ( n6623 ) == ( bv_8_158_n355 )  ;
assign n6625 = state_in[103:96] ;
assign n6626 =  ( n6625 ) == ( bv_8_157_n359 )  ;
assign n6627 = state_in[103:96] ;
assign n6628 =  ( n6627 ) == ( bv_8_156_n279 )  ;
assign n6629 = state_in[103:96] ;
assign n6630 =  ( n6629 ) == ( bv_8_155_n364 )  ;
assign n6631 = state_in[103:96] ;
assign n6632 =  ( n6631 ) == ( bv_8_154_n368 )  ;
assign n6633 = state_in[103:96] ;
assign n6634 =  ( n6633 ) == ( bv_8_153_n140 )  ;
assign n6635 = state_in[103:96] ;
assign n6636 =  ( n6635 ) == ( bv_8_152_n374 )  ;
assign n6637 = state_in[103:96] ;
assign n6638 =  ( n6637 ) == ( bv_8_151_n218 )  ;
assign n6639 = state_in[103:96] ;
assign n6640 =  ( n6639 ) == ( bv_8_150_n201 )  ;
assign n6641 = state_in[103:96] ;
assign n6642 =  ( n6641 ) == ( bv_8_149_n384 )  ;
assign n6643 = state_in[103:96] ;
assign n6644 =  ( n6643 ) == ( bv_8_148_n388 )  ;
assign n6645 = state_in[103:96] ;
assign n6646 =  ( n6645 ) == ( bv_8_147_n392 )  ;
assign n6647 = state_in[103:96] ;
assign n6648 =  ( n6647 ) == ( bv_8_146_n337 )  ;
assign n6649 = state_in[103:96] ;
assign n6650 =  ( n6649 ) == ( bv_8_145_n397 )  ;
assign n6651 = state_in[103:96] ;
assign n6652 =  ( n6651 ) == ( bv_8_144_n173 )  ;
assign n6653 = state_in[103:96] ;
assign n6654 =  ( n6653 ) == ( bv_8_143_n403 )  ;
assign n6655 = state_in[103:96] ;
assign n6656 =  ( n6655 ) == ( bv_8_142_n406 )  ;
assign n6657 = state_in[103:96] ;
assign n6658 =  ( n6657 ) == ( bv_8_141_n410 )  ;
assign n6659 = state_in[103:96] ;
assign n6660 =  ( n6659 ) == ( bv_8_140_n376 )  ;
assign n6661 = state_in[103:96] ;
assign n6662 =  ( n6661 ) == ( bv_8_139_n297 )  ;
assign n6663 = state_in[103:96] ;
assign n6664 =  ( n6663 ) == ( bv_8_138_n418 )  ;
assign n6665 = state_in[103:96] ;
assign n6666 =  ( n6665 ) == ( bv_8_137_n421 )  ;
assign n6667 = state_in[103:96] ;
assign n6668 =  ( n6667 ) == ( bv_8_136_n425 )  ;
assign n6669 = state_in[103:96] ;
assign n6670 =  ( n6669 ) == ( bv_8_135_n81 )  ;
assign n6671 = state_in[103:96] ;
assign n6672 =  ( n6671 ) == ( bv_8_134_n431 )  ;
assign n6673 = state_in[103:96] ;
assign n6674 =  ( n6673 ) == ( bv_8_133_n434 )  ;
assign n6675 = state_in[103:96] ;
assign n6676 =  ( n6675 ) == ( bv_8_132_n41 )  ;
assign n6677 = state_in[103:96] ;
assign n6678 =  ( n6677 ) == ( bv_8_131_n440 )  ;
assign n6679 = state_in[103:96] ;
assign n6680 =  ( n6679 ) == ( bv_8_130_n33 )  ;
assign n6681 = state_in[103:96] ;
assign n6682 =  ( n6681 ) == ( bv_8_129_n446 )  ;
assign n6683 = state_in[103:96] ;
assign n6684 =  ( n6683 ) == ( bv_8_128_n450 )  ;
assign n6685 = state_in[103:96] ;
assign n6686 =  ( n6685 ) == ( bv_8_127_n453 )  ;
assign n6687 = state_in[103:96] ;
assign n6688 =  ( n6687 ) == ( bv_8_126_n456 )  ;
assign n6689 = state_in[103:96] ;
assign n6690 =  ( n6689 ) == ( bv_8_125_n459 )  ;
assign n6691 = state_in[103:96] ;
assign n6692 =  ( n6691 ) == ( bv_8_124_n184 )  ;
assign n6693 = state_in[103:96] ;
assign n6694 =  ( n6693 ) == ( bv_8_123_n17 )  ;
assign n6695 = state_in[103:96] ;
assign n6696 =  ( n6695 ) == ( bv_8_122_n416 )  ;
assign n6697 = state_in[103:96] ;
assign n6698 =  ( n6697 ) == ( bv_8_121_n470 )  ;
assign n6699 = state_in[103:96] ;
assign n6700 =  ( n6699 ) == ( bv_8_120_n474 )  ;
assign n6701 = state_in[103:96] ;
assign n6702 =  ( n6701 ) == ( bv_8_119_n472 )  ;
assign n6703 = state_in[103:96] ;
assign n6704 =  ( n6703 ) == ( bv_8_118_n480 )  ;
assign n6705 = state_in[103:96] ;
assign n6706 =  ( n6705 ) == ( bv_8_117_n484 )  ;
assign n6707 = state_in[103:96] ;
assign n6708 =  ( n6707 ) == ( bv_8_116_n345 )  ;
assign n6709 = state_in[103:96] ;
assign n6710 =  ( n6709 ) == ( bv_8_115_n222 )  ;
assign n6711 = state_in[103:96] ;
assign n6712 =  ( n6711 ) == ( bv_8_114_n494 )  ;
assign n6713 = state_in[103:96] ;
assign n6714 =  ( n6713 ) == ( bv_8_113_n180 )  ;
assign n6715 = state_in[103:96] ;
assign n6716 =  ( n6715 ) == ( bv_8_112_n482 )  ;
assign n6717 = state_in[103:96] ;
assign n6718 =  ( n6717 ) == ( bv_8_111_n244 )  ;
assign n6719 = state_in[103:96] ;
assign n6720 =  ( n6719 ) == ( bv_8_110_n294 )  ;
assign n6721 = state_in[103:96] ;
assign n6722 =  ( n6721 ) == ( bv_8_109_n9 )  ;
assign n6723 = state_in[103:96] ;
assign n6724 =  ( n6723 ) == ( bv_8_108_n510 )  ;
assign n6725 = state_in[103:96] ;
assign n6726 =  ( n6725 ) == ( bv_8_107_n370 )  ;
assign n6727 = state_in[103:96] ;
assign n6728 =  ( n6727 ) == ( bv_8_106_n155 )  ;
assign n6729 = state_in[103:96] ;
assign n6730 =  ( n6729 ) == ( bv_8_105_n148 )  ;
assign n6731 = state_in[103:96] ;
assign n6732 =  ( n6731 ) == ( bv_8_104_n520 )  ;
assign n6733 = state_in[103:96] ;
assign n6734 =  ( n6733 ) == ( bv_8_103_n523 )  ;
assign n6735 = state_in[103:96] ;
assign n6736 =  ( n6735 ) == ( bv_8_102_n527 )  ;
assign n6737 = state_in[103:96] ;
assign n6738 =  ( n6737 ) == ( bv_8_101_n49 )  ;
assign n6739 = state_in[103:96] ;
assign n6740 =  ( n6739 ) == ( bv_8_100_n348 )  ;
assign n6741 = state_in[103:96] ;
assign n6742 =  ( n6741 ) == ( bv_8_99_n476 )  ;
assign n6743 = state_in[103:96] ;
assign n6744 =  ( n6743 ) == ( bv_8_98_n536 )  ;
assign n6745 = state_in[103:96] ;
assign n6746 =  ( n6745 ) == ( bv_8_97_n198 )  ;
assign n6747 = state_in[103:96] ;
assign n6748 =  ( n6747 ) == ( bv_8_96_n542 )  ;
assign n6749 = state_in[103:96] ;
assign n6750 =  ( n6749 ) == ( bv_8_95_n545 )  ;
assign n6751 = state_in[103:96] ;
assign n6752 =  ( n6751 ) == ( bv_8_94_n548 )  ;
assign n6753 = state_in[103:96] ;
assign n6754 =  ( n6753 ) == ( bv_8_93_n498 )  ;
assign n6755 = state_in[103:96] ;
assign n6756 =  ( n6755 ) == ( bv_8_92_n234 )  ;
assign n6757 = state_in[103:96] ;
assign n6758 =  ( n6757 ) == ( bv_8_91_n555 )  ;
assign n6759 = state_in[103:96] ;
assign n6760 =  ( n6759 ) == ( bv_8_90_n25 )  ;
assign n6761 = state_in[103:96] ;
assign n6762 =  ( n6761 ) == ( bv_8_89_n61 )  ;
assign n6763 = state_in[103:96] ;
assign n6764 =  ( n6763 ) == ( bv_8_88_n562 )  ;
assign n6765 = state_in[103:96] ;
assign n6766 =  ( n6765 ) == ( bv_8_87_n226 )  ;
assign n6767 = state_in[103:96] ;
assign n6768 =  ( n6767 ) == ( bv_8_86_n567 )  ;
assign n6769 = state_in[103:96] ;
assign n6770 =  ( n6769 ) == ( bv_8_85_n423 )  ;
assign n6771 = state_in[103:96] ;
assign n6772 =  ( n6771 ) == ( bv_8_84_n386 )  ;
assign n6773 = state_in[103:96] ;
assign n6774 =  ( n6773 ) == ( bv_8_83_n575 )  ;
assign n6775 = state_in[103:96] ;
assign n6776 =  ( n6775 ) == ( bv_8_82_n578 )  ;
assign n6777 = state_in[103:96] ;
assign n6778 =  ( n6777 ) == ( bv_8_81_n582 )  ;
assign n6779 = state_in[103:96] ;
assign n6780 =  ( n6779 ) == ( bv_8_80_n73 )  ;
assign n6781 = state_in[103:96] ;
assign n6782 =  ( n6781 ) == ( bv_8_79_n538 )  ;
assign n6783 = state_in[103:96] ;
assign n6784 =  ( n6783 ) == ( bv_8_78_n590 )  ;
assign n6785 = state_in[103:96] ;
assign n6786 =  ( n6785 ) == ( bv_8_77_n593 )  ;
assign n6787 = state_in[103:96] ;
assign n6788 =  ( n6787 ) == ( bv_8_76_n596 )  ;
assign n6789 = state_in[103:96] ;
assign n6790 =  ( n6789 ) == ( bv_8_75_n503 )  ;
assign n6791 = state_in[103:96] ;
assign n6792 =  ( n6791 ) == ( bv_8_74_n237 )  ;
assign n6793 = state_in[103:96] ;
assign n6794 =  ( n6793 ) == ( bv_8_73_n275 )  ;
assign n6795 = state_in[103:96] ;
assign n6796 =  ( n6795 ) == ( bv_8_72_n330 )  ;
assign n6797 = state_in[103:96] ;
assign n6798 =  ( n6797 ) == ( bv_8_71_n252 )  ;
assign n6799 = state_in[103:96] ;
assign n6800 =  ( n6799 ) == ( bv_8_70_n609 )  ;
assign n6801 = state_in[103:96] ;
assign n6802 =  ( n6801 ) == ( bv_8_69_n612 )  ;
assign n6803 = state_in[103:96] ;
assign n6804 =  ( n6803 ) == ( bv_8_68_n390 )  ;
assign n6805 = state_in[103:96] ;
assign n6806 =  ( n6805 ) == ( bv_8_67_n318 )  ;
assign n6807 = state_in[103:96] ;
assign n6808 =  ( n6807 ) == ( bv_8_66_n466 )  ;
assign n6809 = state_in[103:96] ;
assign n6810 =  ( n6809 ) == ( bv_8_65_n623 )  ;
assign n6811 = state_in[103:96] ;
assign n6812 =  ( n6811 ) == ( bv_8_64_n573 )  ;
assign n6813 = state_in[103:96] ;
assign n6814 =  ( n6813 ) == ( bv_8_63_n489 )  ;
assign n6815 = state_in[103:96] ;
assign n6816 =  ( n6815 ) == ( bv_8_62_n205 )  ;
assign n6817 = state_in[103:96] ;
assign n6818 =  ( n6817 ) == ( bv_8_61_n634 )  ;
assign n6819 = state_in[103:96] ;
assign n6820 =  ( n6819 ) == ( bv_8_60_n93 )  ;
assign n6821 = state_in[103:96] ;
assign n6822 =  ( n6821 ) == ( bv_8_59_n382 )  ;
assign n6823 = state_in[103:96] ;
assign n6824 =  ( n6823 ) == ( bv_8_58_n136 )  ;
assign n6825 = state_in[103:96] ;
assign n6826 =  ( n6825 ) == ( bv_8_57_n312 )  ;
assign n6827 = state_in[103:96] ;
assign n6828 =  ( n6827 ) == ( bv_8_56_n230 )  ;
assign n6829 = state_in[103:96] ;
assign n6830 =  ( n6829 ) == ( bv_8_55_n650 )  ;
assign n6831 = state_in[103:96] ;
assign n6832 =  ( n6831 ) == ( bv_8_54_n616 )  ;
assign n6833 = state_in[103:96] ;
assign n6834 =  ( n6833 ) == ( bv_8_53_n436 )  ;
assign n6835 = state_in[103:96] ;
assign n6836 =  ( n6835 ) == ( bv_8_52_n619 )  ;
assign n6837 = state_in[103:96] ;
assign n6838 =  ( n6837 ) == ( bv_8_51_n101 )  ;
assign n6839 = state_in[103:96] ;
assign n6840 =  ( n6839 ) == ( bv_8_50_n408 )  ;
assign n6841 = state_in[103:96] ;
assign n6842 =  ( n6841 ) == ( bv_8_49_n309 )  ;
assign n6843 = state_in[103:96] ;
assign n6844 =  ( n6843 ) == ( bv_8_48_n660 )  ;
assign n6845 = state_in[103:96] ;
assign n6846 =  ( n6845 ) == ( bv_8_47_n652 )  ;
assign n6847 = state_in[103:96] ;
assign n6848 =  ( n6847 ) == ( bv_8_46_n429 )  ;
assign n6849 = state_in[103:96] ;
assign n6850 =  ( n6849 ) == ( bv_8_45_n97 )  ;
assign n6851 = state_in[103:96] ;
assign n6852 =  ( n6851 ) == ( bv_8_44_n5 )  ;
assign n6853 = state_in[103:96] ;
assign n6854 =  ( n6853 ) == ( bv_8_43_n121 )  ;
assign n6855 = state_in[103:96] ;
assign n6856 =  ( n6855 ) == ( bv_8_42_n672 )  ;
assign n6857 = state_in[103:96] ;
assign n6858 =  ( n6857 ) == ( bv_8_41_n29 )  ;
assign n6859 = state_in[103:96] ;
assign n6860 =  ( n6859 ) == ( bv_8_40_n366 )  ;
assign n6861 = state_in[103:96] ;
assign n6862 =  ( n6861 ) == ( bv_8_39_n132 )  ;
assign n6863 = state_in[103:96] ;
assign n6864 =  ( n6863 ) == ( bv_8_38_n444 )  ;
assign n6865 = state_in[103:96] ;
assign n6866 =  ( n6865 ) == ( bv_8_37_n506 )  ;
assign n6867 = state_in[103:96] ;
assign n6868 =  ( n6867 ) == ( bv_8_36_n645 )  ;
assign n6869 = state_in[103:96] ;
assign n6870 =  ( n6869 ) == ( bv_8_35_n696 )  ;
assign n6871 = state_in[103:96] ;
assign n6872 =  ( n6871 ) == ( bv_8_34_n117 )  ;
assign n6873 = state_in[103:96] ;
assign n6874 =  ( n6873 ) == ( bv_8_33_n486 )  ;
assign n6875 = state_in[103:96] ;
assign n6876 =  ( n6875 ) == ( bv_8_32_n463 )  ;
assign n6877 = state_in[103:96] ;
assign n6878 =  ( n6877 ) == ( bv_8_31_n705 )  ;
assign n6879 = state_in[103:96] ;
assign n6880 =  ( n6879 ) == ( bv_8_30_n21 )  ;
assign n6881 = state_in[103:96] ;
assign n6882 =  ( n6881 ) == ( bv_8_29_n625 )  ;
assign n6883 = state_in[103:96] ;
assign n6884 =  ( n6883 ) == ( bv_8_28_n162 )  ;
assign n6885 = state_in[103:96] ;
assign n6886 =  ( n6885 ) == ( bv_8_27_n642 )  ;
assign n6887 = state_in[103:96] ;
assign n6888 =  ( n6887 ) == ( bv_8_26_n53 )  ;
assign n6889 = state_in[103:96] ;
assign n6890 =  ( n6889 ) == ( bv_8_25_n399 )  ;
assign n6891 = state_in[103:96] ;
assign n6892 =  ( n6891 ) == ( bv_8_24_n448 )  ;
assign n6893 = state_in[103:96] ;
assign n6894 =  ( n6893 ) == ( bv_8_23_n144 )  ;
assign n6895 = state_in[103:96] ;
assign n6896 =  ( n6895 ) == ( bv_8_22_n357 )  ;
assign n6897 = state_in[103:96] ;
assign n6898 =  ( n6897 ) == ( bv_8_21_n89 )  ;
assign n6899 = state_in[103:96] ;
assign n6900 =  ( n6899 ) == ( bv_8_20_n341 )  ;
assign n6901 = state_in[103:96] ;
assign n6902 =  ( n6901 ) == ( bv_8_19_n588 )  ;
assign n6903 = state_in[103:96] ;
assign n6904 =  ( n6903 ) == ( bv_8_18_n628 )  ;
assign n6905 = state_in[103:96] ;
assign n6906 =  ( n6905 ) == ( bv_8_17_n525 )  ;
assign n6907 = state_in[103:96] ;
assign n6908 =  ( n6907 ) == ( bv_8_16_n248 )  ;
assign n6909 = state_in[103:96] ;
assign n6910 =  ( n6909 ) == ( bv_8_15_n190 )  ;
assign n6911 = state_in[103:96] ;
assign n6912 =  ( n6911 ) == ( bv_8_14_n648 )  ;
assign n6913 = state_in[103:96] ;
assign n6914 =  ( n6913 ) == ( bv_8_13_n194 )  ;
assign n6915 = state_in[103:96] ;
assign n6916 =  ( n6915 ) == ( bv_8_12_n333 )  ;
assign n6917 = state_in[103:96] ;
assign n6918 =  ( n6917 ) == ( bv_8_11_n379 )  ;
assign n6919 = state_in[103:96] ;
assign n6920 =  ( n6919 ) == ( bv_8_10_n655 )  ;
assign n6921 = state_in[103:96] ;
assign n6922 =  ( n6921 ) == ( bv_8_9_n57 )  ;
assign n6923 = state_in[103:96] ;
assign n6924 =  ( n6923 ) == ( bv_8_8_n669 )  ;
assign n6925 = state_in[103:96] ;
assign n6926 =  ( n6925 ) == ( bv_8_7_n105 )  ;
assign n6927 = state_in[103:96] ;
assign n6928 =  ( n6927 ) == ( bv_8_6_n169 )  ;
assign n6929 = state_in[103:96] ;
assign n6930 =  ( n6929 ) == ( bv_8_5_n492 )  ;
assign n6931 = state_in[103:96] ;
assign n6932 =  ( n6931 ) == ( bv_8_4_n516 )  ;
assign n6933 = state_in[103:96] ;
assign n6934 =  ( n6933 ) == ( bv_8_3_n65 )  ;
assign n6935 = state_in[103:96] ;
assign n6936 =  ( n6935 ) == ( bv_8_2_n751 )  ;
assign n6937 = state_in[103:96] ;
assign n6938 =  ( n6937 ) == ( bv_8_1_n287 )  ;
assign n6939 = state_in[103:96] ;
assign n6940 =  ( n6939 ) == ( bv_8_0_n580 )  ;
assign n6941 =  ( n6940 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n6942 =  ( n6938 ) ? ( bv_8_124_n184 ) : ( n6941 ) ;
assign n6943 =  ( n6936 ) ? ( bv_8_119_n472 ) : ( n6942 ) ;
assign n6944 =  ( n6934 ) ? ( bv_8_123_n17 ) : ( n6943 ) ;
assign n6945 =  ( n6932 ) ? ( bv_8_242_n55 ) : ( n6944 ) ;
assign n6946 =  ( n6930 ) ? ( bv_8_107_n370 ) : ( n6945 ) ;
assign n6947 =  ( n6928 ) ? ( bv_8_111_n244 ) : ( n6946 ) ;
assign n6948 =  ( n6926 ) ? ( bv_8_197_n224 ) : ( n6947 ) ;
assign n6949 =  ( n6924 ) ? ( bv_8_48_n660 ) : ( n6948 ) ;
assign n6950 =  ( n6922 ) ? ( bv_8_1_n287 ) : ( n6949 ) ;
assign n6951 =  ( n6920 ) ? ( bv_8_103_n523 ) : ( n6950 ) ;
assign n6952 =  ( n6918 ) ? ( bv_8_43_n121 ) : ( n6951 ) ;
assign n6953 =  ( n6916 ) ? ( bv_8_254_n7 ) : ( n6952 ) ;
assign n6954 =  ( n6914 ) ? ( bv_8_215_n45 ) : ( n6953 ) ;
assign n6955 =  ( n6912 ) ? ( bv_8_171_n314 ) : ( n6954 ) ;
assign n6956 =  ( n6910 ) ? ( bv_8_118_n480 ) : ( n6955 ) ;
assign n6957 =  ( n6908 ) ? ( bv_8_202_n207 ) : ( n6956 ) ;
assign n6958 =  ( n6906 ) ? ( bv_8_130_n33 ) : ( n6957 ) ;
assign n6959 =  ( n6904 ) ? ( bv_8_201_n85 ) : ( n6958 ) ;
assign n6960 =  ( n6902 ) ? ( bv_8_125_n459 ) : ( n6959 ) ;
assign n6961 =  ( n6900 ) ? ( bv_8_250_n23 ) : ( n6960 ) ;
assign n6962 =  ( n6898 ) ? ( bv_8_89_n61 ) : ( n6961 ) ;
assign n6963 =  ( n6896 ) ? ( bv_8_71_n252 ) : ( n6962 ) ;
assign n6964 =  ( n6894 ) ? ( bv_8_240_n63 ) : ( n6963 ) ;
assign n6965 =  ( n6892 ) ? ( bv_8_173_n307 ) : ( n6964 ) ;
assign n6966 =  ( n6890 ) ? ( bv_8_212_n171 ) : ( n6965 ) ;
assign n6967 =  ( n6888 ) ? ( bv_8_162_n343 ) : ( n6966 ) ;
assign n6968 =  ( n6886 ) ? ( bv_8_175_n302 ) : ( n6967 ) ;
assign n6969 =  ( n6884 ) ? ( bv_8_156_n279 ) : ( n6968 ) ;
assign n6970 =  ( n6882 ) ? ( bv_8_164_n335 ) : ( n6969 ) ;
assign n6971 =  ( n6880 ) ? ( bv_8_114_n494 ) : ( n6970 ) ;
assign n6972 =  ( n6878 ) ? ( bv_8_192_n242 ) : ( n6971 ) ;
assign n6973 =  ( n6876 ) ? ( bv_8_183_n273 ) : ( n6972 ) ;
assign n6974 =  ( n6874 ) ? ( bv_8_253_n11 ) : ( n6973 ) ;
assign n6975 =  ( n6872 ) ? ( bv_8_147_n392 ) : ( n6974 ) ;
assign n6976 =  ( n6870 ) ? ( bv_8_38_n444 ) : ( n6975 ) ;
assign n6977 =  ( n6868 ) ? ( bv_8_54_n616 ) : ( n6976 ) ;
assign n6978 =  ( n6866 ) ? ( bv_8_63_n489 ) : ( n6977 ) ;
assign n6979 =  ( n6864 ) ? ( bv_8_247_n35 ) : ( n6978 ) ;
assign n6980 =  ( n6862 ) ? ( bv_8_204_n177 ) : ( n6979 ) ;
assign n6981 =  ( n6860 ) ? ( bv_8_52_n619 ) : ( n6980 ) ;
assign n6982 =  ( n6858 ) ? ( bv_8_165_n69 ) : ( n6981 ) ;
assign n6983 =  ( n6856 ) ? ( bv_8_229_n107 ) : ( n6982 ) ;
assign n6984 =  ( n6854 ) ? ( bv_8_241_n59 ) : ( n6983 ) ;
assign n6985 =  ( n6852 ) ? ( bv_8_113_n180 ) : ( n6984 ) ;
assign n6986 =  ( n6850 ) ? ( bv_8_216_n157 ) : ( n6985 ) ;
assign n6987 =  ( n6848 ) ? ( bv_8_49_n309 ) : ( n6986 ) ;
assign n6988 =  ( n6846 ) ? ( bv_8_21_n89 ) : ( n6987 ) ;
assign n6989 =  ( n6844 ) ? ( bv_8_4_n516 ) : ( n6988 ) ;
assign n6990 =  ( n6842 ) ? ( bv_8_199_n216 ) : ( n6989 ) ;
assign n6991 =  ( n6840 ) ? ( bv_8_35_n696 ) : ( n6990 ) ;
assign n6992 =  ( n6838 ) ? ( bv_8_195_n232 ) : ( n6991 ) ;
assign n6993 =  ( n6836 ) ? ( bv_8_24_n448 ) : ( n6992 ) ;
assign n6994 =  ( n6834 ) ? ( bv_8_150_n201 ) : ( n6993 ) ;
assign n6995 =  ( n6832 ) ? ( bv_8_5_n492 ) : ( n6994 ) ;
assign n6996 =  ( n6830 ) ? ( bv_8_154_n368 ) : ( n6995 ) ;
assign n6997 =  ( n6828 ) ? ( bv_8_7_n105 ) : ( n6996 ) ;
assign n6998 =  ( n6826 ) ? ( bv_8_18_n628 ) : ( n6997 ) ;
assign n6999 =  ( n6824 ) ? ( bv_8_128_n450 ) : ( n6998 ) ;
assign n7000 =  ( n6822 ) ? ( bv_8_226_n119 ) : ( n6999 ) ;
assign n7001 =  ( n6820 ) ? ( bv_8_235_n83 ) : ( n7000 ) ;
assign n7002 =  ( n6818 ) ? ( bv_8_39_n132 ) : ( n7001 ) ;
assign n7003 =  ( n6816 ) ? ( bv_8_178_n292 ) : ( n7002 ) ;
assign n7004 =  ( n6814 ) ? ( bv_8_117_n484 ) : ( n7003 ) ;
assign n7005 =  ( n6812 ) ? ( bv_8_9_n57 ) : ( n7004 ) ;
assign n7006 =  ( n6810 ) ? ( bv_8_131_n440 ) : ( n7005 ) ;
assign n7007 =  ( n6808 ) ? ( bv_8_44_n5 ) : ( n7006 ) ;
assign n7008 =  ( n6806 ) ? ( bv_8_26_n53 ) : ( n7007 ) ;
assign n7009 =  ( n6804 ) ? ( bv_8_27_n642 ) : ( n7008 ) ;
assign n7010 =  ( n6802 ) ? ( bv_8_110_n294 ) : ( n7009 ) ;
assign n7011 =  ( n6800 ) ? ( bv_8_90_n25 ) : ( n7010 ) ;
assign n7012 =  ( n6798 ) ? ( bv_8_160_n350 ) : ( n7011 ) ;
assign n7013 =  ( n6796 ) ? ( bv_8_82_n578 ) : ( n7012 ) ;
assign n7014 =  ( n6794 ) ? ( bv_8_59_n382 ) : ( n7013 ) ;
assign n7015 =  ( n6792 ) ? ( bv_8_214_n164 ) : ( n7014 ) ;
assign n7016 =  ( n6790 ) ? ( bv_8_179_n289 ) : ( n7015 ) ;
assign n7017 =  ( n6788 ) ? ( bv_8_41_n29 ) : ( n7016 ) ;
assign n7018 =  ( n6786 ) ? ( bv_8_227_n115 ) : ( n7017 ) ;
assign n7019 =  ( n6784 ) ? ( bv_8_47_n652 ) : ( n7018 ) ;
assign n7020 =  ( n6782 ) ? ( bv_8_132_n41 ) : ( n7019 ) ;
assign n7021 =  ( n6780 ) ? ( bv_8_83_n575 ) : ( n7020 ) ;
assign n7022 =  ( n6778 ) ? ( bv_8_209_n182 ) : ( n7021 ) ;
assign n7023 =  ( n6776 ) ? ( bv_8_0_n580 ) : ( n7022 ) ;
assign n7024 =  ( n6774 ) ? ( bv_8_237_n75 ) : ( n7023 ) ;
assign n7025 =  ( n6772 ) ? ( bv_8_32_n463 ) : ( n7024 ) ;
assign n7026 =  ( n6770 ) ? ( bv_8_252_n15 ) : ( n7025 ) ;
assign n7027 =  ( n6768 ) ? ( bv_8_177_n283 ) : ( n7026 ) ;
assign n7028 =  ( n6766 ) ? ( bv_8_91_n555 ) : ( n7027 ) ;
assign n7029 =  ( n6764 ) ? ( bv_8_106_n155 ) : ( n7028 ) ;
assign n7030 =  ( n6762 ) ? ( bv_8_203_n203 ) : ( n7029 ) ;
assign n7031 =  ( n6760 ) ? ( bv_8_190_n250 ) : ( n7030 ) ;
assign n7032 =  ( n6758 ) ? ( bv_8_57_n312 ) : ( n7031 ) ;
assign n7033 =  ( n6756 ) ? ( bv_8_74_n237 ) : ( n7032 ) ;
assign n7034 =  ( n6754 ) ? ( bv_8_76_n596 ) : ( n7033 ) ;
assign n7035 =  ( n6752 ) ? ( bv_8_88_n562 ) : ( n7034 ) ;
assign n7036 =  ( n6750 ) ? ( bv_8_207_n188 ) : ( n7035 ) ;
assign n7037 =  ( n6748 ) ? ( bv_8_208_n37 ) : ( n7036 ) ;
assign n7038 =  ( n6746 ) ? ( bv_8_239_n67 ) : ( n7037 ) ;
assign n7039 =  ( n6744 ) ? ( bv_8_170_n77 ) : ( n7038 ) ;
assign n7040 =  ( n6742 ) ? ( bv_8_251_n19 ) : ( n7039 ) ;
assign n7041 =  ( n6740 ) ? ( bv_8_67_n318 ) : ( n7040 ) ;
assign n7042 =  ( n6738 ) ? ( bv_8_77_n593 ) : ( n7041 ) ;
assign n7043 =  ( n6736 ) ? ( bv_8_51_n101 ) : ( n7042 ) ;
assign n7044 =  ( n6734 ) ? ( bv_8_133_n434 ) : ( n7043 ) ;
assign n7045 =  ( n6732 ) ? ( bv_8_69_n612 ) : ( n7044 ) ;
assign n7046 =  ( n6730 ) ? ( bv_8_249_n27 ) : ( n7045 ) ;
assign n7047 =  ( n6728 ) ? ( bv_8_2_n751 ) : ( n7046 ) ;
assign n7048 =  ( n6726 ) ? ( bv_8_127_n453 ) : ( n7047 ) ;
assign n7049 =  ( n6724 ) ? ( bv_8_80_n73 ) : ( n7048 ) ;
assign n7050 =  ( n6722 ) ? ( bv_8_60_n93 ) : ( n7049 ) ;
assign n7051 =  ( n6720 ) ? ( bv_8_159_n323 ) : ( n7050 ) ;
assign n7052 =  ( n6718 ) ? ( bv_8_168_n13 ) : ( n7051 ) ;
assign n7053 =  ( n6716 ) ? ( bv_8_81_n582 ) : ( n7052 ) ;
assign n7054 =  ( n6714 ) ? ( bv_8_163_n339 ) : ( n7053 ) ;
assign n7055 =  ( n6712 ) ? ( bv_8_64_n573 ) : ( n7054 ) ;
assign n7056 =  ( n6710 ) ? ( bv_8_143_n403 ) : ( n7055 ) ;
assign n7057 =  ( n6708 ) ? ( bv_8_146_n337 ) : ( n7056 ) ;
assign n7058 =  ( n6706 ) ? ( bv_8_157_n359 ) : ( n7057 ) ;
assign n7059 =  ( n6704 ) ? ( bv_8_56_n230 ) : ( n7058 ) ;
assign n7060 =  ( n6702 ) ? ( bv_8_245_n43 ) : ( n7059 ) ;
assign n7061 =  ( n6700 ) ? ( bv_8_188_n257 ) : ( n7060 ) ;
assign n7062 =  ( n6698 ) ? ( bv_8_182_n277 ) : ( n7061 ) ;
assign n7063 =  ( n6696 ) ? ( bv_8_218_n150 ) : ( n7062 ) ;
assign n7064 =  ( n6694 ) ? ( bv_8_33_n486 ) : ( n7063 ) ;
assign n7065 =  ( n6692 ) ? ( bv_8_16_n248 ) : ( n7064 ) ;
assign n7066 =  ( n6690 ) ? ( bv_8_255_n3 ) : ( n7065 ) ;
assign n7067 =  ( n6688 ) ? ( bv_8_243_n51 ) : ( n7066 ) ;
assign n7068 =  ( n6686 ) ? ( bv_8_210_n113 ) : ( n7067 ) ;
assign n7069 =  ( n6684 ) ? ( bv_8_205_n196 ) : ( n7068 ) ;
assign n7070 =  ( n6682 ) ? ( bv_8_12_n333 ) : ( n7069 ) ;
assign n7071 =  ( n6680 ) ? ( bv_8_19_n588 ) : ( n7070 ) ;
assign n7072 =  ( n6678 ) ? ( bv_8_236_n79 ) : ( n7071 ) ;
assign n7073 =  ( n6676 ) ? ( bv_8_95_n545 ) : ( n7072 ) ;
assign n7074 =  ( n6674 ) ? ( bv_8_151_n218 ) : ( n7073 ) ;
assign n7075 =  ( n6672 ) ? ( bv_8_68_n390 ) : ( n7074 ) ;
assign n7076 =  ( n6670 ) ? ( bv_8_23_n144 ) : ( n7075 ) ;
assign n7077 =  ( n6668 ) ? ( bv_8_196_n228 ) : ( n7076 ) ;
assign n7078 =  ( n6666 ) ? ( bv_8_167_n325 ) : ( n7077 ) ;
assign n7079 =  ( n6664 ) ? ( bv_8_126_n456 ) : ( n7078 ) ;
assign n7080 =  ( n6662 ) ? ( bv_8_61_n634 ) : ( n7079 ) ;
assign n7081 =  ( n6660 ) ? ( bv_8_100_n348 ) : ( n7080 ) ;
assign n7082 =  ( n6658 ) ? ( bv_8_93_n498 ) : ( n7081 ) ;
assign n7083 =  ( n6656 ) ? ( bv_8_25_n399 ) : ( n7082 ) ;
assign n7084 =  ( n6654 ) ? ( bv_8_115_n222 ) : ( n7083 ) ;
assign n7085 =  ( n6652 ) ? ( bv_8_96_n542 ) : ( n7084 ) ;
assign n7086 =  ( n6650 ) ? ( bv_8_129_n446 ) : ( n7085 ) ;
assign n7087 =  ( n6648 ) ? ( bv_8_79_n538 ) : ( n7086 ) ;
assign n7088 =  ( n6646 ) ? ( bv_8_220_n142 ) : ( n7087 ) ;
assign n7089 =  ( n6644 ) ? ( bv_8_34_n117 ) : ( n7088 ) ;
assign n7090 =  ( n6642 ) ? ( bv_8_42_n672 ) : ( n7089 ) ;
assign n7091 =  ( n6640 ) ? ( bv_8_144_n173 ) : ( n7090 ) ;
assign n7092 =  ( n6638 ) ? ( bv_8_136_n425 ) : ( n7091 ) ;
assign n7093 =  ( n6636 ) ? ( bv_8_70_n609 ) : ( n7092 ) ;
assign n7094 =  ( n6634 ) ? ( bv_8_238_n71 ) : ( n7093 ) ;
assign n7095 =  ( n6632 ) ? ( bv_8_184_n270 ) : ( n7094 ) ;
assign n7096 =  ( n6630 ) ? ( bv_8_20_n341 ) : ( n7095 ) ;
assign n7097 =  ( n6628 ) ? ( bv_8_222_n134 ) : ( n7096 ) ;
assign n7098 =  ( n6626 ) ? ( bv_8_94_n548 ) : ( n7097 ) ;
assign n7099 =  ( n6624 ) ? ( bv_8_11_n379 ) : ( n7098 ) ;
assign n7100 =  ( n6622 ) ? ( bv_8_219_n146 ) : ( n7099 ) ;
assign n7101 =  ( n6620 ) ? ( bv_8_224_n126 ) : ( n7100 ) ;
assign n7102 =  ( n6618 ) ? ( bv_8_50_n408 ) : ( n7101 ) ;
assign n7103 =  ( n6616 ) ? ( bv_8_58_n136 ) : ( n7102 ) ;
assign n7104 =  ( n6614 ) ? ( bv_8_10_n655 ) : ( n7103 ) ;
assign n7105 =  ( n6612 ) ? ( bv_8_73_n275 ) : ( n7104 ) ;
assign n7106 =  ( n6610 ) ? ( bv_8_6_n169 ) : ( n7105 ) ;
assign n7107 =  ( n6608 ) ? ( bv_8_36_n645 ) : ( n7106 ) ;
assign n7108 =  ( n6606 ) ? ( bv_8_92_n234 ) : ( n7107 ) ;
assign n7109 =  ( n6604 ) ? ( bv_8_194_n159 ) : ( n7108 ) ;
assign n7110 =  ( n6602 ) ? ( bv_8_211_n175 ) : ( n7109 ) ;
assign n7111 =  ( n6600 ) ? ( bv_8_172_n268 ) : ( n7110 ) ;
assign n7112 =  ( n6598 ) ? ( bv_8_98_n536 ) : ( n7111 ) ;
assign n7113 =  ( n6596 ) ? ( bv_8_145_n397 ) : ( n7112 ) ;
assign n7114 =  ( n6594 ) ? ( bv_8_149_n384 ) : ( n7113 ) ;
assign n7115 =  ( n6592 ) ? ( bv_8_228_n111 ) : ( n7114 ) ;
assign n7116 =  ( n6590 ) ? ( bv_8_121_n470 ) : ( n7115 ) ;
assign n7117 =  ( n6588 ) ? ( bv_8_231_n99 ) : ( n7116 ) ;
assign n7118 =  ( n6586 ) ? ( bv_8_200_n213 ) : ( n7117 ) ;
assign n7119 =  ( n6584 ) ? ( bv_8_55_n650 ) : ( n7118 ) ;
assign n7120 =  ( n6582 ) ? ( bv_8_109_n9 ) : ( n7119 ) ;
assign n7121 =  ( n6580 ) ? ( bv_8_141_n410 ) : ( n7120 ) ;
assign n7122 =  ( n6578 ) ? ( bv_8_213_n167 ) : ( n7121 ) ;
assign n7123 =  ( n6576 ) ? ( bv_8_78_n590 ) : ( n7122 ) ;
assign n7124 =  ( n6574 ) ? ( bv_8_169_n109 ) : ( n7123 ) ;
assign n7125 =  ( n6572 ) ? ( bv_8_108_n510 ) : ( n7124 ) ;
assign n7126 =  ( n6570 ) ? ( bv_8_86_n567 ) : ( n7125 ) ;
assign n7127 =  ( n6568 ) ? ( bv_8_244_n47 ) : ( n7126 ) ;
assign n7128 =  ( n6566 ) ? ( bv_8_234_n87 ) : ( n7127 ) ;
assign n7129 =  ( n6564 ) ? ( bv_8_101_n49 ) : ( n7128 ) ;
assign n7130 =  ( n6562 ) ? ( bv_8_122_n416 ) : ( n7129 ) ;
assign n7131 =  ( n6560 ) ? ( bv_8_174_n152 ) : ( n7130 ) ;
assign n7132 =  ( n6558 ) ? ( bv_8_8_n669 ) : ( n7131 ) ;
assign n7133 =  ( n6556 ) ? ( bv_8_186_n263 ) : ( n7132 ) ;
assign n7134 =  ( n6554 ) ? ( bv_8_120_n474 ) : ( n7133 ) ;
assign n7135 =  ( n6552 ) ? ( bv_8_37_n506 ) : ( n7134 ) ;
assign n7136 =  ( n6550 ) ? ( bv_8_46_n429 ) : ( n7135 ) ;
assign n7137 =  ( n6548 ) ? ( bv_8_28_n162 ) : ( n7136 ) ;
assign n7138 =  ( n6546 ) ? ( bv_8_166_n328 ) : ( n7137 ) ;
assign n7139 =  ( n6544 ) ? ( bv_8_180_n285 ) : ( n7138 ) ;
assign n7140 =  ( n6542 ) ? ( bv_8_198_n220 ) : ( n7139 ) ;
assign n7141 =  ( n6540 ) ? ( bv_8_232_n95 ) : ( n7140 ) ;
assign n7142 =  ( n6538 ) ? ( bv_8_221_n138 ) : ( n7141 ) ;
assign n7143 =  ( n6536 ) ? ( bv_8_116_n345 ) : ( n7142 ) ;
assign n7144 =  ( n6534 ) ? ( bv_8_31_n705 ) : ( n7143 ) ;
assign n7145 =  ( n6532 ) ? ( bv_8_75_n503 ) : ( n7144 ) ;
assign n7146 =  ( n6530 ) ? ( bv_8_189_n254 ) : ( n7145 ) ;
assign n7147 =  ( n6528 ) ? ( bv_8_139_n297 ) : ( n7146 ) ;
assign n7148 =  ( n6526 ) ? ( bv_8_138_n418 ) : ( n7147 ) ;
assign n7149 =  ( n6524 ) ? ( bv_8_112_n482 ) : ( n7148 ) ;
assign n7150 =  ( n6522 ) ? ( bv_8_62_n205 ) : ( n7149 ) ;
assign n7151 =  ( n6520 ) ? ( bv_8_181_n281 ) : ( n7150 ) ;
assign n7152 =  ( n6518 ) ? ( bv_8_102_n527 ) : ( n7151 ) ;
assign n7153 =  ( n6516 ) ? ( bv_8_72_n330 ) : ( n7152 ) ;
assign n7154 =  ( n6514 ) ? ( bv_8_3_n65 ) : ( n7153 ) ;
assign n7155 =  ( n6512 ) ? ( bv_8_246_n39 ) : ( n7154 ) ;
assign n7156 =  ( n6510 ) ? ( bv_8_14_n648 ) : ( n7155 ) ;
assign n7157 =  ( n6508 ) ? ( bv_8_97_n198 ) : ( n7156 ) ;
assign n7158 =  ( n6506 ) ? ( bv_8_53_n436 ) : ( n7157 ) ;
assign n7159 =  ( n6504 ) ? ( bv_8_87_n226 ) : ( n7158 ) ;
assign n7160 =  ( n6502 ) ? ( bv_8_185_n266 ) : ( n7159 ) ;
assign n7161 =  ( n6500 ) ? ( bv_8_134_n431 ) : ( n7160 ) ;
assign n7162 =  ( n6498 ) ? ( bv_8_193_n239 ) : ( n7161 ) ;
assign n7163 =  ( n6496 ) ? ( bv_8_29_n625 ) : ( n7162 ) ;
assign n7164 =  ( n6494 ) ? ( bv_8_158_n355 ) : ( n7163 ) ;
assign n7165 =  ( n6492 ) ? ( bv_8_225_n123 ) : ( n7164 ) ;
assign n7166 =  ( n6490 ) ? ( bv_8_248_n31 ) : ( n7165 ) ;
assign n7167 =  ( n6488 ) ? ( bv_8_152_n374 ) : ( n7166 ) ;
assign n7168 =  ( n6486 ) ? ( bv_8_17_n525 ) : ( n7167 ) ;
assign n7169 =  ( n6484 ) ? ( bv_8_105_n148 ) : ( n7168 ) ;
assign n7170 =  ( n6482 ) ? ( bv_8_217_n128 ) : ( n7169 ) ;
assign n7171 =  ( n6480 ) ? ( bv_8_142_n406 ) : ( n7170 ) ;
assign n7172 =  ( n6478 ) ? ( bv_8_148_n388 ) : ( n7171 ) ;
assign n7173 =  ( n6476 ) ? ( bv_8_155_n364 ) : ( n7172 ) ;
assign n7174 =  ( n6474 ) ? ( bv_8_30_n21 ) : ( n7173 ) ;
assign n7175 =  ( n6472 ) ? ( bv_8_135_n81 ) : ( n7174 ) ;
assign n7176 =  ( n6470 ) ? ( bv_8_233_n91 ) : ( n7175 ) ;
assign n7177 =  ( n6468 ) ? ( bv_8_206_n192 ) : ( n7176 ) ;
assign n7178 =  ( n6466 ) ? ( bv_8_85_n423 ) : ( n7177 ) ;
assign n7179 =  ( n6464 ) ? ( bv_8_40_n366 ) : ( n7178 ) ;
assign n7180 =  ( n6462 ) ? ( bv_8_223_n130 ) : ( n7179 ) ;
assign n7181 =  ( n6460 ) ? ( bv_8_140_n376 ) : ( n7180 ) ;
assign n7182 =  ( n6458 ) ? ( bv_8_161_n211 ) : ( n7181 ) ;
assign n7183 =  ( n6456 ) ? ( bv_8_137_n421 ) : ( n7182 ) ;
assign n7184 =  ( n6454 ) ? ( bv_8_13_n194 ) : ( n7183 ) ;
assign n7185 =  ( n6452 ) ? ( bv_8_191_n246 ) : ( n7184 ) ;
assign n7186 =  ( n6450 ) ? ( bv_8_230_n103 ) : ( n7185 ) ;
assign n7187 =  ( n6448 ) ? ( bv_8_66_n466 ) : ( n7186 ) ;
assign n7188 =  ( n6446 ) ? ( bv_8_104_n520 ) : ( n7187 ) ;
assign n7189 =  ( n6444 ) ? ( bv_8_65_n623 ) : ( n7188 ) ;
assign n7190 =  ( n6442 ) ? ( bv_8_153_n140 ) : ( n7189 ) ;
assign n7191 =  ( n6440 ) ? ( bv_8_45_n97 ) : ( n7190 ) ;
assign n7192 =  ( n6438 ) ? ( bv_8_15_n190 ) : ( n7191 ) ;
assign n7193 =  ( n6436 ) ? ( bv_8_176_n299 ) : ( n7192 ) ;
assign n7194 =  ( n6434 ) ? ( bv_8_84_n386 ) : ( n7193 ) ;
assign n7195 =  ( n6432 ) ? ( bv_8_187_n260 ) : ( n7194 ) ;
assign n7196 =  ( n6430 ) ? ( bv_8_22_n357 ) : ( n7195 ) ;
assign n7197 = state_in[95:88] ;
assign n7198 =  ( n7197 ) == ( bv_8_255_n3 )  ;
assign n7199 = state_in[95:88] ;
assign n7200 =  ( n7199 ) == ( bv_8_254_n7 )  ;
assign n7201 = state_in[95:88] ;
assign n7202 =  ( n7201 ) == ( bv_8_253_n11 )  ;
assign n7203 = state_in[95:88] ;
assign n7204 =  ( n7203 ) == ( bv_8_252_n15 )  ;
assign n7205 = state_in[95:88] ;
assign n7206 =  ( n7205 ) == ( bv_8_251_n19 )  ;
assign n7207 = state_in[95:88] ;
assign n7208 =  ( n7207 ) == ( bv_8_250_n23 )  ;
assign n7209 = state_in[95:88] ;
assign n7210 =  ( n7209 ) == ( bv_8_249_n27 )  ;
assign n7211 = state_in[95:88] ;
assign n7212 =  ( n7211 ) == ( bv_8_248_n31 )  ;
assign n7213 = state_in[95:88] ;
assign n7214 =  ( n7213 ) == ( bv_8_247_n35 )  ;
assign n7215 = state_in[95:88] ;
assign n7216 =  ( n7215 ) == ( bv_8_246_n39 )  ;
assign n7217 = state_in[95:88] ;
assign n7218 =  ( n7217 ) == ( bv_8_245_n43 )  ;
assign n7219 = state_in[95:88] ;
assign n7220 =  ( n7219 ) == ( bv_8_244_n47 )  ;
assign n7221 = state_in[95:88] ;
assign n7222 =  ( n7221 ) == ( bv_8_243_n51 )  ;
assign n7223 = state_in[95:88] ;
assign n7224 =  ( n7223 ) == ( bv_8_242_n55 )  ;
assign n7225 = state_in[95:88] ;
assign n7226 =  ( n7225 ) == ( bv_8_241_n59 )  ;
assign n7227 = state_in[95:88] ;
assign n7228 =  ( n7227 ) == ( bv_8_240_n63 )  ;
assign n7229 = state_in[95:88] ;
assign n7230 =  ( n7229 ) == ( bv_8_239_n67 )  ;
assign n7231 = state_in[95:88] ;
assign n7232 =  ( n7231 ) == ( bv_8_238_n71 )  ;
assign n7233 = state_in[95:88] ;
assign n7234 =  ( n7233 ) == ( bv_8_237_n75 )  ;
assign n7235 = state_in[95:88] ;
assign n7236 =  ( n7235 ) == ( bv_8_236_n79 )  ;
assign n7237 = state_in[95:88] ;
assign n7238 =  ( n7237 ) == ( bv_8_235_n83 )  ;
assign n7239 = state_in[95:88] ;
assign n7240 =  ( n7239 ) == ( bv_8_234_n87 )  ;
assign n7241 = state_in[95:88] ;
assign n7242 =  ( n7241 ) == ( bv_8_233_n91 )  ;
assign n7243 = state_in[95:88] ;
assign n7244 =  ( n7243 ) == ( bv_8_232_n95 )  ;
assign n7245 = state_in[95:88] ;
assign n7246 =  ( n7245 ) == ( bv_8_231_n99 )  ;
assign n7247 = state_in[95:88] ;
assign n7248 =  ( n7247 ) == ( bv_8_230_n103 )  ;
assign n7249 = state_in[95:88] ;
assign n7250 =  ( n7249 ) == ( bv_8_229_n107 )  ;
assign n7251 = state_in[95:88] ;
assign n7252 =  ( n7251 ) == ( bv_8_228_n111 )  ;
assign n7253 = state_in[95:88] ;
assign n7254 =  ( n7253 ) == ( bv_8_227_n115 )  ;
assign n7255 = state_in[95:88] ;
assign n7256 =  ( n7255 ) == ( bv_8_226_n119 )  ;
assign n7257 = state_in[95:88] ;
assign n7258 =  ( n7257 ) == ( bv_8_225_n123 )  ;
assign n7259 = state_in[95:88] ;
assign n7260 =  ( n7259 ) == ( bv_8_224_n126 )  ;
assign n7261 = state_in[95:88] ;
assign n7262 =  ( n7261 ) == ( bv_8_223_n130 )  ;
assign n7263 = state_in[95:88] ;
assign n7264 =  ( n7263 ) == ( bv_8_222_n134 )  ;
assign n7265 = state_in[95:88] ;
assign n7266 =  ( n7265 ) == ( bv_8_221_n138 )  ;
assign n7267 = state_in[95:88] ;
assign n7268 =  ( n7267 ) == ( bv_8_220_n142 )  ;
assign n7269 = state_in[95:88] ;
assign n7270 =  ( n7269 ) == ( bv_8_219_n146 )  ;
assign n7271 = state_in[95:88] ;
assign n7272 =  ( n7271 ) == ( bv_8_218_n150 )  ;
assign n7273 = state_in[95:88] ;
assign n7274 =  ( n7273 ) == ( bv_8_217_n128 )  ;
assign n7275 = state_in[95:88] ;
assign n7276 =  ( n7275 ) == ( bv_8_216_n157 )  ;
assign n7277 = state_in[95:88] ;
assign n7278 =  ( n7277 ) == ( bv_8_215_n45 )  ;
assign n7279 = state_in[95:88] ;
assign n7280 =  ( n7279 ) == ( bv_8_214_n164 )  ;
assign n7281 = state_in[95:88] ;
assign n7282 =  ( n7281 ) == ( bv_8_213_n167 )  ;
assign n7283 = state_in[95:88] ;
assign n7284 =  ( n7283 ) == ( bv_8_212_n171 )  ;
assign n7285 = state_in[95:88] ;
assign n7286 =  ( n7285 ) == ( bv_8_211_n175 )  ;
assign n7287 = state_in[95:88] ;
assign n7288 =  ( n7287 ) == ( bv_8_210_n113 )  ;
assign n7289 = state_in[95:88] ;
assign n7290 =  ( n7289 ) == ( bv_8_209_n182 )  ;
assign n7291 = state_in[95:88] ;
assign n7292 =  ( n7291 ) == ( bv_8_208_n37 )  ;
assign n7293 = state_in[95:88] ;
assign n7294 =  ( n7293 ) == ( bv_8_207_n188 )  ;
assign n7295 = state_in[95:88] ;
assign n7296 =  ( n7295 ) == ( bv_8_206_n192 )  ;
assign n7297 = state_in[95:88] ;
assign n7298 =  ( n7297 ) == ( bv_8_205_n196 )  ;
assign n7299 = state_in[95:88] ;
assign n7300 =  ( n7299 ) == ( bv_8_204_n177 )  ;
assign n7301 = state_in[95:88] ;
assign n7302 =  ( n7301 ) == ( bv_8_203_n203 )  ;
assign n7303 = state_in[95:88] ;
assign n7304 =  ( n7303 ) == ( bv_8_202_n207 )  ;
assign n7305 = state_in[95:88] ;
assign n7306 =  ( n7305 ) == ( bv_8_201_n85 )  ;
assign n7307 = state_in[95:88] ;
assign n7308 =  ( n7307 ) == ( bv_8_200_n213 )  ;
assign n7309 = state_in[95:88] ;
assign n7310 =  ( n7309 ) == ( bv_8_199_n216 )  ;
assign n7311 = state_in[95:88] ;
assign n7312 =  ( n7311 ) == ( bv_8_198_n220 )  ;
assign n7313 = state_in[95:88] ;
assign n7314 =  ( n7313 ) == ( bv_8_197_n224 )  ;
assign n7315 = state_in[95:88] ;
assign n7316 =  ( n7315 ) == ( bv_8_196_n228 )  ;
assign n7317 = state_in[95:88] ;
assign n7318 =  ( n7317 ) == ( bv_8_195_n232 )  ;
assign n7319 = state_in[95:88] ;
assign n7320 =  ( n7319 ) == ( bv_8_194_n159 )  ;
assign n7321 = state_in[95:88] ;
assign n7322 =  ( n7321 ) == ( bv_8_193_n239 )  ;
assign n7323 = state_in[95:88] ;
assign n7324 =  ( n7323 ) == ( bv_8_192_n242 )  ;
assign n7325 = state_in[95:88] ;
assign n7326 =  ( n7325 ) == ( bv_8_191_n246 )  ;
assign n7327 = state_in[95:88] ;
assign n7328 =  ( n7327 ) == ( bv_8_190_n250 )  ;
assign n7329 = state_in[95:88] ;
assign n7330 =  ( n7329 ) == ( bv_8_189_n254 )  ;
assign n7331 = state_in[95:88] ;
assign n7332 =  ( n7331 ) == ( bv_8_188_n257 )  ;
assign n7333 = state_in[95:88] ;
assign n7334 =  ( n7333 ) == ( bv_8_187_n260 )  ;
assign n7335 = state_in[95:88] ;
assign n7336 =  ( n7335 ) == ( bv_8_186_n263 )  ;
assign n7337 = state_in[95:88] ;
assign n7338 =  ( n7337 ) == ( bv_8_185_n266 )  ;
assign n7339 = state_in[95:88] ;
assign n7340 =  ( n7339 ) == ( bv_8_184_n270 )  ;
assign n7341 = state_in[95:88] ;
assign n7342 =  ( n7341 ) == ( bv_8_183_n273 )  ;
assign n7343 = state_in[95:88] ;
assign n7344 =  ( n7343 ) == ( bv_8_182_n277 )  ;
assign n7345 = state_in[95:88] ;
assign n7346 =  ( n7345 ) == ( bv_8_181_n281 )  ;
assign n7347 = state_in[95:88] ;
assign n7348 =  ( n7347 ) == ( bv_8_180_n285 )  ;
assign n7349 = state_in[95:88] ;
assign n7350 =  ( n7349 ) == ( bv_8_179_n289 )  ;
assign n7351 = state_in[95:88] ;
assign n7352 =  ( n7351 ) == ( bv_8_178_n292 )  ;
assign n7353 = state_in[95:88] ;
assign n7354 =  ( n7353 ) == ( bv_8_177_n283 )  ;
assign n7355 = state_in[95:88] ;
assign n7356 =  ( n7355 ) == ( bv_8_176_n299 )  ;
assign n7357 = state_in[95:88] ;
assign n7358 =  ( n7357 ) == ( bv_8_175_n302 )  ;
assign n7359 = state_in[95:88] ;
assign n7360 =  ( n7359 ) == ( bv_8_174_n152 )  ;
assign n7361 = state_in[95:88] ;
assign n7362 =  ( n7361 ) == ( bv_8_173_n307 )  ;
assign n7363 = state_in[95:88] ;
assign n7364 =  ( n7363 ) == ( bv_8_172_n268 )  ;
assign n7365 = state_in[95:88] ;
assign n7366 =  ( n7365 ) == ( bv_8_171_n314 )  ;
assign n7367 = state_in[95:88] ;
assign n7368 =  ( n7367 ) == ( bv_8_170_n77 )  ;
assign n7369 = state_in[95:88] ;
assign n7370 =  ( n7369 ) == ( bv_8_169_n109 )  ;
assign n7371 = state_in[95:88] ;
assign n7372 =  ( n7371 ) == ( bv_8_168_n13 )  ;
assign n7373 = state_in[95:88] ;
assign n7374 =  ( n7373 ) == ( bv_8_167_n325 )  ;
assign n7375 = state_in[95:88] ;
assign n7376 =  ( n7375 ) == ( bv_8_166_n328 )  ;
assign n7377 = state_in[95:88] ;
assign n7378 =  ( n7377 ) == ( bv_8_165_n69 )  ;
assign n7379 = state_in[95:88] ;
assign n7380 =  ( n7379 ) == ( bv_8_164_n335 )  ;
assign n7381 = state_in[95:88] ;
assign n7382 =  ( n7381 ) == ( bv_8_163_n339 )  ;
assign n7383 = state_in[95:88] ;
assign n7384 =  ( n7383 ) == ( bv_8_162_n343 )  ;
assign n7385 = state_in[95:88] ;
assign n7386 =  ( n7385 ) == ( bv_8_161_n211 )  ;
assign n7387 = state_in[95:88] ;
assign n7388 =  ( n7387 ) == ( bv_8_160_n350 )  ;
assign n7389 = state_in[95:88] ;
assign n7390 =  ( n7389 ) == ( bv_8_159_n323 )  ;
assign n7391 = state_in[95:88] ;
assign n7392 =  ( n7391 ) == ( bv_8_158_n355 )  ;
assign n7393 = state_in[95:88] ;
assign n7394 =  ( n7393 ) == ( bv_8_157_n359 )  ;
assign n7395 = state_in[95:88] ;
assign n7396 =  ( n7395 ) == ( bv_8_156_n279 )  ;
assign n7397 = state_in[95:88] ;
assign n7398 =  ( n7397 ) == ( bv_8_155_n364 )  ;
assign n7399 = state_in[95:88] ;
assign n7400 =  ( n7399 ) == ( bv_8_154_n368 )  ;
assign n7401 = state_in[95:88] ;
assign n7402 =  ( n7401 ) == ( bv_8_153_n140 )  ;
assign n7403 = state_in[95:88] ;
assign n7404 =  ( n7403 ) == ( bv_8_152_n374 )  ;
assign n7405 = state_in[95:88] ;
assign n7406 =  ( n7405 ) == ( bv_8_151_n218 )  ;
assign n7407 = state_in[95:88] ;
assign n7408 =  ( n7407 ) == ( bv_8_150_n201 )  ;
assign n7409 = state_in[95:88] ;
assign n7410 =  ( n7409 ) == ( bv_8_149_n384 )  ;
assign n7411 = state_in[95:88] ;
assign n7412 =  ( n7411 ) == ( bv_8_148_n388 )  ;
assign n7413 = state_in[95:88] ;
assign n7414 =  ( n7413 ) == ( bv_8_147_n392 )  ;
assign n7415 = state_in[95:88] ;
assign n7416 =  ( n7415 ) == ( bv_8_146_n337 )  ;
assign n7417 = state_in[95:88] ;
assign n7418 =  ( n7417 ) == ( bv_8_145_n397 )  ;
assign n7419 = state_in[95:88] ;
assign n7420 =  ( n7419 ) == ( bv_8_144_n173 )  ;
assign n7421 = state_in[95:88] ;
assign n7422 =  ( n7421 ) == ( bv_8_143_n403 )  ;
assign n7423 = state_in[95:88] ;
assign n7424 =  ( n7423 ) == ( bv_8_142_n406 )  ;
assign n7425 = state_in[95:88] ;
assign n7426 =  ( n7425 ) == ( bv_8_141_n410 )  ;
assign n7427 = state_in[95:88] ;
assign n7428 =  ( n7427 ) == ( bv_8_140_n376 )  ;
assign n7429 = state_in[95:88] ;
assign n7430 =  ( n7429 ) == ( bv_8_139_n297 )  ;
assign n7431 = state_in[95:88] ;
assign n7432 =  ( n7431 ) == ( bv_8_138_n418 )  ;
assign n7433 = state_in[95:88] ;
assign n7434 =  ( n7433 ) == ( bv_8_137_n421 )  ;
assign n7435 = state_in[95:88] ;
assign n7436 =  ( n7435 ) == ( bv_8_136_n425 )  ;
assign n7437 = state_in[95:88] ;
assign n7438 =  ( n7437 ) == ( bv_8_135_n81 )  ;
assign n7439 = state_in[95:88] ;
assign n7440 =  ( n7439 ) == ( bv_8_134_n431 )  ;
assign n7441 = state_in[95:88] ;
assign n7442 =  ( n7441 ) == ( bv_8_133_n434 )  ;
assign n7443 = state_in[95:88] ;
assign n7444 =  ( n7443 ) == ( bv_8_132_n41 )  ;
assign n7445 = state_in[95:88] ;
assign n7446 =  ( n7445 ) == ( bv_8_131_n440 )  ;
assign n7447 = state_in[95:88] ;
assign n7448 =  ( n7447 ) == ( bv_8_130_n33 )  ;
assign n7449 = state_in[95:88] ;
assign n7450 =  ( n7449 ) == ( bv_8_129_n446 )  ;
assign n7451 = state_in[95:88] ;
assign n7452 =  ( n7451 ) == ( bv_8_128_n450 )  ;
assign n7453 = state_in[95:88] ;
assign n7454 =  ( n7453 ) == ( bv_8_127_n453 )  ;
assign n7455 = state_in[95:88] ;
assign n7456 =  ( n7455 ) == ( bv_8_126_n456 )  ;
assign n7457 = state_in[95:88] ;
assign n7458 =  ( n7457 ) == ( bv_8_125_n459 )  ;
assign n7459 = state_in[95:88] ;
assign n7460 =  ( n7459 ) == ( bv_8_124_n184 )  ;
assign n7461 = state_in[95:88] ;
assign n7462 =  ( n7461 ) == ( bv_8_123_n17 )  ;
assign n7463 = state_in[95:88] ;
assign n7464 =  ( n7463 ) == ( bv_8_122_n416 )  ;
assign n7465 = state_in[95:88] ;
assign n7466 =  ( n7465 ) == ( bv_8_121_n470 )  ;
assign n7467 = state_in[95:88] ;
assign n7468 =  ( n7467 ) == ( bv_8_120_n474 )  ;
assign n7469 = state_in[95:88] ;
assign n7470 =  ( n7469 ) == ( bv_8_119_n472 )  ;
assign n7471 = state_in[95:88] ;
assign n7472 =  ( n7471 ) == ( bv_8_118_n480 )  ;
assign n7473 = state_in[95:88] ;
assign n7474 =  ( n7473 ) == ( bv_8_117_n484 )  ;
assign n7475 = state_in[95:88] ;
assign n7476 =  ( n7475 ) == ( bv_8_116_n345 )  ;
assign n7477 = state_in[95:88] ;
assign n7478 =  ( n7477 ) == ( bv_8_115_n222 )  ;
assign n7479 = state_in[95:88] ;
assign n7480 =  ( n7479 ) == ( bv_8_114_n494 )  ;
assign n7481 = state_in[95:88] ;
assign n7482 =  ( n7481 ) == ( bv_8_113_n180 )  ;
assign n7483 = state_in[95:88] ;
assign n7484 =  ( n7483 ) == ( bv_8_112_n482 )  ;
assign n7485 = state_in[95:88] ;
assign n7486 =  ( n7485 ) == ( bv_8_111_n244 )  ;
assign n7487 = state_in[95:88] ;
assign n7488 =  ( n7487 ) == ( bv_8_110_n294 )  ;
assign n7489 = state_in[95:88] ;
assign n7490 =  ( n7489 ) == ( bv_8_109_n9 )  ;
assign n7491 = state_in[95:88] ;
assign n7492 =  ( n7491 ) == ( bv_8_108_n510 )  ;
assign n7493 = state_in[95:88] ;
assign n7494 =  ( n7493 ) == ( bv_8_107_n370 )  ;
assign n7495 = state_in[95:88] ;
assign n7496 =  ( n7495 ) == ( bv_8_106_n155 )  ;
assign n7497 = state_in[95:88] ;
assign n7498 =  ( n7497 ) == ( bv_8_105_n148 )  ;
assign n7499 = state_in[95:88] ;
assign n7500 =  ( n7499 ) == ( bv_8_104_n520 )  ;
assign n7501 = state_in[95:88] ;
assign n7502 =  ( n7501 ) == ( bv_8_103_n523 )  ;
assign n7503 = state_in[95:88] ;
assign n7504 =  ( n7503 ) == ( bv_8_102_n527 )  ;
assign n7505 = state_in[95:88] ;
assign n7506 =  ( n7505 ) == ( bv_8_101_n49 )  ;
assign n7507 = state_in[95:88] ;
assign n7508 =  ( n7507 ) == ( bv_8_100_n348 )  ;
assign n7509 = state_in[95:88] ;
assign n7510 =  ( n7509 ) == ( bv_8_99_n476 )  ;
assign n7511 = state_in[95:88] ;
assign n7512 =  ( n7511 ) == ( bv_8_98_n536 )  ;
assign n7513 = state_in[95:88] ;
assign n7514 =  ( n7513 ) == ( bv_8_97_n198 )  ;
assign n7515 = state_in[95:88] ;
assign n7516 =  ( n7515 ) == ( bv_8_96_n542 )  ;
assign n7517 = state_in[95:88] ;
assign n7518 =  ( n7517 ) == ( bv_8_95_n545 )  ;
assign n7519 = state_in[95:88] ;
assign n7520 =  ( n7519 ) == ( bv_8_94_n548 )  ;
assign n7521 = state_in[95:88] ;
assign n7522 =  ( n7521 ) == ( bv_8_93_n498 )  ;
assign n7523 = state_in[95:88] ;
assign n7524 =  ( n7523 ) == ( bv_8_92_n234 )  ;
assign n7525 = state_in[95:88] ;
assign n7526 =  ( n7525 ) == ( bv_8_91_n555 )  ;
assign n7527 = state_in[95:88] ;
assign n7528 =  ( n7527 ) == ( bv_8_90_n25 )  ;
assign n7529 = state_in[95:88] ;
assign n7530 =  ( n7529 ) == ( bv_8_89_n61 )  ;
assign n7531 = state_in[95:88] ;
assign n7532 =  ( n7531 ) == ( bv_8_88_n562 )  ;
assign n7533 = state_in[95:88] ;
assign n7534 =  ( n7533 ) == ( bv_8_87_n226 )  ;
assign n7535 = state_in[95:88] ;
assign n7536 =  ( n7535 ) == ( bv_8_86_n567 )  ;
assign n7537 = state_in[95:88] ;
assign n7538 =  ( n7537 ) == ( bv_8_85_n423 )  ;
assign n7539 = state_in[95:88] ;
assign n7540 =  ( n7539 ) == ( bv_8_84_n386 )  ;
assign n7541 = state_in[95:88] ;
assign n7542 =  ( n7541 ) == ( bv_8_83_n575 )  ;
assign n7543 = state_in[95:88] ;
assign n7544 =  ( n7543 ) == ( bv_8_82_n578 )  ;
assign n7545 = state_in[95:88] ;
assign n7546 =  ( n7545 ) == ( bv_8_81_n582 )  ;
assign n7547 = state_in[95:88] ;
assign n7548 =  ( n7547 ) == ( bv_8_80_n73 )  ;
assign n7549 = state_in[95:88] ;
assign n7550 =  ( n7549 ) == ( bv_8_79_n538 )  ;
assign n7551 = state_in[95:88] ;
assign n7552 =  ( n7551 ) == ( bv_8_78_n590 )  ;
assign n7553 = state_in[95:88] ;
assign n7554 =  ( n7553 ) == ( bv_8_77_n593 )  ;
assign n7555 = state_in[95:88] ;
assign n7556 =  ( n7555 ) == ( bv_8_76_n596 )  ;
assign n7557 = state_in[95:88] ;
assign n7558 =  ( n7557 ) == ( bv_8_75_n503 )  ;
assign n7559 = state_in[95:88] ;
assign n7560 =  ( n7559 ) == ( bv_8_74_n237 )  ;
assign n7561 = state_in[95:88] ;
assign n7562 =  ( n7561 ) == ( bv_8_73_n275 )  ;
assign n7563 = state_in[95:88] ;
assign n7564 =  ( n7563 ) == ( bv_8_72_n330 )  ;
assign n7565 = state_in[95:88] ;
assign n7566 =  ( n7565 ) == ( bv_8_71_n252 )  ;
assign n7567 = state_in[95:88] ;
assign n7568 =  ( n7567 ) == ( bv_8_70_n609 )  ;
assign n7569 = state_in[95:88] ;
assign n7570 =  ( n7569 ) == ( bv_8_69_n612 )  ;
assign n7571 = state_in[95:88] ;
assign n7572 =  ( n7571 ) == ( bv_8_68_n390 )  ;
assign n7573 = state_in[95:88] ;
assign n7574 =  ( n7573 ) == ( bv_8_67_n318 )  ;
assign n7575 = state_in[95:88] ;
assign n7576 =  ( n7575 ) == ( bv_8_66_n466 )  ;
assign n7577 = state_in[95:88] ;
assign n7578 =  ( n7577 ) == ( bv_8_65_n623 )  ;
assign n7579 = state_in[95:88] ;
assign n7580 =  ( n7579 ) == ( bv_8_64_n573 )  ;
assign n7581 = state_in[95:88] ;
assign n7582 =  ( n7581 ) == ( bv_8_63_n489 )  ;
assign n7583 = state_in[95:88] ;
assign n7584 =  ( n7583 ) == ( bv_8_62_n205 )  ;
assign n7585 = state_in[95:88] ;
assign n7586 =  ( n7585 ) == ( bv_8_61_n634 )  ;
assign n7587 = state_in[95:88] ;
assign n7588 =  ( n7587 ) == ( bv_8_60_n93 )  ;
assign n7589 = state_in[95:88] ;
assign n7590 =  ( n7589 ) == ( bv_8_59_n382 )  ;
assign n7591 = state_in[95:88] ;
assign n7592 =  ( n7591 ) == ( bv_8_58_n136 )  ;
assign n7593 = state_in[95:88] ;
assign n7594 =  ( n7593 ) == ( bv_8_57_n312 )  ;
assign n7595 = state_in[95:88] ;
assign n7596 =  ( n7595 ) == ( bv_8_56_n230 )  ;
assign n7597 = state_in[95:88] ;
assign n7598 =  ( n7597 ) == ( bv_8_55_n650 )  ;
assign n7599 = state_in[95:88] ;
assign n7600 =  ( n7599 ) == ( bv_8_54_n616 )  ;
assign n7601 = state_in[95:88] ;
assign n7602 =  ( n7601 ) == ( bv_8_53_n436 )  ;
assign n7603 = state_in[95:88] ;
assign n7604 =  ( n7603 ) == ( bv_8_52_n619 )  ;
assign n7605 = state_in[95:88] ;
assign n7606 =  ( n7605 ) == ( bv_8_51_n101 )  ;
assign n7607 = state_in[95:88] ;
assign n7608 =  ( n7607 ) == ( bv_8_50_n408 )  ;
assign n7609 = state_in[95:88] ;
assign n7610 =  ( n7609 ) == ( bv_8_49_n309 )  ;
assign n7611 = state_in[95:88] ;
assign n7612 =  ( n7611 ) == ( bv_8_48_n660 )  ;
assign n7613 = state_in[95:88] ;
assign n7614 =  ( n7613 ) == ( bv_8_47_n652 )  ;
assign n7615 = state_in[95:88] ;
assign n7616 =  ( n7615 ) == ( bv_8_46_n429 )  ;
assign n7617 = state_in[95:88] ;
assign n7618 =  ( n7617 ) == ( bv_8_45_n97 )  ;
assign n7619 = state_in[95:88] ;
assign n7620 =  ( n7619 ) == ( bv_8_44_n5 )  ;
assign n7621 = state_in[95:88] ;
assign n7622 =  ( n7621 ) == ( bv_8_43_n121 )  ;
assign n7623 = state_in[95:88] ;
assign n7624 =  ( n7623 ) == ( bv_8_42_n672 )  ;
assign n7625 = state_in[95:88] ;
assign n7626 =  ( n7625 ) == ( bv_8_41_n29 )  ;
assign n7627 = state_in[95:88] ;
assign n7628 =  ( n7627 ) == ( bv_8_40_n366 )  ;
assign n7629 = state_in[95:88] ;
assign n7630 =  ( n7629 ) == ( bv_8_39_n132 )  ;
assign n7631 = state_in[95:88] ;
assign n7632 =  ( n7631 ) == ( bv_8_38_n444 )  ;
assign n7633 = state_in[95:88] ;
assign n7634 =  ( n7633 ) == ( bv_8_37_n506 )  ;
assign n7635 = state_in[95:88] ;
assign n7636 =  ( n7635 ) == ( bv_8_36_n645 )  ;
assign n7637 = state_in[95:88] ;
assign n7638 =  ( n7637 ) == ( bv_8_35_n696 )  ;
assign n7639 = state_in[95:88] ;
assign n7640 =  ( n7639 ) == ( bv_8_34_n117 )  ;
assign n7641 = state_in[95:88] ;
assign n7642 =  ( n7641 ) == ( bv_8_33_n486 )  ;
assign n7643 = state_in[95:88] ;
assign n7644 =  ( n7643 ) == ( bv_8_32_n463 )  ;
assign n7645 = state_in[95:88] ;
assign n7646 =  ( n7645 ) == ( bv_8_31_n705 )  ;
assign n7647 = state_in[95:88] ;
assign n7648 =  ( n7647 ) == ( bv_8_30_n21 )  ;
assign n7649 = state_in[95:88] ;
assign n7650 =  ( n7649 ) == ( bv_8_29_n625 )  ;
assign n7651 = state_in[95:88] ;
assign n7652 =  ( n7651 ) == ( bv_8_28_n162 )  ;
assign n7653 = state_in[95:88] ;
assign n7654 =  ( n7653 ) == ( bv_8_27_n642 )  ;
assign n7655 = state_in[95:88] ;
assign n7656 =  ( n7655 ) == ( bv_8_26_n53 )  ;
assign n7657 = state_in[95:88] ;
assign n7658 =  ( n7657 ) == ( bv_8_25_n399 )  ;
assign n7659 = state_in[95:88] ;
assign n7660 =  ( n7659 ) == ( bv_8_24_n448 )  ;
assign n7661 = state_in[95:88] ;
assign n7662 =  ( n7661 ) == ( bv_8_23_n144 )  ;
assign n7663 = state_in[95:88] ;
assign n7664 =  ( n7663 ) == ( bv_8_22_n357 )  ;
assign n7665 = state_in[95:88] ;
assign n7666 =  ( n7665 ) == ( bv_8_21_n89 )  ;
assign n7667 = state_in[95:88] ;
assign n7668 =  ( n7667 ) == ( bv_8_20_n341 )  ;
assign n7669 = state_in[95:88] ;
assign n7670 =  ( n7669 ) == ( bv_8_19_n588 )  ;
assign n7671 = state_in[95:88] ;
assign n7672 =  ( n7671 ) == ( bv_8_18_n628 )  ;
assign n7673 = state_in[95:88] ;
assign n7674 =  ( n7673 ) == ( bv_8_17_n525 )  ;
assign n7675 = state_in[95:88] ;
assign n7676 =  ( n7675 ) == ( bv_8_16_n248 )  ;
assign n7677 = state_in[95:88] ;
assign n7678 =  ( n7677 ) == ( bv_8_15_n190 )  ;
assign n7679 = state_in[95:88] ;
assign n7680 =  ( n7679 ) == ( bv_8_14_n648 )  ;
assign n7681 = state_in[95:88] ;
assign n7682 =  ( n7681 ) == ( bv_8_13_n194 )  ;
assign n7683 = state_in[95:88] ;
assign n7684 =  ( n7683 ) == ( bv_8_12_n333 )  ;
assign n7685 = state_in[95:88] ;
assign n7686 =  ( n7685 ) == ( bv_8_11_n379 )  ;
assign n7687 = state_in[95:88] ;
assign n7688 =  ( n7687 ) == ( bv_8_10_n655 )  ;
assign n7689 = state_in[95:88] ;
assign n7690 =  ( n7689 ) == ( bv_8_9_n57 )  ;
assign n7691 = state_in[95:88] ;
assign n7692 =  ( n7691 ) == ( bv_8_8_n669 )  ;
assign n7693 = state_in[95:88] ;
assign n7694 =  ( n7693 ) == ( bv_8_7_n105 )  ;
assign n7695 = state_in[95:88] ;
assign n7696 =  ( n7695 ) == ( bv_8_6_n169 )  ;
assign n7697 = state_in[95:88] ;
assign n7698 =  ( n7697 ) == ( bv_8_5_n492 )  ;
assign n7699 = state_in[95:88] ;
assign n7700 =  ( n7699 ) == ( bv_8_4_n516 )  ;
assign n7701 = state_in[95:88] ;
assign n7702 =  ( n7701 ) == ( bv_8_3_n65 )  ;
assign n7703 = state_in[95:88] ;
assign n7704 =  ( n7703 ) == ( bv_8_2_n751 )  ;
assign n7705 = state_in[95:88] ;
assign n7706 =  ( n7705 ) == ( bv_8_1_n287 )  ;
assign n7707 = state_in[95:88] ;
assign n7708 =  ( n7707 ) == ( bv_8_0_n580 )  ;
assign n7709 =  ( n7708 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n7710 =  ( n7706 ) ? ( bv_8_248_n31 ) : ( n7709 ) ;
assign n7711 =  ( n7704 ) ? ( bv_8_238_n71 ) : ( n7710 ) ;
assign n7712 =  ( n7702 ) ? ( bv_8_246_n39 ) : ( n7711 ) ;
assign n7713 =  ( n7700 ) ? ( bv_8_255_n3 ) : ( n7712 ) ;
assign n7714 =  ( n7698 ) ? ( bv_8_214_n164 ) : ( n7713 ) ;
assign n7715 =  ( n7696 ) ? ( bv_8_222_n134 ) : ( n7714 ) ;
assign n7716 =  ( n7694 ) ? ( bv_8_145_n397 ) : ( n7715 ) ;
assign n7717 =  ( n7692 ) ? ( bv_8_96_n542 ) : ( n7716 ) ;
assign n7718 =  ( n7690 ) ? ( bv_8_2_n751 ) : ( n7717 ) ;
assign n7719 =  ( n7688 ) ? ( bv_8_206_n192 ) : ( n7718 ) ;
assign n7720 =  ( n7686 ) ? ( bv_8_86_n567 ) : ( n7719 ) ;
assign n7721 =  ( n7684 ) ? ( bv_8_231_n99 ) : ( n7720 ) ;
assign n7722 =  ( n7682 ) ? ( bv_8_181_n281 ) : ( n7721 ) ;
assign n7723 =  ( n7680 ) ? ( bv_8_77_n593 ) : ( n7722 ) ;
assign n7724 =  ( n7678 ) ? ( bv_8_236_n79 ) : ( n7723 ) ;
assign n7725 =  ( n7676 ) ? ( bv_8_143_n403 ) : ( n7724 ) ;
assign n7726 =  ( n7674 ) ? ( bv_8_31_n705 ) : ( n7725 ) ;
assign n7727 =  ( n7672 ) ? ( bv_8_137_n421 ) : ( n7726 ) ;
assign n7728 =  ( n7670 ) ? ( bv_8_250_n23 ) : ( n7727 ) ;
assign n7729 =  ( n7668 ) ? ( bv_8_239_n67 ) : ( n7728 ) ;
assign n7730 =  ( n7666 ) ? ( bv_8_178_n292 ) : ( n7729 ) ;
assign n7731 =  ( n7664 ) ? ( bv_8_142_n406 ) : ( n7730 ) ;
assign n7732 =  ( n7662 ) ? ( bv_8_251_n19 ) : ( n7731 ) ;
assign n7733 =  ( n7660 ) ? ( bv_8_65_n623 ) : ( n7732 ) ;
assign n7734 =  ( n7658 ) ? ( bv_8_179_n289 ) : ( n7733 ) ;
assign n7735 =  ( n7656 ) ? ( bv_8_95_n545 ) : ( n7734 ) ;
assign n7736 =  ( n7654 ) ? ( bv_8_69_n612 ) : ( n7735 ) ;
assign n7737 =  ( n7652 ) ? ( bv_8_35_n696 ) : ( n7736 ) ;
assign n7738 =  ( n7650 ) ? ( bv_8_83_n575 ) : ( n7737 ) ;
assign n7739 =  ( n7648 ) ? ( bv_8_228_n111 ) : ( n7738 ) ;
assign n7740 =  ( n7646 ) ? ( bv_8_155_n364 ) : ( n7739 ) ;
assign n7741 =  ( n7644 ) ? ( bv_8_117_n484 ) : ( n7740 ) ;
assign n7742 =  ( n7642 ) ? ( bv_8_225_n123 ) : ( n7741 ) ;
assign n7743 =  ( n7640 ) ? ( bv_8_61_n634 ) : ( n7742 ) ;
assign n7744 =  ( n7638 ) ? ( bv_8_76_n596 ) : ( n7743 ) ;
assign n7745 =  ( n7636 ) ? ( bv_8_108_n510 ) : ( n7744 ) ;
assign n7746 =  ( n7634 ) ? ( bv_8_126_n456 ) : ( n7745 ) ;
assign n7747 =  ( n7632 ) ? ( bv_8_245_n43 ) : ( n7746 ) ;
assign n7748 =  ( n7630 ) ? ( bv_8_131_n440 ) : ( n7747 ) ;
assign n7749 =  ( n7628 ) ? ( bv_8_104_n520 ) : ( n7748 ) ;
assign n7750 =  ( n7626 ) ? ( bv_8_81_n582 ) : ( n7749 ) ;
assign n7751 =  ( n7624 ) ? ( bv_8_209_n182 ) : ( n7750 ) ;
assign n7752 =  ( n7622 ) ? ( bv_8_249_n27 ) : ( n7751 ) ;
assign n7753 =  ( n7620 ) ? ( bv_8_226_n119 ) : ( n7752 ) ;
assign n7754 =  ( n7618 ) ? ( bv_8_171_n314 ) : ( n7753 ) ;
assign n7755 =  ( n7616 ) ? ( bv_8_98_n536 ) : ( n7754 ) ;
assign n7756 =  ( n7614 ) ? ( bv_8_42_n672 ) : ( n7755 ) ;
assign n7757 =  ( n7612 ) ? ( bv_8_8_n669 ) : ( n7756 ) ;
assign n7758 =  ( n7610 ) ? ( bv_8_149_n384 ) : ( n7757 ) ;
assign n7759 =  ( n7608 ) ? ( bv_8_70_n609 ) : ( n7758 ) ;
assign n7760 =  ( n7606 ) ? ( bv_8_157_n359 ) : ( n7759 ) ;
assign n7761 =  ( n7604 ) ? ( bv_8_48_n660 ) : ( n7760 ) ;
assign n7762 =  ( n7602 ) ? ( bv_8_55_n650 ) : ( n7761 ) ;
assign n7763 =  ( n7600 ) ? ( bv_8_10_n655 ) : ( n7762 ) ;
assign n7764 =  ( n7598 ) ? ( bv_8_47_n652 ) : ( n7763 ) ;
assign n7765 =  ( n7596 ) ? ( bv_8_14_n648 ) : ( n7764 ) ;
assign n7766 =  ( n7594 ) ? ( bv_8_36_n645 ) : ( n7765 ) ;
assign n7767 =  ( n7592 ) ? ( bv_8_27_n642 ) : ( n7766 ) ;
assign n7768 =  ( n7590 ) ? ( bv_8_223_n130 ) : ( n7767 ) ;
assign n7769 =  ( n7588 ) ? ( bv_8_205_n196 ) : ( n7768 ) ;
assign n7770 =  ( n7586 ) ? ( bv_8_78_n590 ) : ( n7769 ) ;
assign n7771 =  ( n7584 ) ? ( bv_8_127_n453 ) : ( n7770 ) ;
assign n7772 =  ( n7582 ) ? ( bv_8_234_n87 ) : ( n7771 ) ;
assign n7773 =  ( n7580 ) ? ( bv_8_18_n628 ) : ( n7772 ) ;
assign n7774 =  ( n7578 ) ? ( bv_8_29_n625 ) : ( n7773 ) ;
assign n7775 =  ( n7576 ) ? ( bv_8_88_n562 ) : ( n7774 ) ;
assign n7776 =  ( n7574 ) ? ( bv_8_52_n619 ) : ( n7775 ) ;
assign n7777 =  ( n7572 ) ? ( bv_8_54_n616 ) : ( n7776 ) ;
assign n7778 =  ( n7570 ) ? ( bv_8_220_n142 ) : ( n7777 ) ;
assign n7779 =  ( n7568 ) ? ( bv_8_180_n285 ) : ( n7778 ) ;
assign n7780 =  ( n7566 ) ? ( bv_8_91_n555 ) : ( n7779 ) ;
assign n7781 =  ( n7564 ) ? ( bv_8_164_n335 ) : ( n7780 ) ;
assign n7782 =  ( n7562 ) ? ( bv_8_118_n480 ) : ( n7781 ) ;
assign n7783 =  ( n7560 ) ? ( bv_8_183_n273 ) : ( n7782 ) ;
assign n7784 =  ( n7558 ) ? ( bv_8_125_n459 ) : ( n7783 ) ;
assign n7785 =  ( n7556 ) ? ( bv_8_82_n578 ) : ( n7784 ) ;
assign n7786 =  ( n7554 ) ? ( bv_8_221_n138 ) : ( n7785 ) ;
assign n7787 =  ( n7552 ) ? ( bv_8_94_n548 ) : ( n7786 ) ;
assign n7788 =  ( n7550 ) ? ( bv_8_19_n588 ) : ( n7787 ) ;
assign n7789 =  ( n7548 ) ? ( bv_8_166_n328 ) : ( n7788 ) ;
assign n7790 =  ( n7546 ) ? ( bv_8_185_n266 ) : ( n7789 ) ;
assign n7791 =  ( n7544 ) ? ( bv_8_0_n580 ) : ( n7790 ) ;
assign n7792 =  ( n7542 ) ? ( bv_8_193_n239 ) : ( n7791 ) ;
assign n7793 =  ( n7540 ) ? ( bv_8_64_n573 ) : ( n7792 ) ;
assign n7794 =  ( n7538 ) ? ( bv_8_227_n115 ) : ( n7793 ) ;
assign n7795 =  ( n7536 ) ? ( bv_8_121_n470 ) : ( n7794 ) ;
assign n7796 =  ( n7534 ) ? ( bv_8_182_n277 ) : ( n7795 ) ;
assign n7797 =  ( n7532 ) ? ( bv_8_212_n171 ) : ( n7796 ) ;
assign n7798 =  ( n7530 ) ? ( bv_8_141_n410 ) : ( n7797 ) ;
assign n7799 =  ( n7528 ) ? ( bv_8_103_n523 ) : ( n7798 ) ;
assign n7800 =  ( n7526 ) ? ( bv_8_114_n494 ) : ( n7799 ) ;
assign n7801 =  ( n7524 ) ? ( bv_8_148_n388 ) : ( n7800 ) ;
assign n7802 =  ( n7522 ) ? ( bv_8_152_n374 ) : ( n7801 ) ;
assign n7803 =  ( n7520 ) ? ( bv_8_176_n299 ) : ( n7802 ) ;
assign n7804 =  ( n7518 ) ? ( bv_8_133_n434 ) : ( n7803 ) ;
assign n7805 =  ( n7516 ) ? ( bv_8_187_n260 ) : ( n7804 ) ;
assign n7806 =  ( n7514 ) ? ( bv_8_197_n224 ) : ( n7805 ) ;
assign n7807 =  ( n7512 ) ? ( bv_8_79_n538 ) : ( n7806 ) ;
assign n7808 =  ( n7510 ) ? ( bv_8_237_n75 ) : ( n7807 ) ;
assign n7809 =  ( n7508 ) ? ( bv_8_134_n431 ) : ( n7808 ) ;
assign n7810 =  ( n7506 ) ? ( bv_8_154_n368 ) : ( n7809 ) ;
assign n7811 =  ( n7504 ) ? ( bv_8_102_n527 ) : ( n7810 ) ;
assign n7812 =  ( n7502 ) ? ( bv_8_17_n525 ) : ( n7811 ) ;
assign n7813 =  ( n7500 ) ? ( bv_8_138_n418 ) : ( n7812 ) ;
assign n7814 =  ( n7498 ) ? ( bv_8_233_n91 ) : ( n7813 ) ;
assign n7815 =  ( n7496 ) ? ( bv_8_4_n516 ) : ( n7814 ) ;
assign n7816 =  ( n7494 ) ? ( bv_8_254_n7 ) : ( n7815 ) ;
assign n7817 =  ( n7492 ) ? ( bv_8_160_n350 ) : ( n7816 ) ;
assign n7818 =  ( n7490 ) ? ( bv_8_120_n474 ) : ( n7817 ) ;
assign n7819 =  ( n7488 ) ? ( bv_8_37_n506 ) : ( n7818 ) ;
assign n7820 =  ( n7486 ) ? ( bv_8_75_n503 ) : ( n7819 ) ;
assign n7821 =  ( n7484 ) ? ( bv_8_162_n343 ) : ( n7820 ) ;
assign n7822 =  ( n7482 ) ? ( bv_8_93_n498 ) : ( n7821 ) ;
assign n7823 =  ( n7480 ) ? ( bv_8_128_n450 ) : ( n7822 ) ;
assign n7824 =  ( n7478 ) ? ( bv_8_5_n492 ) : ( n7823 ) ;
assign n7825 =  ( n7476 ) ? ( bv_8_63_n489 ) : ( n7824 ) ;
assign n7826 =  ( n7474 ) ? ( bv_8_33_n486 ) : ( n7825 ) ;
assign n7827 =  ( n7472 ) ? ( bv_8_112_n482 ) : ( n7826 ) ;
assign n7828 =  ( n7470 ) ? ( bv_8_241_n59 ) : ( n7827 ) ;
assign n7829 =  ( n7468 ) ? ( bv_8_99_n476 ) : ( n7828 ) ;
assign n7830 =  ( n7466 ) ? ( bv_8_119_n472 ) : ( n7829 ) ;
assign n7831 =  ( n7464 ) ? ( bv_8_175_n302 ) : ( n7830 ) ;
assign n7832 =  ( n7462 ) ? ( bv_8_66_n466 ) : ( n7831 ) ;
assign n7833 =  ( n7460 ) ? ( bv_8_32_n463 ) : ( n7832 ) ;
assign n7834 =  ( n7458 ) ? ( bv_8_229_n107 ) : ( n7833 ) ;
assign n7835 =  ( n7456 ) ? ( bv_8_253_n11 ) : ( n7834 ) ;
assign n7836 =  ( n7454 ) ? ( bv_8_191_n246 ) : ( n7835 ) ;
assign n7837 =  ( n7452 ) ? ( bv_8_129_n446 ) : ( n7836 ) ;
assign n7838 =  ( n7450 ) ? ( bv_8_24_n448 ) : ( n7837 ) ;
assign n7839 =  ( n7448 ) ? ( bv_8_38_n444 ) : ( n7838 ) ;
assign n7840 =  ( n7446 ) ? ( bv_8_195_n232 ) : ( n7839 ) ;
assign n7841 =  ( n7444 ) ? ( bv_8_190_n250 ) : ( n7840 ) ;
assign n7842 =  ( n7442 ) ? ( bv_8_53_n436 ) : ( n7841 ) ;
assign n7843 =  ( n7440 ) ? ( bv_8_136_n425 ) : ( n7842 ) ;
assign n7844 =  ( n7438 ) ? ( bv_8_46_n429 ) : ( n7843 ) ;
assign n7845 =  ( n7436 ) ? ( bv_8_147_n392 ) : ( n7844 ) ;
assign n7846 =  ( n7434 ) ? ( bv_8_85_n423 ) : ( n7845 ) ;
assign n7847 =  ( n7432 ) ? ( bv_8_252_n15 ) : ( n7846 ) ;
assign n7848 =  ( n7430 ) ? ( bv_8_122_n416 ) : ( n7847 ) ;
assign n7849 =  ( n7428 ) ? ( bv_8_200_n213 ) : ( n7848 ) ;
assign n7850 =  ( n7426 ) ? ( bv_8_186_n263 ) : ( n7849 ) ;
assign n7851 =  ( n7424 ) ? ( bv_8_50_n408 ) : ( n7850 ) ;
assign n7852 =  ( n7422 ) ? ( bv_8_230_n103 ) : ( n7851 ) ;
assign n7853 =  ( n7420 ) ? ( bv_8_192_n242 ) : ( n7852 ) ;
assign n7854 =  ( n7418 ) ? ( bv_8_25_n399 ) : ( n7853 ) ;
assign n7855 =  ( n7416 ) ? ( bv_8_158_n355 ) : ( n7854 ) ;
assign n7856 =  ( n7414 ) ? ( bv_8_163_n339 ) : ( n7855 ) ;
assign n7857 =  ( n7412 ) ? ( bv_8_68_n390 ) : ( n7856 ) ;
assign n7858 =  ( n7410 ) ? ( bv_8_84_n386 ) : ( n7857 ) ;
assign n7859 =  ( n7408 ) ? ( bv_8_59_n382 ) : ( n7858 ) ;
assign n7860 =  ( n7406 ) ? ( bv_8_11_n379 ) : ( n7859 ) ;
assign n7861 =  ( n7404 ) ? ( bv_8_140_n376 ) : ( n7860 ) ;
assign n7862 =  ( n7402 ) ? ( bv_8_199_n216 ) : ( n7861 ) ;
assign n7863 =  ( n7400 ) ? ( bv_8_107_n370 ) : ( n7862 ) ;
assign n7864 =  ( n7398 ) ? ( bv_8_40_n366 ) : ( n7863 ) ;
assign n7865 =  ( n7396 ) ? ( bv_8_167_n325 ) : ( n7864 ) ;
assign n7866 =  ( n7394 ) ? ( bv_8_188_n257 ) : ( n7865 ) ;
assign n7867 =  ( n7392 ) ? ( bv_8_22_n357 ) : ( n7866 ) ;
assign n7868 =  ( n7390 ) ? ( bv_8_173_n307 ) : ( n7867 ) ;
assign n7869 =  ( n7388 ) ? ( bv_8_219_n146 ) : ( n7868 ) ;
assign n7870 =  ( n7386 ) ? ( bv_8_100_n348 ) : ( n7869 ) ;
assign n7871 =  ( n7384 ) ? ( bv_8_116_n345 ) : ( n7870 ) ;
assign n7872 =  ( n7382 ) ? ( bv_8_20_n341 ) : ( n7871 ) ;
assign n7873 =  ( n7380 ) ? ( bv_8_146_n337 ) : ( n7872 ) ;
assign n7874 =  ( n7378 ) ? ( bv_8_12_n333 ) : ( n7873 ) ;
assign n7875 =  ( n7376 ) ? ( bv_8_72_n330 ) : ( n7874 ) ;
assign n7876 =  ( n7374 ) ? ( bv_8_184_n270 ) : ( n7875 ) ;
assign n7877 =  ( n7372 ) ? ( bv_8_159_n323 ) : ( n7876 ) ;
assign n7878 =  ( n7370 ) ? ( bv_8_189_n254 ) : ( n7877 ) ;
assign n7879 =  ( n7368 ) ? ( bv_8_67_n318 ) : ( n7878 ) ;
assign n7880 =  ( n7366 ) ? ( bv_8_196_n228 ) : ( n7879 ) ;
assign n7881 =  ( n7364 ) ? ( bv_8_57_n312 ) : ( n7880 ) ;
assign n7882 =  ( n7362 ) ? ( bv_8_49_n309 ) : ( n7881 ) ;
assign n7883 =  ( n7360 ) ? ( bv_8_211_n175 ) : ( n7882 ) ;
assign n7884 =  ( n7358 ) ? ( bv_8_242_n55 ) : ( n7883 ) ;
assign n7885 =  ( n7356 ) ? ( bv_8_213_n167 ) : ( n7884 ) ;
assign n7886 =  ( n7354 ) ? ( bv_8_139_n297 ) : ( n7885 ) ;
assign n7887 =  ( n7352 ) ? ( bv_8_110_n294 ) : ( n7886 ) ;
assign n7888 =  ( n7350 ) ? ( bv_8_218_n150 ) : ( n7887 ) ;
assign n7889 =  ( n7348 ) ? ( bv_8_1_n287 ) : ( n7888 ) ;
assign n7890 =  ( n7346 ) ? ( bv_8_177_n283 ) : ( n7889 ) ;
assign n7891 =  ( n7344 ) ? ( bv_8_156_n279 ) : ( n7890 ) ;
assign n7892 =  ( n7342 ) ? ( bv_8_73_n275 ) : ( n7891 ) ;
assign n7893 =  ( n7340 ) ? ( bv_8_216_n157 ) : ( n7892 ) ;
assign n7894 =  ( n7338 ) ? ( bv_8_172_n268 ) : ( n7893 ) ;
assign n7895 =  ( n7336 ) ? ( bv_8_243_n51 ) : ( n7894 ) ;
assign n7896 =  ( n7334 ) ? ( bv_8_207_n188 ) : ( n7895 ) ;
assign n7897 =  ( n7332 ) ? ( bv_8_202_n207 ) : ( n7896 ) ;
assign n7898 =  ( n7330 ) ? ( bv_8_244_n47 ) : ( n7897 ) ;
assign n7899 =  ( n7328 ) ? ( bv_8_71_n252 ) : ( n7898 ) ;
assign n7900 =  ( n7326 ) ? ( bv_8_16_n248 ) : ( n7899 ) ;
assign n7901 =  ( n7324 ) ? ( bv_8_111_n244 ) : ( n7900 ) ;
assign n7902 =  ( n7322 ) ? ( bv_8_240_n63 ) : ( n7901 ) ;
assign n7903 =  ( n7320 ) ? ( bv_8_74_n237 ) : ( n7902 ) ;
assign n7904 =  ( n7318 ) ? ( bv_8_92_n234 ) : ( n7903 ) ;
assign n7905 =  ( n7316 ) ? ( bv_8_56_n230 ) : ( n7904 ) ;
assign n7906 =  ( n7314 ) ? ( bv_8_87_n226 ) : ( n7905 ) ;
assign n7907 =  ( n7312 ) ? ( bv_8_115_n222 ) : ( n7906 ) ;
assign n7908 =  ( n7310 ) ? ( bv_8_151_n218 ) : ( n7907 ) ;
assign n7909 =  ( n7308 ) ? ( bv_8_203_n203 ) : ( n7908 ) ;
assign n7910 =  ( n7306 ) ? ( bv_8_161_n211 ) : ( n7909 ) ;
assign n7911 =  ( n7304 ) ? ( bv_8_232_n95 ) : ( n7910 ) ;
assign n7912 =  ( n7302 ) ? ( bv_8_62_n205 ) : ( n7911 ) ;
assign n7913 =  ( n7300 ) ? ( bv_8_150_n201 ) : ( n7912 ) ;
assign n7914 =  ( n7298 ) ? ( bv_8_97_n198 ) : ( n7913 ) ;
assign n7915 =  ( n7296 ) ? ( bv_8_13_n194 ) : ( n7914 ) ;
assign n7916 =  ( n7294 ) ? ( bv_8_15_n190 ) : ( n7915 ) ;
assign n7917 =  ( n7292 ) ? ( bv_8_224_n126 ) : ( n7916 ) ;
assign n7918 =  ( n7290 ) ? ( bv_8_124_n184 ) : ( n7917 ) ;
assign n7919 =  ( n7288 ) ? ( bv_8_113_n180 ) : ( n7918 ) ;
assign n7920 =  ( n7286 ) ? ( bv_8_204_n177 ) : ( n7919 ) ;
assign n7921 =  ( n7284 ) ? ( bv_8_144_n173 ) : ( n7920 ) ;
assign n7922 =  ( n7282 ) ? ( bv_8_6_n169 ) : ( n7921 ) ;
assign n7923 =  ( n7280 ) ? ( bv_8_247_n35 ) : ( n7922 ) ;
assign n7924 =  ( n7278 ) ? ( bv_8_28_n162 ) : ( n7923 ) ;
assign n7925 =  ( n7276 ) ? ( bv_8_194_n159 ) : ( n7924 ) ;
assign n7926 =  ( n7274 ) ? ( bv_8_106_n155 ) : ( n7925 ) ;
assign n7927 =  ( n7272 ) ? ( bv_8_174_n152 ) : ( n7926 ) ;
assign n7928 =  ( n7270 ) ? ( bv_8_105_n148 ) : ( n7927 ) ;
assign n7929 =  ( n7268 ) ? ( bv_8_23_n144 ) : ( n7928 ) ;
assign n7930 =  ( n7266 ) ? ( bv_8_153_n140 ) : ( n7929 ) ;
assign n7931 =  ( n7264 ) ? ( bv_8_58_n136 ) : ( n7930 ) ;
assign n7932 =  ( n7262 ) ? ( bv_8_39_n132 ) : ( n7931 ) ;
assign n7933 =  ( n7260 ) ? ( bv_8_217_n128 ) : ( n7932 ) ;
assign n7934 =  ( n7258 ) ? ( bv_8_235_n83 ) : ( n7933 ) ;
assign n7935 =  ( n7256 ) ? ( bv_8_43_n121 ) : ( n7934 ) ;
assign n7936 =  ( n7254 ) ? ( bv_8_34_n117 ) : ( n7935 ) ;
assign n7937 =  ( n7252 ) ? ( bv_8_210_n113 ) : ( n7936 ) ;
assign n7938 =  ( n7250 ) ? ( bv_8_169_n109 ) : ( n7937 ) ;
assign n7939 =  ( n7248 ) ? ( bv_8_7_n105 ) : ( n7938 ) ;
assign n7940 =  ( n7246 ) ? ( bv_8_51_n101 ) : ( n7939 ) ;
assign n7941 =  ( n7244 ) ? ( bv_8_45_n97 ) : ( n7940 ) ;
assign n7942 =  ( n7242 ) ? ( bv_8_60_n93 ) : ( n7941 ) ;
assign n7943 =  ( n7240 ) ? ( bv_8_21_n89 ) : ( n7942 ) ;
assign n7944 =  ( n7238 ) ? ( bv_8_201_n85 ) : ( n7943 ) ;
assign n7945 =  ( n7236 ) ? ( bv_8_135_n81 ) : ( n7944 ) ;
assign n7946 =  ( n7234 ) ? ( bv_8_170_n77 ) : ( n7945 ) ;
assign n7947 =  ( n7232 ) ? ( bv_8_80_n73 ) : ( n7946 ) ;
assign n7948 =  ( n7230 ) ? ( bv_8_165_n69 ) : ( n7947 ) ;
assign n7949 =  ( n7228 ) ? ( bv_8_3_n65 ) : ( n7948 ) ;
assign n7950 =  ( n7226 ) ? ( bv_8_89_n61 ) : ( n7949 ) ;
assign n7951 =  ( n7224 ) ? ( bv_8_9_n57 ) : ( n7950 ) ;
assign n7952 =  ( n7222 ) ? ( bv_8_26_n53 ) : ( n7951 ) ;
assign n7953 =  ( n7220 ) ? ( bv_8_101_n49 ) : ( n7952 ) ;
assign n7954 =  ( n7218 ) ? ( bv_8_215_n45 ) : ( n7953 ) ;
assign n7955 =  ( n7216 ) ? ( bv_8_132_n41 ) : ( n7954 ) ;
assign n7956 =  ( n7214 ) ? ( bv_8_208_n37 ) : ( n7955 ) ;
assign n7957 =  ( n7212 ) ? ( bv_8_130_n33 ) : ( n7956 ) ;
assign n7958 =  ( n7210 ) ? ( bv_8_41_n29 ) : ( n7957 ) ;
assign n7959 =  ( n7208 ) ? ( bv_8_90_n25 ) : ( n7958 ) ;
assign n7960 =  ( n7206 ) ? ( bv_8_30_n21 ) : ( n7959 ) ;
assign n7961 =  ( n7204 ) ? ( bv_8_123_n17 ) : ( n7960 ) ;
assign n7962 =  ( n7202 ) ? ( bv_8_168_n13 ) : ( n7961 ) ;
assign n7963 =  ( n7200 ) ? ( bv_8_109_n9 ) : ( n7962 ) ;
assign n7964 =  ( n7198 ) ? ( bv_8_44_n5 ) : ( n7963 ) ;
assign n7965 =  ( n7196 ) ^ ( n7964 )  ;
assign n7966 = state_in[55:48] ;
assign n7967 =  ( n7966 ) == ( bv_8_255_n3 )  ;
assign n7968 = state_in[55:48] ;
assign n7969 =  ( n7968 ) == ( bv_8_254_n7 )  ;
assign n7970 = state_in[55:48] ;
assign n7971 =  ( n7970 ) == ( bv_8_253_n11 )  ;
assign n7972 = state_in[55:48] ;
assign n7973 =  ( n7972 ) == ( bv_8_252_n15 )  ;
assign n7974 = state_in[55:48] ;
assign n7975 =  ( n7974 ) == ( bv_8_251_n19 )  ;
assign n7976 = state_in[55:48] ;
assign n7977 =  ( n7976 ) == ( bv_8_250_n23 )  ;
assign n7978 = state_in[55:48] ;
assign n7979 =  ( n7978 ) == ( bv_8_249_n27 )  ;
assign n7980 = state_in[55:48] ;
assign n7981 =  ( n7980 ) == ( bv_8_248_n31 )  ;
assign n7982 = state_in[55:48] ;
assign n7983 =  ( n7982 ) == ( bv_8_247_n35 )  ;
assign n7984 = state_in[55:48] ;
assign n7985 =  ( n7984 ) == ( bv_8_246_n39 )  ;
assign n7986 = state_in[55:48] ;
assign n7987 =  ( n7986 ) == ( bv_8_245_n43 )  ;
assign n7988 = state_in[55:48] ;
assign n7989 =  ( n7988 ) == ( bv_8_244_n47 )  ;
assign n7990 = state_in[55:48] ;
assign n7991 =  ( n7990 ) == ( bv_8_243_n51 )  ;
assign n7992 = state_in[55:48] ;
assign n7993 =  ( n7992 ) == ( bv_8_242_n55 )  ;
assign n7994 = state_in[55:48] ;
assign n7995 =  ( n7994 ) == ( bv_8_241_n59 )  ;
assign n7996 = state_in[55:48] ;
assign n7997 =  ( n7996 ) == ( bv_8_240_n63 )  ;
assign n7998 = state_in[55:48] ;
assign n7999 =  ( n7998 ) == ( bv_8_239_n67 )  ;
assign n8000 = state_in[55:48] ;
assign n8001 =  ( n8000 ) == ( bv_8_238_n71 )  ;
assign n8002 = state_in[55:48] ;
assign n8003 =  ( n8002 ) == ( bv_8_237_n75 )  ;
assign n8004 = state_in[55:48] ;
assign n8005 =  ( n8004 ) == ( bv_8_236_n79 )  ;
assign n8006 = state_in[55:48] ;
assign n8007 =  ( n8006 ) == ( bv_8_235_n83 )  ;
assign n8008 = state_in[55:48] ;
assign n8009 =  ( n8008 ) == ( bv_8_234_n87 )  ;
assign n8010 = state_in[55:48] ;
assign n8011 =  ( n8010 ) == ( bv_8_233_n91 )  ;
assign n8012 = state_in[55:48] ;
assign n8013 =  ( n8012 ) == ( bv_8_232_n95 )  ;
assign n8014 = state_in[55:48] ;
assign n8015 =  ( n8014 ) == ( bv_8_231_n99 )  ;
assign n8016 = state_in[55:48] ;
assign n8017 =  ( n8016 ) == ( bv_8_230_n103 )  ;
assign n8018 = state_in[55:48] ;
assign n8019 =  ( n8018 ) == ( bv_8_229_n107 )  ;
assign n8020 = state_in[55:48] ;
assign n8021 =  ( n8020 ) == ( bv_8_228_n111 )  ;
assign n8022 = state_in[55:48] ;
assign n8023 =  ( n8022 ) == ( bv_8_227_n115 )  ;
assign n8024 = state_in[55:48] ;
assign n8025 =  ( n8024 ) == ( bv_8_226_n119 )  ;
assign n8026 = state_in[55:48] ;
assign n8027 =  ( n8026 ) == ( bv_8_225_n123 )  ;
assign n8028 = state_in[55:48] ;
assign n8029 =  ( n8028 ) == ( bv_8_224_n126 )  ;
assign n8030 = state_in[55:48] ;
assign n8031 =  ( n8030 ) == ( bv_8_223_n130 )  ;
assign n8032 = state_in[55:48] ;
assign n8033 =  ( n8032 ) == ( bv_8_222_n134 )  ;
assign n8034 = state_in[55:48] ;
assign n8035 =  ( n8034 ) == ( bv_8_221_n138 )  ;
assign n8036 = state_in[55:48] ;
assign n8037 =  ( n8036 ) == ( bv_8_220_n142 )  ;
assign n8038 = state_in[55:48] ;
assign n8039 =  ( n8038 ) == ( bv_8_219_n146 )  ;
assign n8040 = state_in[55:48] ;
assign n8041 =  ( n8040 ) == ( bv_8_218_n150 )  ;
assign n8042 = state_in[55:48] ;
assign n8043 =  ( n8042 ) == ( bv_8_217_n128 )  ;
assign n8044 = state_in[55:48] ;
assign n8045 =  ( n8044 ) == ( bv_8_216_n157 )  ;
assign n8046 = state_in[55:48] ;
assign n8047 =  ( n8046 ) == ( bv_8_215_n45 )  ;
assign n8048 = state_in[55:48] ;
assign n8049 =  ( n8048 ) == ( bv_8_214_n164 )  ;
assign n8050 = state_in[55:48] ;
assign n8051 =  ( n8050 ) == ( bv_8_213_n167 )  ;
assign n8052 = state_in[55:48] ;
assign n8053 =  ( n8052 ) == ( bv_8_212_n171 )  ;
assign n8054 = state_in[55:48] ;
assign n8055 =  ( n8054 ) == ( bv_8_211_n175 )  ;
assign n8056 = state_in[55:48] ;
assign n8057 =  ( n8056 ) == ( bv_8_210_n113 )  ;
assign n8058 = state_in[55:48] ;
assign n8059 =  ( n8058 ) == ( bv_8_209_n182 )  ;
assign n8060 = state_in[55:48] ;
assign n8061 =  ( n8060 ) == ( bv_8_208_n37 )  ;
assign n8062 = state_in[55:48] ;
assign n8063 =  ( n8062 ) == ( bv_8_207_n188 )  ;
assign n8064 = state_in[55:48] ;
assign n8065 =  ( n8064 ) == ( bv_8_206_n192 )  ;
assign n8066 = state_in[55:48] ;
assign n8067 =  ( n8066 ) == ( bv_8_205_n196 )  ;
assign n8068 = state_in[55:48] ;
assign n8069 =  ( n8068 ) == ( bv_8_204_n177 )  ;
assign n8070 = state_in[55:48] ;
assign n8071 =  ( n8070 ) == ( bv_8_203_n203 )  ;
assign n8072 = state_in[55:48] ;
assign n8073 =  ( n8072 ) == ( bv_8_202_n207 )  ;
assign n8074 = state_in[55:48] ;
assign n8075 =  ( n8074 ) == ( bv_8_201_n85 )  ;
assign n8076 = state_in[55:48] ;
assign n8077 =  ( n8076 ) == ( bv_8_200_n213 )  ;
assign n8078 = state_in[55:48] ;
assign n8079 =  ( n8078 ) == ( bv_8_199_n216 )  ;
assign n8080 = state_in[55:48] ;
assign n8081 =  ( n8080 ) == ( bv_8_198_n220 )  ;
assign n8082 = state_in[55:48] ;
assign n8083 =  ( n8082 ) == ( bv_8_197_n224 )  ;
assign n8084 = state_in[55:48] ;
assign n8085 =  ( n8084 ) == ( bv_8_196_n228 )  ;
assign n8086 = state_in[55:48] ;
assign n8087 =  ( n8086 ) == ( bv_8_195_n232 )  ;
assign n8088 = state_in[55:48] ;
assign n8089 =  ( n8088 ) == ( bv_8_194_n159 )  ;
assign n8090 = state_in[55:48] ;
assign n8091 =  ( n8090 ) == ( bv_8_193_n239 )  ;
assign n8092 = state_in[55:48] ;
assign n8093 =  ( n8092 ) == ( bv_8_192_n242 )  ;
assign n8094 = state_in[55:48] ;
assign n8095 =  ( n8094 ) == ( bv_8_191_n246 )  ;
assign n8096 = state_in[55:48] ;
assign n8097 =  ( n8096 ) == ( bv_8_190_n250 )  ;
assign n8098 = state_in[55:48] ;
assign n8099 =  ( n8098 ) == ( bv_8_189_n254 )  ;
assign n8100 = state_in[55:48] ;
assign n8101 =  ( n8100 ) == ( bv_8_188_n257 )  ;
assign n8102 = state_in[55:48] ;
assign n8103 =  ( n8102 ) == ( bv_8_187_n260 )  ;
assign n8104 = state_in[55:48] ;
assign n8105 =  ( n8104 ) == ( bv_8_186_n263 )  ;
assign n8106 = state_in[55:48] ;
assign n8107 =  ( n8106 ) == ( bv_8_185_n266 )  ;
assign n8108 = state_in[55:48] ;
assign n8109 =  ( n8108 ) == ( bv_8_184_n270 )  ;
assign n8110 = state_in[55:48] ;
assign n8111 =  ( n8110 ) == ( bv_8_183_n273 )  ;
assign n8112 = state_in[55:48] ;
assign n8113 =  ( n8112 ) == ( bv_8_182_n277 )  ;
assign n8114 = state_in[55:48] ;
assign n8115 =  ( n8114 ) == ( bv_8_181_n281 )  ;
assign n8116 = state_in[55:48] ;
assign n8117 =  ( n8116 ) == ( bv_8_180_n285 )  ;
assign n8118 = state_in[55:48] ;
assign n8119 =  ( n8118 ) == ( bv_8_179_n289 )  ;
assign n8120 = state_in[55:48] ;
assign n8121 =  ( n8120 ) == ( bv_8_178_n292 )  ;
assign n8122 = state_in[55:48] ;
assign n8123 =  ( n8122 ) == ( bv_8_177_n283 )  ;
assign n8124 = state_in[55:48] ;
assign n8125 =  ( n8124 ) == ( bv_8_176_n299 )  ;
assign n8126 = state_in[55:48] ;
assign n8127 =  ( n8126 ) == ( bv_8_175_n302 )  ;
assign n8128 = state_in[55:48] ;
assign n8129 =  ( n8128 ) == ( bv_8_174_n152 )  ;
assign n8130 = state_in[55:48] ;
assign n8131 =  ( n8130 ) == ( bv_8_173_n307 )  ;
assign n8132 = state_in[55:48] ;
assign n8133 =  ( n8132 ) == ( bv_8_172_n268 )  ;
assign n8134 = state_in[55:48] ;
assign n8135 =  ( n8134 ) == ( bv_8_171_n314 )  ;
assign n8136 = state_in[55:48] ;
assign n8137 =  ( n8136 ) == ( bv_8_170_n77 )  ;
assign n8138 = state_in[55:48] ;
assign n8139 =  ( n8138 ) == ( bv_8_169_n109 )  ;
assign n8140 = state_in[55:48] ;
assign n8141 =  ( n8140 ) == ( bv_8_168_n13 )  ;
assign n8142 = state_in[55:48] ;
assign n8143 =  ( n8142 ) == ( bv_8_167_n325 )  ;
assign n8144 = state_in[55:48] ;
assign n8145 =  ( n8144 ) == ( bv_8_166_n328 )  ;
assign n8146 = state_in[55:48] ;
assign n8147 =  ( n8146 ) == ( bv_8_165_n69 )  ;
assign n8148 = state_in[55:48] ;
assign n8149 =  ( n8148 ) == ( bv_8_164_n335 )  ;
assign n8150 = state_in[55:48] ;
assign n8151 =  ( n8150 ) == ( bv_8_163_n339 )  ;
assign n8152 = state_in[55:48] ;
assign n8153 =  ( n8152 ) == ( bv_8_162_n343 )  ;
assign n8154 = state_in[55:48] ;
assign n8155 =  ( n8154 ) == ( bv_8_161_n211 )  ;
assign n8156 = state_in[55:48] ;
assign n8157 =  ( n8156 ) == ( bv_8_160_n350 )  ;
assign n8158 = state_in[55:48] ;
assign n8159 =  ( n8158 ) == ( bv_8_159_n323 )  ;
assign n8160 = state_in[55:48] ;
assign n8161 =  ( n8160 ) == ( bv_8_158_n355 )  ;
assign n8162 = state_in[55:48] ;
assign n8163 =  ( n8162 ) == ( bv_8_157_n359 )  ;
assign n8164 = state_in[55:48] ;
assign n8165 =  ( n8164 ) == ( bv_8_156_n279 )  ;
assign n8166 = state_in[55:48] ;
assign n8167 =  ( n8166 ) == ( bv_8_155_n364 )  ;
assign n8168 = state_in[55:48] ;
assign n8169 =  ( n8168 ) == ( bv_8_154_n368 )  ;
assign n8170 = state_in[55:48] ;
assign n8171 =  ( n8170 ) == ( bv_8_153_n140 )  ;
assign n8172 = state_in[55:48] ;
assign n8173 =  ( n8172 ) == ( bv_8_152_n374 )  ;
assign n8174 = state_in[55:48] ;
assign n8175 =  ( n8174 ) == ( bv_8_151_n218 )  ;
assign n8176 = state_in[55:48] ;
assign n8177 =  ( n8176 ) == ( bv_8_150_n201 )  ;
assign n8178 = state_in[55:48] ;
assign n8179 =  ( n8178 ) == ( bv_8_149_n384 )  ;
assign n8180 = state_in[55:48] ;
assign n8181 =  ( n8180 ) == ( bv_8_148_n388 )  ;
assign n8182 = state_in[55:48] ;
assign n8183 =  ( n8182 ) == ( bv_8_147_n392 )  ;
assign n8184 = state_in[55:48] ;
assign n8185 =  ( n8184 ) == ( bv_8_146_n337 )  ;
assign n8186 = state_in[55:48] ;
assign n8187 =  ( n8186 ) == ( bv_8_145_n397 )  ;
assign n8188 = state_in[55:48] ;
assign n8189 =  ( n8188 ) == ( bv_8_144_n173 )  ;
assign n8190 = state_in[55:48] ;
assign n8191 =  ( n8190 ) == ( bv_8_143_n403 )  ;
assign n8192 = state_in[55:48] ;
assign n8193 =  ( n8192 ) == ( bv_8_142_n406 )  ;
assign n8194 = state_in[55:48] ;
assign n8195 =  ( n8194 ) == ( bv_8_141_n410 )  ;
assign n8196 = state_in[55:48] ;
assign n8197 =  ( n8196 ) == ( bv_8_140_n376 )  ;
assign n8198 = state_in[55:48] ;
assign n8199 =  ( n8198 ) == ( bv_8_139_n297 )  ;
assign n8200 = state_in[55:48] ;
assign n8201 =  ( n8200 ) == ( bv_8_138_n418 )  ;
assign n8202 = state_in[55:48] ;
assign n8203 =  ( n8202 ) == ( bv_8_137_n421 )  ;
assign n8204 = state_in[55:48] ;
assign n8205 =  ( n8204 ) == ( bv_8_136_n425 )  ;
assign n8206 = state_in[55:48] ;
assign n8207 =  ( n8206 ) == ( bv_8_135_n81 )  ;
assign n8208 = state_in[55:48] ;
assign n8209 =  ( n8208 ) == ( bv_8_134_n431 )  ;
assign n8210 = state_in[55:48] ;
assign n8211 =  ( n8210 ) == ( bv_8_133_n434 )  ;
assign n8212 = state_in[55:48] ;
assign n8213 =  ( n8212 ) == ( bv_8_132_n41 )  ;
assign n8214 = state_in[55:48] ;
assign n8215 =  ( n8214 ) == ( bv_8_131_n440 )  ;
assign n8216 = state_in[55:48] ;
assign n8217 =  ( n8216 ) == ( bv_8_130_n33 )  ;
assign n8218 = state_in[55:48] ;
assign n8219 =  ( n8218 ) == ( bv_8_129_n446 )  ;
assign n8220 = state_in[55:48] ;
assign n8221 =  ( n8220 ) == ( bv_8_128_n450 )  ;
assign n8222 = state_in[55:48] ;
assign n8223 =  ( n8222 ) == ( bv_8_127_n453 )  ;
assign n8224 = state_in[55:48] ;
assign n8225 =  ( n8224 ) == ( bv_8_126_n456 )  ;
assign n8226 = state_in[55:48] ;
assign n8227 =  ( n8226 ) == ( bv_8_125_n459 )  ;
assign n8228 = state_in[55:48] ;
assign n8229 =  ( n8228 ) == ( bv_8_124_n184 )  ;
assign n8230 = state_in[55:48] ;
assign n8231 =  ( n8230 ) == ( bv_8_123_n17 )  ;
assign n8232 = state_in[55:48] ;
assign n8233 =  ( n8232 ) == ( bv_8_122_n416 )  ;
assign n8234 = state_in[55:48] ;
assign n8235 =  ( n8234 ) == ( bv_8_121_n470 )  ;
assign n8236 = state_in[55:48] ;
assign n8237 =  ( n8236 ) == ( bv_8_120_n474 )  ;
assign n8238 = state_in[55:48] ;
assign n8239 =  ( n8238 ) == ( bv_8_119_n472 )  ;
assign n8240 = state_in[55:48] ;
assign n8241 =  ( n8240 ) == ( bv_8_118_n480 )  ;
assign n8242 = state_in[55:48] ;
assign n8243 =  ( n8242 ) == ( bv_8_117_n484 )  ;
assign n8244 = state_in[55:48] ;
assign n8245 =  ( n8244 ) == ( bv_8_116_n345 )  ;
assign n8246 = state_in[55:48] ;
assign n8247 =  ( n8246 ) == ( bv_8_115_n222 )  ;
assign n8248 = state_in[55:48] ;
assign n8249 =  ( n8248 ) == ( bv_8_114_n494 )  ;
assign n8250 = state_in[55:48] ;
assign n8251 =  ( n8250 ) == ( bv_8_113_n180 )  ;
assign n8252 = state_in[55:48] ;
assign n8253 =  ( n8252 ) == ( bv_8_112_n482 )  ;
assign n8254 = state_in[55:48] ;
assign n8255 =  ( n8254 ) == ( bv_8_111_n244 )  ;
assign n8256 = state_in[55:48] ;
assign n8257 =  ( n8256 ) == ( bv_8_110_n294 )  ;
assign n8258 = state_in[55:48] ;
assign n8259 =  ( n8258 ) == ( bv_8_109_n9 )  ;
assign n8260 = state_in[55:48] ;
assign n8261 =  ( n8260 ) == ( bv_8_108_n510 )  ;
assign n8262 = state_in[55:48] ;
assign n8263 =  ( n8262 ) == ( bv_8_107_n370 )  ;
assign n8264 = state_in[55:48] ;
assign n8265 =  ( n8264 ) == ( bv_8_106_n155 )  ;
assign n8266 = state_in[55:48] ;
assign n8267 =  ( n8266 ) == ( bv_8_105_n148 )  ;
assign n8268 = state_in[55:48] ;
assign n8269 =  ( n8268 ) == ( bv_8_104_n520 )  ;
assign n8270 = state_in[55:48] ;
assign n8271 =  ( n8270 ) == ( bv_8_103_n523 )  ;
assign n8272 = state_in[55:48] ;
assign n8273 =  ( n8272 ) == ( bv_8_102_n527 )  ;
assign n8274 = state_in[55:48] ;
assign n8275 =  ( n8274 ) == ( bv_8_101_n49 )  ;
assign n8276 = state_in[55:48] ;
assign n8277 =  ( n8276 ) == ( bv_8_100_n348 )  ;
assign n8278 = state_in[55:48] ;
assign n8279 =  ( n8278 ) == ( bv_8_99_n476 )  ;
assign n8280 = state_in[55:48] ;
assign n8281 =  ( n8280 ) == ( bv_8_98_n536 )  ;
assign n8282 = state_in[55:48] ;
assign n8283 =  ( n8282 ) == ( bv_8_97_n198 )  ;
assign n8284 = state_in[55:48] ;
assign n8285 =  ( n8284 ) == ( bv_8_96_n542 )  ;
assign n8286 = state_in[55:48] ;
assign n8287 =  ( n8286 ) == ( bv_8_95_n545 )  ;
assign n8288 = state_in[55:48] ;
assign n8289 =  ( n8288 ) == ( bv_8_94_n548 )  ;
assign n8290 = state_in[55:48] ;
assign n8291 =  ( n8290 ) == ( bv_8_93_n498 )  ;
assign n8292 = state_in[55:48] ;
assign n8293 =  ( n8292 ) == ( bv_8_92_n234 )  ;
assign n8294 = state_in[55:48] ;
assign n8295 =  ( n8294 ) == ( bv_8_91_n555 )  ;
assign n8296 = state_in[55:48] ;
assign n8297 =  ( n8296 ) == ( bv_8_90_n25 )  ;
assign n8298 = state_in[55:48] ;
assign n8299 =  ( n8298 ) == ( bv_8_89_n61 )  ;
assign n8300 = state_in[55:48] ;
assign n8301 =  ( n8300 ) == ( bv_8_88_n562 )  ;
assign n8302 = state_in[55:48] ;
assign n8303 =  ( n8302 ) == ( bv_8_87_n226 )  ;
assign n8304 = state_in[55:48] ;
assign n8305 =  ( n8304 ) == ( bv_8_86_n567 )  ;
assign n8306 = state_in[55:48] ;
assign n8307 =  ( n8306 ) == ( bv_8_85_n423 )  ;
assign n8308 = state_in[55:48] ;
assign n8309 =  ( n8308 ) == ( bv_8_84_n386 )  ;
assign n8310 = state_in[55:48] ;
assign n8311 =  ( n8310 ) == ( bv_8_83_n575 )  ;
assign n8312 = state_in[55:48] ;
assign n8313 =  ( n8312 ) == ( bv_8_82_n578 )  ;
assign n8314 = state_in[55:48] ;
assign n8315 =  ( n8314 ) == ( bv_8_81_n582 )  ;
assign n8316 = state_in[55:48] ;
assign n8317 =  ( n8316 ) == ( bv_8_80_n73 )  ;
assign n8318 = state_in[55:48] ;
assign n8319 =  ( n8318 ) == ( bv_8_79_n538 )  ;
assign n8320 = state_in[55:48] ;
assign n8321 =  ( n8320 ) == ( bv_8_78_n590 )  ;
assign n8322 = state_in[55:48] ;
assign n8323 =  ( n8322 ) == ( bv_8_77_n593 )  ;
assign n8324 = state_in[55:48] ;
assign n8325 =  ( n8324 ) == ( bv_8_76_n596 )  ;
assign n8326 = state_in[55:48] ;
assign n8327 =  ( n8326 ) == ( bv_8_75_n503 )  ;
assign n8328 = state_in[55:48] ;
assign n8329 =  ( n8328 ) == ( bv_8_74_n237 )  ;
assign n8330 = state_in[55:48] ;
assign n8331 =  ( n8330 ) == ( bv_8_73_n275 )  ;
assign n8332 = state_in[55:48] ;
assign n8333 =  ( n8332 ) == ( bv_8_72_n330 )  ;
assign n8334 = state_in[55:48] ;
assign n8335 =  ( n8334 ) == ( bv_8_71_n252 )  ;
assign n8336 = state_in[55:48] ;
assign n8337 =  ( n8336 ) == ( bv_8_70_n609 )  ;
assign n8338 = state_in[55:48] ;
assign n8339 =  ( n8338 ) == ( bv_8_69_n612 )  ;
assign n8340 = state_in[55:48] ;
assign n8341 =  ( n8340 ) == ( bv_8_68_n390 )  ;
assign n8342 = state_in[55:48] ;
assign n8343 =  ( n8342 ) == ( bv_8_67_n318 )  ;
assign n8344 = state_in[55:48] ;
assign n8345 =  ( n8344 ) == ( bv_8_66_n466 )  ;
assign n8346 = state_in[55:48] ;
assign n8347 =  ( n8346 ) == ( bv_8_65_n623 )  ;
assign n8348 = state_in[55:48] ;
assign n8349 =  ( n8348 ) == ( bv_8_64_n573 )  ;
assign n8350 = state_in[55:48] ;
assign n8351 =  ( n8350 ) == ( bv_8_63_n489 )  ;
assign n8352 = state_in[55:48] ;
assign n8353 =  ( n8352 ) == ( bv_8_62_n205 )  ;
assign n8354 = state_in[55:48] ;
assign n8355 =  ( n8354 ) == ( bv_8_61_n634 )  ;
assign n8356 = state_in[55:48] ;
assign n8357 =  ( n8356 ) == ( bv_8_60_n93 )  ;
assign n8358 = state_in[55:48] ;
assign n8359 =  ( n8358 ) == ( bv_8_59_n382 )  ;
assign n8360 = state_in[55:48] ;
assign n8361 =  ( n8360 ) == ( bv_8_58_n136 )  ;
assign n8362 = state_in[55:48] ;
assign n8363 =  ( n8362 ) == ( bv_8_57_n312 )  ;
assign n8364 = state_in[55:48] ;
assign n8365 =  ( n8364 ) == ( bv_8_56_n230 )  ;
assign n8366 = state_in[55:48] ;
assign n8367 =  ( n8366 ) == ( bv_8_55_n650 )  ;
assign n8368 = state_in[55:48] ;
assign n8369 =  ( n8368 ) == ( bv_8_54_n616 )  ;
assign n8370 = state_in[55:48] ;
assign n8371 =  ( n8370 ) == ( bv_8_53_n436 )  ;
assign n8372 = state_in[55:48] ;
assign n8373 =  ( n8372 ) == ( bv_8_52_n619 )  ;
assign n8374 = state_in[55:48] ;
assign n8375 =  ( n8374 ) == ( bv_8_51_n101 )  ;
assign n8376 = state_in[55:48] ;
assign n8377 =  ( n8376 ) == ( bv_8_50_n408 )  ;
assign n8378 = state_in[55:48] ;
assign n8379 =  ( n8378 ) == ( bv_8_49_n309 )  ;
assign n8380 = state_in[55:48] ;
assign n8381 =  ( n8380 ) == ( bv_8_48_n660 )  ;
assign n8382 = state_in[55:48] ;
assign n8383 =  ( n8382 ) == ( bv_8_47_n652 )  ;
assign n8384 = state_in[55:48] ;
assign n8385 =  ( n8384 ) == ( bv_8_46_n429 )  ;
assign n8386 = state_in[55:48] ;
assign n8387 =  ( n8386 ) == ( bv_8_45_n97 )  ;
assign n8388 = state_in[55:48] ;
assign n8389 =  ( n8388 ) == ( bv_8_44_n5 )  ;
assign n8390 = state_in[55:48] ;
assign n8391 =  ( n8390 ) == ( bv_8_43_n121 )  ;
assign n8392 = state_in[55:48] ;
assign n8393 =  ( n8392 ) == ( bv_8_42_n672 )  ;
assign n8394 = state_in[55:48] ;
assign n8395 =  ( n8394 ) == ( bv_8_41_n29 )  ;
assign n8396 = state_in[55:48] ;
assign n8397 =  ( n8396 ) == ( bv_8_40_n366 )  ;
assign n8398 = state_in[55:48] ;
assign n8399 =  ( n8398 ) == ( bv_8_39_n132 )  ;
assign n8400 = state_in[55:48] ;
assign n8401 =  ( n8400 ) == ( bv_8_38_n444 )  ;
assign n8402 = state_in[55:48] ;
assign n8403 =  ( n8402 ) == ( bv_8_37_n506 )  ;
assign n8404 = state_in[55:48] ;
assign n8405 =  ( n8404 ) == ( bv_8_36_n645 )  ;
assign n8406 = state_in[55:48] ;
assign n8407 =  ( n8406 ) == ( bv_8_35_n696 )  ;
assign n8408 = state_in[55:48] ;
assign n8409 =  ( n8408 ) == ( bv_8_34_n117 )  ;
assign n8410 = state_in[55:48] ;
assign n8411 =  ( n8410 ) == ( bv_8_33_n486 )  ;
assign n8412 = state_in[55:48] ;
assign n8413 =  ( n8412 ) == ( bv_8_32_n463 )  ;
assign n8414 = state_in[55:48] ;
assign n8415 =  ( n8414 ) == ( bv_8_31_n705 )  ;
assign n8416 = state_in[55:48] ;
assign n8417 =  ( n8416 ) == ( bv_8_30_n21 )  ;
assign n8418 = state_in[55:48] ;
assign n8419 =  ( n8418 ) == ( bv_8_29_n625 )  ;
assign n8420 = state_in[55:48] ;
assign n8421 =  ( n8420 ) == ( bv_8_28_n162 )  ;
assign n8422 = state_in[55:48] ;
assign n8423 =  ( n8422 ) == ( bv_8_27_n642 )  ;
assign n8424 = state_in[55:48] ;
assign n8425 =  ( n8424 ) == ( bv_8_26_n53 )  ;
assign n8426 = state_in[55:48] ;
assign n8427 =  ( n8426 ) == ( bv_8_25_n399 )  ;
assign n8428 = state_in[55:48] ;
assign n8429 =  ( n8428 ) == ( bv_8_24_n448 )  ;
assign n8430 = state_in[55:48] ;
assign n8431 =  ( n8430 ) == ( bv_8_23_n144 )  ;
assign n8432 = state_in[55:48] ;
assign n8433 =  ( n8432 ) == ( bv_8_22_n357 )  ;
assign n8434 = state_in[55:48] ;
assign n8435 =  ( n8434 ) == ( bv_8_21_n89 )  ;
assign n8436 = state_in[55:48] ;
assign n8437 =  ( n8436 ) == ( bv_8_20_n341 )  ;
assign n8438 = state_in[55:48] ;
assign n8439 =  ( n8438 ) == ( bv_8_19_n588 )  ;
assign n8440 = state_in[55:48] ;
assign n8441 =  ( n8440 ) == ( bv_8_18_n628 )  ;
assign n8442 = state_in[55:48] ;
assign n8443 =  ( n8442 ) == ( bv_8_17_n525 )  ;
assign n8444 = state_in[55:48] ;
assign n8445 =  ( n8444 ) == ( bv_8_16_n248 )  ;
assign n8446 = state_in[55:48] ;
assign n8447 =  ( n8446 ) == ( bv_8_15_n190 )  ;
assign n8448 = state_in[55:48] ;
assign n8449 =  ( n8448 ) == ( bv_8_14_n648 )  ;
assign n8450 = state_in[55:48] ;
assign n8451 =  ( n8450 ) == ( bv_8_13_n194 )  ;
assign n8452 = state_in[55:48] ;
assign n8453 =  ( n8452 ) == ( bv_8_12_n333 )  ;
assign n8454 = state_in[55:48] ;
assign n8455 =  ( n8454 ) == ( bv_8_11_n379 )  ;
assign n8456 = state_in[55:48] ;
assign n8457 =  ( n8456 ) == ( bv_8_10_n655 )  ;
assign n8458 = state_in[55:48] ;
assign n8459 =  ( n8458 ) == ( bv_8_9_n57 )  ;
assign n8460 = state_in[55:48] ;
assign n8461 =  ( n8460 ) == ( bv_8_8_n669 )  ;
assign n8462 = state_in[55:48] ;
assign n8463 =  ( n8462 ) == ( bv_8_7_n105 )  ;
assign n8464 = state_in[55:48] ;
assign n8465 =  ( n8464 ) == ( bv_8_6_n169 )  ;
assign n8466 = state_in[55:48] ;
assign n8467 =  ( n8466 ) == ( bv_8_5_n492 )  ;
assign n8468 = state_in[55:48] ;
assign n8469 =  ( n8468 ) == ( bv_8_4_n516 )  ;
assign n8470 = state_in[55:48] ;
assign n8471 =  ( n8470 ) == ( bv_8_3_n65 )  ;
assign n8472 = state_in[55:48] ;
assign n8473 =  ( n8472 ) == ( bv_8_2_n751 )  ;
assign n8474 = state_in[55:48] ;
assign n8475 =  ( n8474 ) == ( bv_8_1_n287 )  ;
assign n8476 = state_in[55:48] ;
assign n8477 =  ( n8476 ) == ( bv_8_0_n580 )  ;
assign n8478 =  ( n8477 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n8479 =  ( n8475 ) ? ( bv_8_124_n184 ) : ( n8478 ) ;
assign n8480 =  ( n8473 ) ? ( bv_8_119_n472 ) : ( n8479 ) ;
assign n8481 =  ( n8471 ) ? ( bv_8_123_n17 ) : ( n8480 ) ;
assign n8482 =  ( n8469 ) ? ( bv_8_242_n55 ) : ( n8481 ) ;
assign n8483 =  ( n8467 ) ? ( bv_8_107_n370 ) : ( n8482 ) ;
assign n8484 =  ( n8465 ) ? ( bv_8_111_n244 ) : ( n8483 ) ;
assign n8485 =  ( n8463 ) ? ( bv_8_197_n224 ) : ( n8484 ) ;
assign n8486 =  ( n8461 ) ? ( bv_8_48_n660 ) : ( n8485 ) ;
assign n8487 =  ( n8459 ) ? ( bv_8_1_n287 ) : ( n8486 ) ;
assign n8488 =  ( n8457 ) ? ( bv_8_103_n523 ) : ( n8487 ) ;
assign n8489 =  ( n8455 ) ? ( bv_8_43_n121 ) : ( n8488 ) ;
assign n8490 =  ( n8453 ) ? ( bv_8_254_n7 ) : ( n8489 ) ;
assign n8491 =  ( n8451 ) ? ( bv_8_215_n45 ) : ( n8490 ) ;
assign n8492 =  ( n8449 ) ? ( bv_8_171_n314 ) : ( n8491 ) ;
assign n8493 =  ( n8447 ) ? ( bv_8_118_n480 ) : ( n8492 ) ;
assign n8494 =  ( n8445 ) ? ( bv_8_202_n207 ) : ( n8493 ) ;
assign n8495 =  ( n8443 ) ? ( bv_8_130_n33 ) : ( n8494 ) ;
assign n8496 =  ( n8441 ) ? ( bv_8_201_n85 ) : ( n8495 ) ;
assign n8497 =  ( n8439 ) ? ( bv_8_125_n459 ) : ( n8496 ) ;
assign n8498 =  ( n8437 ) ? ( bv_8_250_n23 ) : ( n8497 ) ;
assign n8499 =  ( n8435 ) ? ( bv_8_89_n61 ) : ( n8498 ) ;
assign n8500 =  ( n8433 ) ? ( bv_8_71_n252 ) : ( n8499 ) ;
assign n8501 =  ( n8431 ) ? ( bv_8_240_n63 ) : ( n8500 ) ;
assign n8502 =  ( n8429 ) ? ( bv_8_173_n307 ) : ( n8501 ) ;
assign n8503 =  ( n8427 ) ? ( bv_8_212_n171 ) : ( n8502 ) ;
assign n8504 =  ( n8425 ) ? ( bv_8_162_n343 ) : ( n8503 ) ;
assign n8505 =  ( n8423 ) ? ( bv_8_175_n302 ) : ( n8504 ) ;
assign n8506 =  ( n8421 ) ? ( bv_8_156_n279 ) : ( n8505 ) ;
assign n8507 =  ( n8419 ) ? ( bv_8_164_n335 ) : ( n8506 ) ;
assign n8508 =  ( n8417 ) ? ( bv_8_114_n494 ) : ( n8507 ) ;
assign n8509 =  ( n8415 ) ? ( bv_8_192_n242 ) : ( n8508 ) ;
assign n8510 =  ( n8413 ) ? ( bv_8_183_n273 ) : ( n8509 ) ;
assign n8511 =  ( n8411 ) ? ( bv_8_253_n11 ) : ( n8510 ) ;
assign n8512 =  ( n8409 ) ? ( bv_8_147_n392 ) : ( n8511 ) ;
assign n8513 =  ( n8407 ) ? ( bv_8_38_n444 ) : ( n8512 ) ;
assign n8514 =  ( n8405 ) ? ( bv_8_54_n616 ) : ( n8513 ) ;
assign n8515 =  ( n8403 ) ? ( bv_8_63_n489 ) : ( n8514 ) ;
assign n8516 =  ( n8401 ) ? ( bv_8_247_n35 ) : ( n8515 ) ;
assign n8517 =  ( n8399 ) ? ( bv_8_204_n177 ) : ( n8516 ) ;
assign n8518 =  ( n8397 ) ? ( bv_8_52_n619 ) : ( n8517 ) ;
assign n8519 =  ( n8395 ) ? ( bv_8_165_n69 ) : ( n8518 ) ;
assign n8520 =  ( n8393 ) ? ( bv_8_229_n107 ) : ( n8519 ) ;
assign n8521 =  ( n8391 ) ? ( bv_8_241_n59 ) : ( n8520 ) ;
assign n8522 =  ( n8389 ) ? ( bv_8_113_n180 ) : ( n8521 ) ;
assign n8523 =  ( n8387 ) ? ( bv_8_216_n157 ) : ( n8522 ) ;
assign n8524 =  ( n8385 ) ? ( bv_8_49_n309 ) : ( n8523 ) ;
assign n8525 =  ( n8383 ) ? ( bv_8_21_n89 ) : ( n8524 ) ;
assign n8526 =  ( n8381 ) ? ( bv_8_4_n516 ) : ( n8525 ) ;
assign n8527 =  ( n8379 ) ? ( bv_8_199_n216 ) : ( n8526 ) ;
assign n8528 =  ( n8377 ) ? ( bv_8_35_n696 ) : ( n8527 ) ;
assign n8529 =  ( n8375 ) ? ( bv_8_195_n232 ) : ( n8528 ) ;
assign n8530 =  ( n8373 ) ? ( bv_8_24_n448 ) : ( n8529 ) ;
assign n8531 =  ( n8371 ) ? ( bv_8_150_n201 ) : ( n8530 ) ;
assign n8532 =  ( n8369 ) ? ( bv_8_5_n492 ) : ( n8531 ) ;
assign n8533 =  ( n8367 ) ? ( bv_8_154_n368 ) : ( n8532 ) ;
assign n8534 =  ( n8365 ) ? ( bv_8_7_n105 ) : ( n8533 ) ;
assign n8535 =  ( n8363 ) ? ( bv_8_18_n628 ) : ( n8534 ) ;
assign n8536 =  ( n8361 ) ? ( bv_8_128_n450 ) : ( n8535 ) ;
assign n8537 =  ( n8359 ) ? ( bv_8_226_n119 ) : ( n8536 ) ;
assign n8538 =  ( n8357 ) ? ( bv_8_235_n83 ) : ( n8537 ) ;
assign n8539 =  ( n8355 ) ? ( bv_8_39_n132 ) : ( n8538 ) ;
assign n8540 =  ( n8353 ) ? ( bv_8_178_n292 ) : ( n8539 ) ;
assign n8541 =  ( n8351 ) ? ( bv_8_117_n484 ) : ( n8540 ) ;
assign n8542 =  ( n8349 ) ? ( bv_8_9_n57 ) : ( n8541 ) ;
assign n8543 =  ( n8347 ) ? ( bv_8_131_n440 ) : ( n8542 ) ;
assign n8544 =  ( n8345 ) ? ( bv_8_44_n5 ) : ( n8543 ) ;
assign n8545 =  ( n8343 ) ? ( bv_8_26_n53 ) : ( n8544 ) ;
assign n8546 =  ( n8341 ) ? ( bv_8_27_n642 ) : ( n8545 ) ;
assign n8547 =  ( n8339 ) ? ( bv_8_110_n294 ) : ( n8546 ) ;
assign n8548 =  ( n8337 ) ? ( bv_8_90_n25 ) : ( n8547 ) ;
assign n8549 =  ( n8335 ) ? ( bv_8_160_n350 ) : ( n8548 ) ;
assign n8550 =  ( n8333 ) ? ( bv_8_82_n578 ) : ( n8549 ) ;
assign n8551 =  ( n8331 ) ? ( bv_8_59_n382 ) : ( n8550 ) ;
assign n8552 =  ( n8329 ) ? ( bv_8_214_n164 ) : ( n8551 ) ;
assign n8553 =  ( n8327 ) ? ( bv_8_179_n289 ) : ( n8552 ) ;
assign n8554 =  ( n8325 ) ? ( bv_8_41_n29 ) : ( n8553 ) ;
assign n8555 =  ( n8323 ) ? ( bv_8_227_n115 ) : ( n8554 ) ;
assign n8556 =  ( n8321 ) ? ( bv_8_47_n652 ) : ( n8555 ) ;
assign n8557 =  ( n8319 ) ? ( bv_8_132_n41 ) : ( n8556 ) ;
assign n8558 =  ( n8317 ) ? ( bv_8_83_n575 ) : ( n8557 ) ;
assign n8559 =  ( n8315 ) ? ( bv_8_209_n182 ) : ( n8558 ) ;
assign n8560 =  ( n8313 ) ? ( bv_8_0_n580 ) : ( n8559 ) ;
assign n8561 =  ( n8311 ) ? ( bv_8_237_n75 ) : ( n8560 ) ;
assign n8562 =  ( n8309 ) ? ( bv_8_32_n463 ) : ( n8561 ) ;
assign n8563 =  ( n8307 ) ? ( bv_8_252_n15 ) : ( n8562 ) ;
assign n8564 =  ( n8305 ) ? ( bv_8_177_n283 ) : ( n8563 ) ;
assign n8565 =  ( n8303 ) ? ( bv_8_91_n555 ) : ( n8564 ) ;
assign n8566 =  ( n8301 ) ? ( bv_8_106_n155 ) : ( n8565 ) ;
assign n8567 =  ( n8299 ) ? ( bv_8_203_n203 ) : ( n8566 ) ;
assign n8568 =  ( n8297 ) ? ( bv_8_190_n250 ) : ( n8567 ) ;
assign n8569 =  ( n8295 ) ? ( bv_8_57_n312 ) : ( n8568 ) ;
assign n8570 =  ( n8293 ) ? ( bv_8_74_n237 ) : ( n8569 ) ;
assign n8571 =  ( n8291 ) ? ( bv_8_76_n596 ) : ( n8570 ) ;
assign n8572 =  ( n8289 ) ? ( bv_8_88_n562 ) : ( n8571 ) ;
assign n8573 =  ( n8287 ) ? ( bv_8_207_n188 ) : ( n8572 ) ;
assign n8574 =  ( n8285 ) ? ( bv_8_208_n37 ) : ( n8573 ) ;
assign n8575 =  ( n8283 ) ? ( bv_8_239_n67 ) : ( n8574 ) ;
assign n8576 =  ( n8281 ) ? ( bv_8_170_n77 ) : ( n8575 ) ;
assign n8577 =  ( n8279 ) ? ( bv_8_251_n19 ) : ( n8576 ) ;
assign n8578 =  ( n8277 ) ? ( bv_8_67_n318 ) : ( n8577 ) ;
assign n8579 =  ( n8275 ) ? ( bv_8_77_n593 ) : ( n8578 ) ;
assign n8580 =  ( n8273 ) ? ( bv_8_51_n101 ) : ( n8579 ) ;
assign n8581 =  ( n8271 ) ? ( bv_8_133_n434 ) : ( n8580 ) ;
assign n8582 =  ( n8269 ) ? ( bv_8_69_n612 ) : ( n8581 ) ;
assign n8583 =  ( n8267 ) ? ( bv_8_249_n27 ) : ( n8582 ) ;
assign n8584 =  ( n8265 ) ? ( bv_8_2_n751 ) : ( n8583 ) ;
assign n8585 =  ( n8263 ) ? ( bv_8_127_n453 ) : ( n8584 ) ;
assign n8586 =  ( n8261 ) ? ( bv_8_80_n73 ) : ( n8585 ) ;
assign n8587 =  ( n8259 ) ? ( bv_8_60_n93 ) : ( n8586 ) ;
assign n8588 =  ( n8257 ) ? ( bv_8_159_n323 ) : ( n8587 ) ;
assign n8589 =  ( n8255 ) ? ( bv_8_168_n13 ) : ( n8588 ) ;
assign n8590 =  ( n8253 ) ? ( bv_8_81_n582 ) : ( n8589 ) ;
assign n8591 =  ( n8251 ) ? ( bv_8_163_n339 ) : ( n8590 ) ;
assign n8592 =  ( n8249 ) ? ( bv_8_64_n573 ) : ( n8591 ) ;
assign n8593 =  ( n8247 ) ? ( bv_8_143_n403 ) : ( n8592 ) ;
assign n8594 =  ( n8245 ) ? ( bv_8_146_n337 ) : ( n8593 ) ;
assign n8595 =  ( n8243 ) ? ( bv_8_157_n359 ) : ( n8594 ) ;
assign n8596 =  ( n8241 ) ? ( bv_8_56_n230 ) : ( n8595 ) ;
assign n8597 =  ( n8239 ) ? ( bv_8_245_n43 ) : ( n8596 ) ;
assign n8598 =  ( n8237 ) ? ( bv_8_188_n257 ) : ( n8597 ) ;
assign n8599 =  ( n8235 ) ? ( bv_8_182_n277 ) : ( n8598 ) ;
assign n8600 =  ( n8233 ) ? ( bv_8_218_n150 ) : ( n8599 ) ;
assign n8601 =  ( n8231 ) ? ( bv_8_33_n486 ) : ( n8600 ) ;
assign n8602 =  ( n8229 ) ? ( bv_8_16_n248 ) : ( n8601 ) ;
assign n8603 =  ( n8227 ) ? ( bv_8_255_n3 ) : ( n8602 ) ;
assign n8604 =  ( n8225 ) ? ( bv_8_243_n51 ) : ( n8603 ) ;
assign n8605 =  ( n8223 ) ? ( bv_8_210_n113 ) : ( n8604 ) ;
assign n8606 =  ( n8221 ) ? ( bv_8_205_n196 ) : ( n8605 ) ;
assign n8607 =  ( n8219 ) ? ( bv_8_12_n333 ) : ( n8606 ) ;
assign n8608 =  ( n8217 ) ? ( bv_8_19_n588 ) : ( n8607 ) ;
assign n8609 =  ( n8215 ) ? ( bv_8_236_n79 ) : ( n8608 ) ;
assign n8610 =  ( n8213 ) ? ( bv_8_95_n545 ) : ( n8609 ) ;
assign n8611 =  ( n8211 ) ? ( bv_8_151_n218 ) : ( n8610 ) ;
assign n8612 =  ( n8209 ) ? ( bv_8_68_n390 ) : ( n8611 ) ;
assign n8613 =  ( n8207 ) ? ( bv_8_23_n144 ) : ( n8612 ) ;
assign n8614 =  ( n8205 ) ? ( bv_8_196_n228 ) : ( n8613 ) ;
assign n8615 =  ( n8203 ) ? ( bv_8_167_n325 ) : ( n8614 ) ;
assign n8616 =  ( n8201 ) ? ( bv_8_126_n456 ) : ( n8615 ) ;
assign n8617 =  ( n8199 ) ? ( bv_8_61_n634 ) : ( n8616 ) ;
assign n8618 =  ( n8197 ) ? ( bv_8_100_n348 ) : ( n8617 ) ;
assign n8619 =  ( n8195 ) ? ( bv_8_93_n498 ) : ( n8618 ) ;
assign n8620 =  ( n8193 ) ? ( bv_8_25_n399 ) : ( n8619 ) ;
assign n8621 =  ( n8191 ) ? ( bv_8_115_n222 ) : ( n8620 ) ;
assign n8622 =  ( n8189 ) ? ( bv_8_96_n542 ) : ( n8621 ) ;
assign n8623 =  ( n8187 ) ? ( bv_8_129_n446 ) : ( n8622 ) ;
assign n8624 =  ( n8185 ) ? ( bv_8_79_n538 ) : ( n8623 ) ;
assign n8625 =  ( n8183 ) ? ( bv_8_220_n142 ) : ( n8624 ) ;
assign n8626 =  ( n8181 ) ? ( bv_8_34_n117 ) : ( n8625 ) ;
assign n8627 =  ( n8179 ) ? ( bv_8_42_n672 ) : ( n8626 ) ;
assign n8628 =  ( n8177 ) ? ( bv_8_144_n173 ) : ( n8627 ) ;
assign n8629 =  ( n8175 ) ? ( bv_8_136_n425 ) : ( n8628 ) ;
assign n8630 =  ( n8173 ) ? ( bv_8_70_n609 ) : ( n8629 ) ;
assign n8631 =  ( n8171 ) ? ( bv_8_238_n71 ) : ( n8630 ) ;
assign n8632 =  ( n8169 ) ? ( bv_8_184_n270 ) : ( n8631 ) ;
assign n8633 =  ( n8167 ) ? ( bv_8_20_n341 ) : ( n8632 ) ;
assign n8634 =  ( n8165 ) ? ( bv_8_222_n134 ) : ( n8633 ) ;
assign n8635 =  ( n8163 ) ? ( bv_8_94_n548 ) : ( n8634 ) ;
assign n8636 =  ( n8161 ) ? ( bv_8_11_n379 ) : ( n8635 ) ;
assign n8637 =  ( n8159 ) ? ( bv_8_219_n146 ) : ( n8636 ) ;
assign n8638 =  ( n8157 ) ? ( bv_8_224_n126 ) : ( n8637 ) ;
assign n8639 =  ( n8155 ) ? ( bv_8_50_n408 ) : ( n8638 ) ;
assign n8640 =  ( n8153 ) ? ( bv_8_58_n136 ) : ( n8639 ) ;
assign n8641 =  ( n8151 ) ? ( bv_8_10_n655 ) : ( n8640 ) ;
assign n8642 =  ( n8149 ) ? ( bv_8_73_n275 ) : ( n8641 ) ;
assign n8643 =  ( n8147 ) ? ( bv_8_6_n169 ) : ( n8642 ) ;
assign n8644 =  ( n8145 ) ? ( bv_8_36_n645 ) : ( n8643 ) ;
assign n8645 =  ( n8143 ) ? ( bv_8_92_n234 ) : ( n8644 ) ;
assign n8646 =  ( n8141 ) ? ( bv_8_194_n159 ) : ( n8645 ) ;
assign n8647 =  ( n8139 ) ? ( bv_8_211_n175 ) : ( n8646 ) ;
assign n8648 =  ( n8137 ) ? ( bv_8_172_n268 ) : ( n8647 ) ;
assign n8649 =  ( n8135 ) ? ( bv_8_98_n536 ) : ( n8648 ) ;
assign n8650 =  ( n8133 ) ? ( bv_8_145_n397 ) : ( n8649 ) ;
assign n8651 =  ( n8131 ) ? ( bv_8_149_n384 ) : ( n8650 ) ;
assign n8652 =  ( n8129 ) ? ( bv_8_228_n111 ) : ( n8651 ) ;
assign n8653 =  ( n8127 ) ? ( bv_8_121_n470 ) : ( n8652 ) ;
assign n8654 =  ( n8125 ) ? ( bv_8_231_n99 ) : ( n8653 ) ;
assign n8655 =  ( n8123 ) ? ( bv_8_200_n213 ) : ( n8654 ) ;
assign n8656 =  ( n8121 ) ? ( bv_8_55_n650 ) : ( n8655 ) ;
assign n8657 =  ( n8119 ) ? ( bv_8_109_n9 ) : ( n8656 ) ;
assign n8658 =  ( n8117 ) ? ( bv_8_141_n410 ) : ( n8657 ) ;
assign n8659 =  ( n8115 ) ? ( bv_8_213_n167 ) : ( n8658 ) ;
assign n8660 =  ( n8113 ) ? ( bv_8_78_n590 ) : ( n8659 ) ;
assign n8661 =  ( n8111 ) ? ( bv_8_169_n109 ) : ( n8660 ) ;
assign n8662 =  ( n8109 ) ? ( bv_8_108_n510 ) : ( n8661 ) ;
assign n8663 =  ( n8107 ) ? ( bv_8_86_n567 ) : ( n8662 ) ;
assign n8664 =  ( n8105 ) ? ( bv_8_244_n47 ) : ( n8663 ) ;
assign n8665 =  ( n8103 ) ? ( bv_8_234_n87 ) : ( n8664 ) ;
assign n8666 =  ( n8101 ) ? ( bv_8_101_n49 ) : ( n8665 ) ;
assign n8667 =  ( n8099 ) ? ( bv_8_122_n416 ) : ( n8666 ) ;
assign n8668 =  ( n8097 ) ? ( bv_8_174_n152 ) : ( n8667 ) ;
assign n8669 =  ( n8095 ) ? ( bv_8_8_n669 ) : ( n8668 ) ;
assign n8670 =  ( n8093 ) ? ( bv_8_186_n263 ) : ( n8669 ) ;
assign n8671 =  ( n8091 ) ? ( bv_8_120_n474 ) : ( n8670 ) ;
assign n8672 =  ( n8089 ) ? ( bv_8_37_n506 ) : ( n8671 ) ;
assign n8673 =  ( n8087 ) ? ( bv_8_46_n429 ) : ( n8672 ) ;
assign n8674 =  ( n8085 ) ? ( bv_8_28_n162 ) : ( n8673 ) ;
assign n8675 =  ( n8083 ) ? ( bv_8_166_n328 ) : ( n8674 ) ;
assign n8676 =  ( n8081 ) ? ( bv_8_180_n285 ) : ( n8675 ) ;
assign n8677 =  ( n8079 ) ? ( bv_8_198_n220 ) : ( n8676 ) ;
assign n8678 =  ( n8077 ) ? ( bv_8_232_n95 ) : ( n8677 ) ;
assign n8679 =  ( n8075 ) ? ( bv_8_221_n138 ) : ( n8678 ) ;
assign n8680 =  ( n8073 ) ? ( bv_8_116_n345 ) : ( n8679 ) ;
assign n8681 =  ( n8071 ) ? ( bv_8_31_n705 ) : ( n8680 ) ;
assign n8682 =  ( n8069 ) ? ( bv_8_75_n503 ) : ( n8681 ) ;
assign n8683 =  ( n8067 ) ? ( bv_8_189_n254 ) : ( n8682 ) ;
assign n8684 =  ( n8065 ) ? ( bv_8_139_n297 ) : ( n8683 ) ;
assign n8685 =  ( n8063 ) ? ( bv_8_138_n418 ) : ( n8684 ) ;
assign n8686 =  ( n8061 ) ? ( bv_8_112_n482 ) : ( n8685 ) ;
assign n8687 =  ( n8059 ) ? ( bv_8_62_n205 ) : ( n8686 ) ;
assign n8688 =  ( n8057 ) ? ( bv_8_181_n281 ) : ( n8687 ) ;
assign n8689 =  ( n8055 ) ? ( bv_8_102_n527 ) : ( n8688 ) ;
assign n8690 =  ( n8053 ) ? ( bv_8_72_n330 ) : ( n8689 ) ;
assign n8691 =  ( n8051 ) ? ( bv_8_3_n65 ) : ( n8690 ) ;
assign n8692 =  ( n8049 ) ? ( bv_8_246_n39 ) : ( n8691 ) ;
assign n8693 =  ( n8047 ) ? ( bv_8_14_n648 ) : ( n8692 ) ;
assign n8694 =  ( n8045 ) ? ( bv_8_97_n198 ) : ( n8693 ) ;
assign n8695 =  ( n8043 ) ? ( bv_8_53_n436 ) : ( n8694 ) ;
assign n8696 =  ( n8041 ) ? ( bv_8_87_n226 ) : ( n8695 ) ;
assign n8697 =  ( n8039 ) ? ( bv_8_185_n266 ) : ( n8696 ) ;
assign n8698 =  ( n8037 ) ? ( bv_8_134_n431 ) : ( n8697 ) ;
assign n8699 =  ( n8035 ) ? ( bv_8_193_n239 ) : ( n8698 ) ;
assign n8700 =  ( n8033 ) ? ( bv_8_29_n625 ) : ( n8699 ) ;
assign n8701 =  ( n8031 ) ? ( bv_8_158_n355 ) : ( n8700 ) ;
assign n8702 =  ( n8029 ) ? ( bv_8_225_n123 ) : ( n8701 ) ;
assign n8703 =  ( n8027 ) ? ( bv_8_248_n31 ) : ( n8702 ) ;
assign n8704 =  ( n8025 ) ? ( bv_8_152_n374 ) : ( n8703 ) ;
assign n8705 =  ( n8023 ) ? ( bv_8_17_n525 ) : ( n8704 ) ;
assign n8706 =  ( n8021 ) ? ( bv_8_105_n148 ) : ( n8705 ) ;
assign n8707 =  ( n8019 ) ? ( bv_8_217_n128 ) : ( n8706 ) ;
assign n8708 =  ( n8017 ) ? ( bv_8_142_n406 ) : ( n8707 ) ;
assign n8709 =  ( n8015 ) ? ( bv_8_148_n388 ) : ( n8708 ) ;
assign n8710 =  ( n8013 ) ? ( bv_8_155_n364 ) : ( n8709 ) ;
assign n8711 =  ( n8011 ) ? ( bv_8_30_n21 ) : ( n8710 ) ;
assign n8712 =  ( n8009 ) ? ( bv_8_135_n81 ) : ( n8711 ) ;
assign n8713 =  ( n8007 ) ? ( bv_8_233_n91 ) : ( n8712 ) ;
assign n8714 =  ( n8005 ) ? ( bv_8_206_n192 ) : ( n8713 ) ;
assign n8715 =  ( n8003 ) ? ( bv_8_85_n423 ) : ( n8714 ) ;
assign n8716 =  ( n8001 ) ? ( bv_8_40_n366 ) : ( n8715 ) ;
assign n8717 =  ( n7999 ) ? ( bv_8_223_n130 ) : ( n8716 ) ;
assign n8718 =  ( n7997 ) ? ( bv_8_140_n376 ) : ( n8717 ) ;
assign n8719 =  ( n7995 ) ? ( bv_8_161_n211 ) : ( n8718 ) ;
assign n8720 =  ( n7993 ) ? ( bv_8_137_n421 ) : ( n8719 ) ;
assign n8721 =  ( n7991 ) ? ( bv_8_13_n194 ) : ( n8720 ) ;
assign n8722 =  ( n7989 ) ? ( bv_8_191_n246 ) : ( n8721 ) ;
assign n8723 =  ( n7987 ) ? ( bv_8_230_n103 ) : ( n8722 ) ;
assign n8724 =  ( n7985 ) ? ( bv_8_66_n466 ) : ( n8723 ) ;
assign n8725 =  ( n7983 ) ? ( bv_8_104_n520 ) : ( n8724 ) ;
assign n8726 =  ( n7981 ) ? ( bv_8_65_n623 ) : ( n8725 ) ;
assign n8727 =  ( n7979 ) ? ( bv_8_153_n140 ) : ( n8726 ) ;
assign n8728 =  ( n7977 ) ? ( bv_8_45_n97 ) : ( n8727 ) ;
assign n8729 =  ( n7975 ) ? ( bv_8_15_n190 ) : ( n8728 ) ;
assign n8730 =  ( n7973 ) ? ( bv_8_176_n299 ) : ( n8729 ) ;
assign n8731 =  ( n7971 ) ? ( bv_8_84_n386 ) : ( n8730 ) ;
assign n8732 =  ( n7969 ) ? ( bv_8_187_n260 ) : ( n8731 ) ;
assign n8733 =  ( n7967 ) ? ( bv_8_22_n357 ) : ( n8732 ) ;
assign n8734 =  ( n7965 ) ^ ( n8733 )  ;
assign n8735 = state_in[55:48] ;
assign n8736 =  ( n8735 ) == ( bv_8_255_n3 )  ;
assign n8737 = state_in[55:48] ;
assign n8738 =  ( n8737 ) == ( bv_8_254_n7 )  ;
assign n8739 = state_in[55:48] ;
assign n8740 =  ( n8739 ) == ( bv_8_253_n11 )  ;
assign n8741 = state_in[55:48] ;
assign n8742 =  ( n8741 ) == ( bv_8_252_n15 )  ;
assign n8743 = state_in[55:48] ;
assign n8744 =  ( n8743 ) == ( bv_8_251_n19 )  ;
assign n8745 = state_in[55:48] ;
assign n8746 =  ( n8745 ) == ( bv_8_250_n23 )  ;
assign n8747 = state_in[55:48] ;
assign n8748 =  ( n8747 ) == ( bv_8_249_n27 )  ;
assign n8749 = state_in[55:48] ;
assign n8750 =  ( n8749 ) == ( bv_8_248_n31 )  ;
assign n8751 = state_in[55:48] ;
assign n8752 =  ( n8751 ) == ( bv_8_247_n35 )  ;
assign n8753 = state_in[55:48] ;
assign n8754 =  ( n8753 ) == ( bv_8_246_n39 )  ;
assign n8755 = state_in[55:48] ;
assign n8756 =  ( n8755 ) == ( bv_8_245_n43 )  ;
assign n8757 = state_in[55:48] ;
assign n8758 =  ( n8757 ) == ( bv_8_244_n47 )  ;
assign n8759 = state_in[55:48] ;
assign n8760 =  ( n8759 ) == ( bv_8_243_n51 )  ;
assign n8761 = state_in[55:48] ;
assign n8762 =  ( n8761 ) == ( bv_8_242_n55 )  ;
assign n8763 = state_in[55:48] ;
assign n8764 =  ( n8763 ) == ( bv_8_241_n59 )  ;
assign n8765 = state_in[55:48] ;
assign n8766 =  ( n8765 ) == ( bv_8_240_n63 )  ;
assign n8767 = state_in[55:48] ;
assign n8768 =  ( n8767 ) == ( bv_8_239_n67 )  ;
assign n8769 = state_in[55:48] ;
assign n8770 =  ( n8769 ) == ( bv_8_238_n71 )  ;
assign n8771 = state_in[55:48] ;
assign n8772 =  ( n8771 ) == ( bv_8_237_n75 )  ;
assign n8773 = state_in[55:48] ;
assign n8774 =  ( n8773 ) == ( bv_8_236_n79 )  ;
assign n8775 = state_in[55:48] ;
assign n8776 =  ( n8775 ) == ( bv_8_235_n83 )  ;
assign n8777 = state_in[55:48] ;
assign n8778 =  ( n8777 ) == ( bv_8_234_n87 )  ;
assign n8779 = state_in[55:48] ;
assign n8780 =  ( n8779 ) == ( bv_8_233_n91 )  ;
assign n8781 = state_in[55:48] ;
assign n8782 =  ( n8781 ) == ( bv_8_232_n95 )  ;
assign n8783 = state_in[55:48] ;
assign n8784 =  ( n8783 ) == ( bv_8_231_n99 )  ;
assign n8785 = state_in[55:48] ;
assign n8786 =  ( n8785 ) == ( bv_8_230_n103 )  ;
assign n8787 = state_in[55:48] ;
assign n8788 =  ( n8787 ) == ( bv_8_229_n107 )  ;
assign n8789 = state_in[55:48] ;
assign n8790 =  ( n8789 ) == ( bv_8_228_n111 )  ;
assign n8791 = state_in[55:48] ;
assign n8792 =  ( n8791 ) == ( bv_8_227_n115 )  ;
assign n8793 = state_in[55:48] ;
assign n8794 =  ( n8793 ) == ( bv_8_226_n119 )  ;
assign n8795 = state_in[55:48] ;
assign n8796 =  ( n8795 ) == ( bv_8_225_n123 )  ;
assign n8797 = state_in[55:48] ;
assign n8798 =  ( n8797 ) == ( bv_8_224_n126 )  ;
assign n8799 = state_in[55:48] ;
assign n8800 =  ( n8799 ) == ( bv_8_223_n130 )  ;
assign n8801 = state_in[55:48] ;
assign n8802 =  ( n8801 ) == ( bv_8_222_n134 )  ;
assign n8803 = state_in[55:48] ;
assign n8804 =  ( n8803 ) == ( bv_8_221_n138 )  ;
assign n8805 = state_in[55:48] ;
assign n8806 =  ( n8805 ) == ( bv_8_220_n142 )  ;
assign n8807 = state_in[55:48] ;
assign n8808 =  ( n8807 ) == ( bv_8_219_n146 )  ;
assign n8809 = state_in[55:48] ;
assign n8810 =  ( n8809 ) == ( bv_8_218_n150 )  ;
assign n8811 = state_in[55:48] ;
assign n8812 =  ( n8811 ) == ( bv_8_217_n128 )  ;
assign n8813 = state_in[55:48] ;
assign n8814 =  ( n8813 ) == ( bv_8_216_n157 )  ;
assign n8815 = state_in[55:48] ;
assign n8816 =  ( n8815 ) == ( bv_8_215_n45 )  ;
assign n8817 = state_in[55:48] ;
assign n8818 =  ( n8817 ) == ( bv_8_214_n164 )  ;
assign n8819 = state_in[55:48] ;
assign n8820 =  ( n8819 ) == ( bv_8_213_n167 )  ;
assign n8821 = state_in[55:48] ;
assign n8822 =  ( n8821 ) == ( bv_8_212_n171 )  ;
assign n8823 = state_in[55:48] ;
assign n8824 =  ( n8823 ) == ( bv_8_211_n175 )  ;
assign n8825 = state_in[55:48] ;
assign n8826 =  ( n8825 ) == ( bv_8_210_n113 )  ;
assign n8827 = state_in[55:48] ;
assign n8828 =  ( n8827 ) == ( bv_8_209_n182 )  ;
assign n8829 = state_in[55:48] ;
assign n8830 =  ( n8829 ) == ( bv_8_208_n37 )  ;
assign n8831 = state_in[55:48] ;
assign n8832 =  ( n8831 ) == ( bv_8_207_n188 )  ;
assign n8833 = state_in[55:48] ;
assign n8834 =  ( n8833 ) == ( bv_8_206_n192 )  ;
assign n8835 = state_in[55:48] ;
assign n8836 =  ( n8835 ) == ( bv_8_205_n196 )  ;
assign n8837 = state_in[55:48] ;
assign n8838 =  ( n8837 ) == ( bv_8_204_n177 )  ;
assign n8839 = state_in[55:48] ;
assign n8840 =  ( n8839 ) == ( bv_8_203_n203 )  ;
assign n8841 = state_in[55:48] ;
assign n8842 =  ( n8841 ) == ( bv_8_202_n207 )  ;
assign n8843 = state_in[55:48] ;
assign n8844 =  ( n8843 ) == ( bv_8_201_n85 )  ;
assign n8845 = state_in[55:48] ;
assign n8846 =  ( n8845 ) == ( bv_8_200_n213 )  ;
assign n8847 = state_in[55:48] ;
assign n8848 =  ( n8847 ) == ( bv_8_199_n216 )  ;
assign n8849 = state_in[55:48] ;
assign n8850 =  ( n8849 ) == ( bv_8_198_n220 )  ;
assign n8851 = state_in[55:48] ;
assign n8852 =  ( n8851 ) == ( bv_8_197_n224 )  ;
assign n8853 = state_in[55:48] ;
assign n8854 =  ( n8853 ) == ( bv_8_196_n228 )  ;
assign n8855 = state_in[55:48] ;
assign n8856 =  ( n8855 ) == ( bv_8_195_n232 )  ;
assign n8857 = state_in[55:48] ;
assign n8858 =  ( n8857 ) == ( bv_8_194_n159 )  ;
assign n8859 = state_in[55:48] ;
assign n8860 =  ( n8859 ) == ( bv_8_193_n239 )  ;
assign n8861 = state_in[55:48] ;
assign n8862 =  ( n8861 ) == ( bv_8_192_n242 )  ;
assign n8863 = state_in[55:48] ;
assign n8864 =  ( n8863 ) == ( bv_8_191_n246 )  ;
assign n8865 = state_in[55:48] ;
assign n8866 =  ( n8865 ) == ( bv_8_190_n250 )  ;
assign n8867 = state_in[55:48] ;
assign n8868 =  ( n8867 ) == ( bv_8_189_n254 )  ;
assign n8869 = state_in[55:48] ;
assign n8870 =  ( n8869 ) == ( bv_8_188_n257 )  ;
assign n8871 = state_in[55:48] ;
assign n8872 =  ( n8871 ) == ( bv_8_187_n260 )  ;
assign n8873 = state_in[55:48] ;
assign n8874 =  ( n8873 ) == ( bv_8_186_n263 )  ;
assign n8875 = state_in[55:48] ;
assign n8876 =  ( n8875 ) == ( bv_8_185_n266 )  ;
assign n8877 = state_in[55:48] ;
assign n8878 =  ( n8877 ) == ( bv_8_184_n270 )  ;
assign n8879 = state_in[55:48] ;
assign n8880 =  ( n8879 ) == ( bv_8_183_n273 )  ;
assign n8881 = state_in[55:48] ;
assign n8882 =  ( n8881 ) == ( bv_8_182_n277 )  ;
assign n8883 = state_in[55:48] ;
assign n8884 =  ( n8883 ) == ( bv_8_181_n281 )  ;
assign n8885 = state_in[55:48] ;
assign n8886 =  ( n8885 ) == ( bv_8_180_n285 )  ;
assign n8887 = state_in[55:48] ;
assign n8888 =  ( n8887 ) == ( bv_8_179_n289 )  ;
assign n8889 = state_in[55:48] ;
assign n8890 =  ( n8889 ) == ( bv_8_178_n292 )  ;
assign n8891 = state_in[55:48] ;
assign n8892 =  ( n8891 ) == ( bv_8_177_n283 )  ;
assign n8893 = state_in[55:48] ;
assign n8894 =  ( n8893 ) == ( bv_8_176_n299 )  ;
assign n8895 = state_in[55:48] ;
assign n8896 =  ( n8895 ) == ( bv_8_175_n302 )  ;
assign n8897 = state_in[55:48] ;
assign n8898 =  ( n8897 ) == ( bv_8_174_n152 )  ;
assign n8899 = state_in[55:48] ;
assign n8900 =  ( n8899 ) == ( bv_8_173_n307 )  ;
assign n8901 = state_in[55:48] ;
assign n8902 =  ( n8901 ) == ( bv_8_172_n268 )  ;
assign n8903 = state_in[55:48] ;
assign n8904 =  ( n8903 ) == ( bv_8_171_n314 )  ;
assign n8905 = state_in[55:48] ;
assign n8906 =  ( n8905 ) == ( bv_8_170_n77 )  ;
assign n8907 = state_in[55:48] ;
assign n8908 =  ( n8907 ) == ( bv_8_169_n109 )  ;
assign n8909 = state_in[55:48] ;
assign n8910 =  ( n8909 ) == ( bv_8_168_n13 )  ;
assign n8911 = state_in[55:48] ;
assign n8912 =  ( n8911 ) == ( bv_8_167_n325 )  ;
assign n8913 = state_in[55:48] ;
assign n8914 =  ( n8913 ) == ( bv_8_166_n328 )  ;
assign n8915 = state_in[55:48] ;
assign n8916 =  ( n8915 ) == ( bv_8_165_n69 )  ;
assign n8917 = state_in[55:48] ;
assign n8918 =  ( n8917 ) == ( bv_8_164_n335 )  ;
assign n8919 = state_in[55:48] ;
assign n8920 =  ( n8919 ) == ( bv_8_163_n339 )  ;
assign n8921 = state_in[55:48] ;
assign n8922 =  ( n8921 ) == ( bv_8_162_n343 )  ;
assign n8923 = state_in[55:48] ;
assign n8924 =  ( n8923 ) == ( bv_8_161_n211 )  ;
assign n8925 = state_in[55:48] ;
assign n8926 =  ( n8925 ) == ( bv_8_160_n350 )  ;
assign n8927 = state_in[55:48] ;
assign n8928 =  ( n8927 ) == ( bv_8_159_n323 )  ;
assign n8929 = state_in[55:48] ;
assign n8930 =  ( n8929 ) == ( bv_8_158_n355 )  ;
assign n8931 = state_in[55:48] ;
assign n8932 =  ( n8931 ) == ( bv_8_157_n359 )  ;
assign n8933 = state_in[55:48] ;
assign n8934 =  ( n8933 ) == ( bv_8_156_n279 )  ;
assign n8935 = state_in[55:48] ;
assign n8936 =  ( n8935 ) == ( bv_8_155_n364 )  ;
assign n8937 = state_in[55:48] ;
assign n8938 =  ( n8937 ) == ( bv_8_154_n368 )  ;
assign n8939 = state_in[55:48] ;
assign n8940 =  ( n8939 ) == ( bv_8_153_n140 )  ;
assign n8941 = state_in[55:48] ;
assign n8942 =  ( n8941 ) == ( bv_8_152_n374 )  ;
assign n8943 = state_in[55:48] ;
assign n8944 =  ( n8943 ) == ( bv_8_151_n218 )  ;
assign n8945 = state_in[55:48] ;
assign n8946 =  ( n8945 ) == ( bv_8_150_n201 )  ;
assign n8947 = state_in[55:48] ;
assign n8948 =  ( n8947 ) == ( bv_8_149_n384 )  ;
assign n8949 = state_in[55:48] ;
assign n8950 =  ( n8949 ) == ( bv_8_148_n388 )  ;
assign n8951 = state_in[55:48] ;
assign n8952 =  ( n8951 ) == ( bv_8_147_n392 )  ;
assign n8953 = state_in[55:48] ;
assign n8954 =  ( n8953 ) == ( bv_8_146_n337 )  ;
assign n8955 = state_in[55:48] ;
assign n8956 =  ( n8955 ) == ( bv_8_145_n397 )  ;
assign n8957 = state_in[55:48] ;
assign n8958 =  ( n8957 ) == ( bv_8_144_n173 )  ;
assign n8959 = state_in[55:48] ;
assign n8960 =  ( n8959 ) == ( bv_8_143_n403 )  ;
assign n8961 = state_in[55:48] ;
assign n8962 =  ( n8961 ) == ( bv_8_142_n406 )  ;
assign n8963 = state_in[55:48] ;
assign n8964 =  ( n8963 ) == ( bv_8_141_n410 )  ;
assign n8965 = state_in[55:48] ;
assign n8966 =  ( n8965 ) == ( bv_8_140_n376 )  ;
assign n8967 = state_in[55:48] ;
assign n8968 =  ( n8967 ) == ( bv_8_139_n297 )  ;
assign n8969 = state_in[55:48] ;
assign n8970 =  ( n8969 ) == ( bv_8_138_n418 )  ;
assign n8971 = state_in[55:48] ;
assign n8972 =  ( n8971 ) == ( bv_8_137_n421 )  ;
assign n8973 = state_in[55:48] ;
assign n8974 =  ( n8973 ) == ( bv_8_136_n425 )  ;
assign n8975 = state_in[55:48] ;
assign n8976 =  ( n8975 ) == ( bv_8_135_n81 )  ;
assign n8977 = state_in[55:48] ;
assign n8978 =  ( n8977 ) == ( bv_8_134_n431 )  ;
assign n8979 = state_in[55:48] ;
assign n8980 =  ( n8979 ) == ( bv_8_133_n434 )  ;
assign n8981 = state_in[55:48] ;
assign n8982 =  ( n8981 ) == ( bv_8_132_n41 )  ;
assign n8983 = state_in[55:48] ;
assign n8984 =  ( n8983 ) == ( bv_8_131_n440 )  ;
assign n8985 = state_in[55:48] ;
assign n8986 =  ( n8985 ) == ( bv_8_130_n33 )  ;
assign n8987 = state_in[55:48] ;
assign n8988 =  ( n8987 ) == ( bv_8_129_n446 )  ;
assign n8989 = state_in[55:48] ;
assign n8990 =  ( n8989 ) == ( bv_8_128_n450 )  ;
assign n8991 = state_in[55:48] ;
assign n8992 =  ( n8991 ) == ( bv_8_127_n453 )  ;
assign n8993 = state_in[55:48] ;
assign n8994 =  ( n8993 ) == ( bv_8_126_n456 )  ;
assign n8995 = state_in[55:48] ;
assign n8996 =  ( n8995 ) == ( bv_8_125_n459 )  ;
assign n8997 = state_in[55:48] ;
assign n8998 =  ( n8997 ) == ( bv_8_124_n184 )  ;
assign n8999 = state_in[55:48] ;
assign n9000 =  ( n8999 ) == ( bv_8_123_n17 )  ;
assign n9001 = state_in[55:48] ;
assign n9002 =  ( n9001 ) == ( bv_8_122_n416 )  ;
assign n9003 = state_in[55:48] ;
assign n9004 =  ( n9003 ) == ( bv_8_121_n470 )  ;
assign n9005 = state_in[55:48] ;
assign n9006 =  ( n9005 ) == ( bv_8_120_n474 )  ;
assign n9007 = state_in[55:48] ;
assign n9008 =  ( n9007 ) == ( bv_8_119_n472 )  ;
assign n9009 = state_in[55:48] ;
assign n9010 =  ( n9009 ) == ( bv_8_118_n480 )  ;
assign n9011 = state_in[55:48] ;
assign n9012 =  ( n9011 ) == ( bv_8_117_n484 )  ;
assign n9013 = state_in[55:48] ;
assign n9014 =  ( n9013 ) == ( bv_8_116_n345 )  ;
assign n9015 = state_in[55:48] ;
assign n9016 =  ( n9015 ) == ( bv_8_115_n222 )  ;
assign n9017 = state_in[55:48] ;
assign n9018 =  ( n9017 ) == ( bv_8_114_n494 )  ;
assign n9019 = state_in[55:48] ;
assign n9020 =  ( n9019 ) == ( bv_8_113_n180 )  ;
assign n9021 = state_in[55:48] ;
assign n9022 =  ( n9021 ) == ( bv_8_112_n482 )  ;
assign n9023 = state_in[55:48] ;
assign n9024 =  ( n9023 ) == ( bv_8_111_n244 )  ;
assign n9025 = state_in[55:48] ;
assign n9026 =  ( n9025 ) == ( bv_8_110_n294 )  ;
assign n9027 = state_in[55:48] ;
assign n9028 =  ( n9027 ) == ( bv_8_109_n9 )  ;
assign n9029 = state_in[55:48] ;
assign n9030 =  ( n9029 ) == ( bv_8_108_n510 )  ;
assign n9031 = state_in[55:48] ;
assign n9032 =  ( n9031 ) == ( bv_8_107_n370 )  ;
assign n9033 = state_in[55:48] ;
assign n9034 =  ( n9033 ) == ( bv_8_106_n155 )  ;
assign n9035 = state_in[55:48] ;
assign n9036 =  ( n9035 ) == ( bv_8_105_n148 )  ;
assign n9037 = state_in[55:48] ;
assign n9038 =  ( n9037 ) == ( bv_8_104_n520 )  ;
assign n9039 = state_in[55:48] ;
assign n9040 =  ( n9039 ) == ( bv_8_103_n523 )  ;
assign n9041 = state_in[55:48] ;
assign n9042 =  ( n9041 ) == ( bv_8_102_n527 )  ;
assign n9043 = state_in[55:48] ;
assign n9044 =  ( n9043 ) == ( bv_8_101_n49 )  ;
assign n9045 = state_in[55:48] ;
assign n9046 =  ( n9045 ) == ( bv_8_100_n348 )  ;
assign n9047 = state_in[55:48] ;
assign n9048 =  ( n9047 ) == ( bv_8_99_n476 )  ;
assign n9049 = state_in[55:48] ;
assign n9050 =  ( n9049 ) == ( bv_8_98_n536 )  ;
assign n9051 = state_in[55:48] ;
assign n9052 =  ( n9051 ) == ( bv_8_97_n198 )  ;
assign n9053 = state_in[55:48] ;
assign n9054 =  ( n9053 ) == ( bv_8_96_n542 )  ;
assign n9055 = state_in[55:48] ;
assign n9056 =  ( n9055 ) == ( bv_8_95_n545 )  ;
assign n9057 = state_in[55:48] ;
assign n9058 =  ( n9057 ) == ( bv_8_94_n548 )  ;
assign n9059 = state_in[55:48] ;
assign n9060 =  ( n9059 ) == ( bv_8_93_n498 )  ;
assign n9061 = state_in[55:48] ;
assign n9062 =  ( n9061 ) == ( bv_8_92_n234 )  ;
assign n9063 = state_in[55:48] ;
assign n9064 =  ( n9063 ) == ( bv_8_91_n555 )  ;
assign n9065 = state_in[55:48] ;
assign n9066 =  ( n9065 ) == ( bv_8_90_n25 )  ;
assign n9067 = state_in[55:48] ;
assign n9068 =  ( n9067 ) == ( bv_8_89_n61 )  ;
assign n9069 = state_in[55:48] ;
assign n9070 =  ( n9069 ) == ( bv_8_88_n562 )  ;
assign n9071 = state_in[55:48] ;
assign n9072 =  ( n9071 ) == ( bv_8_87_n226 )  ;
assign n9073 = state_in[55:48] ;
assign n9074 =  ( n9073 ) == ( bv_8_86_n567 )  ;
assign n9075 = state_in[55:48] ;
assign n9076 =  ( n9075 ) == ( bv_8_85_n423 )  ;
assign n9077 = state_in[55:48] ;
assign n9078 =  ( n9077 ) == ( bv_8_84_n386 )  ;
assign n9079 = state_in[55:48] ;
assign n9080 =  ( n9079 ) == ( bv_8_83_n575 )  ;
assign n9081 = state_in[55:48] ;
assign n9082 =  ( n9081 ) == ( bv_8_82_n578 )  ;
assign n9083 = state_in[55:48] ;
assign n9084 =  ( n9083 ) == ( bv_8_81_n582 )  ;
assign n9085 = state_in[55:48] ;
assign n9086 =  ( n9085 ) == ( bv_8_80_n73 )  ;
assign n9087 = state_in[55:48] ;
assign n9088 =  ( n9087 ) == ( bv_8_79_n538 )  ;
assign n9089 = state_in[55:48] ;
assign n9090 =  ( n9089 ) == ( bv_8_78_n590 )  ;
assign n9091 = state_in[55:48] ;
assign n9092 =  ( n9091 ) == ( bv_8_77_n593 )  ;
assign n9093 = state_in[55:48] ;
assign n9094 =  ( n9093 ) == ( bv_8_76_n596 )  ;
assign n9095 = state_in[55:48] ;
assign n9096 =  ( n9095 ) == ( bv_8_75_n503 )  ;
assign n9097 = state_in[55:48] ;
assign n9098 =  ( n9097 ) == ( bv_8_74_n237 )  ;
assign n9099 = state_in[55:48] ;
assign n9100 =  ( n9099 ) == ( bv_8_73_n275 )  ;
assign n9101 = state_in[55:48] ;
assign n9102 =  ( n9101 ) == ( bv_8_72_n330 )  ;
assign n9103 = state_in[55:48] ;
assign n9104 =  ( n9103 ) == ( bv_8_71_n252 )  ;
assign n9105 = state_in[55:48] ;
assign n9106 =  ( n9105 ) == ( bv_8_70_n609 )  ;
assign n9107 = state_in[55:48] ;
assign n9108 =  ( n9107 ) == ( bv_8_69_n612 )  ;
assign n9109 = state_in[55:48] ;
assign n9110 =  ( n9109 ) == ( bv_8_68_n390 )  ;
assign n9111 = state_in[55:48] ;
assign n9112 =  ( n9111 ) == ( bv_8_67_n318 )  ;
assign n9113 = state_in[55:48] ;
assign n9114 =  ( n9113 ) == ( bv_8_66_n466 )  ;
assign n9115 = state_in[55:48] ;
assign n9116 =  ( n9115 ) == ( bv_8_65_n623 )  ;
assign n9117 = state_in[55:48] ;
assign n9118 =  ( n9117 ) == ( bv_8_64_n573 )  ;
assign n9119 = state_in[55:48] ;
assign n9120 =  ( n9119 ) == ( bv_8_63_n489 )  ;
assign n9121 = state_in[55:48] ;
assign n9122 =  ( n9121 ) == ( bv_8_62_n205 )  ;
assign n9123 = state_in[55:48] ;
assign n9124 =  ( n9123 ) == ( bv_8_61_n634 )  ;
assign n9125 = state_in[55:48] ;
assign n9126 =  ( n9125 ) == ( bv_8_60_n93 )  ;
assign n9127 = state_in[55:48] ;
assign n9128 =  ( n9127 ) == ( bv_8_59_n382 )  ;
assign n9129 = state_in[55:48] ;
assign n9130 =  ( n9129 ) == ( bv_8_58_n136 )  ;
assign n9131 = state_in[55:48] ;
assign n9132 =  ( n9131 ) == ( bv_8_57_n312 )  ;
assign n9133 = state_in[55:48] ;
assign n9134 =  ( n9133 ) == ( bv_8_56_n230 )  ;
assign n9135 = state_in[55:48] ;
assign n9136 =  ( n9135 ) == ( bv_8_55_n650 )  ;
assign n9137 = state_in[55:48] ;
assign n9138 =  ( n9137 ) == ( bv_8_54_n616 )  ;
assign n9139 = state_in[55:48] ;
assign n9140 =  ( n9139 ) == ( bv_8_53_n436 )  ;
assign n9141 = state_in[55:48] ;
assign n9142 =  ( n9141 ) == ( bv_8_52_n619 )  ;
assign n9143 = state_in[55:48] ;
assign n9144 =  ( n9143 ) == ( bv_8_51_n101 )  ;
assign n9145 = state_in[55:48] ;
assign n9146 =  ( n9145 ) == ( bv_8_50_n408 )  ;
assign n9147 = state_in[55:48] ;
assign n9148 =  ( n9147 ) == ( bv_8_49_n309 )  ;
assign n9149 = state_in[55:48] ;
assign n9150 =  ( n9149 ) == ( bv_8_48_n660 )  ;
assign n9151 = state_in[55:48] ;
assign n9152 =  ( n9151 ) == ( bv_8_47_n652 )  ;
assign n9153 = state_in[55:48] ;
assign n9154 =  ( n9153 ) == ( bv_8_46_n429 )  ;
assign n9155 = state_in[55:48] ;
assign n9156 =  ( n9155 ) == ( bv_8_45_n97 )  ;
assign n9157 = state_in[55:48] ;
assign n9158 =  ( n9157 ) == ( bv_8_44_n5 )  ;
assign n9159 = state_in[55:48] ;
assign n9160 =  ( n9159 ) == ( bv_8_43_n121 )  ;
assign n9161 = state_in[55:48] ;
assign n9162 =  ( n9161 ) == ( bv_8_42_n672 )  ;
assign n9163 = state_in[55:48] ;
assign n9164 =  ( n9163 ) == ( bv_8_41_n29 )  ;
assign n9165 = state_in[55:48] ;
assign n9166 =  ( n9165 ) == ( bv_8_40_n366 )  ;
assign n9167 = state_in[55:48] ;
assign n9168 =  ( n9167 ) == ( bv_8_39_n132 )  ;
assign n9169 = state_in[55:48] ;
assign n9170 =  ( n9169 ) == ( bv_8_38_n444 )  ;
assign n9171 = state_in[55:48] ;
assign n9172 =  ( n9171 ) == ( bv_8_37_n506 )  ;
assign n9173 = state_in[55:48] ;
assign n9174 =  ( n9173 ) == ( bv_8_36_n645 )  ;
assign n9175 = state_in[55:48] ;
assign n9176 =  ( n9175 ) == ( bv_8_35_n696 )  ;
assign n9177 = state_in[55:48] ;
assign n9178 =  ( n9177 ) == ( bv_8_34_n117 )  ;
assign n9179 = state_in[55:48] ;
assign n9180 =  ( n9179 ) == ( bv_8_33_n486 )  ;
assign n9181 = state_in[55:48] ;
assign n9182 =  ( n9181 ) == ( bv_8_32_n463 )  ;
assign n9183 = state_in[55:48] ;
assign n9184 =  ( n9183 ) == ( bv_8_31_n705 )  ;
assign n9185 = state_in[55:48] ;
assign n9186 =  ( n9185 ) == ( bv_8_30_n21 )  ;
assign n9187 = state_in[55:48] ;
assign n9188 =  ( n9187 ) == ( bv_8_29_n625 )  ;
assign n9189 = state_in[55:48] ;
assign n9190 =  ( n9189 ) == ( bv_8_28_n162 )  ;
assign n9191 = state_in[55:48] ;
assign n9192 =  ( n9191 ) == ( bv_8_27_n642 )  ;
assign n9193 = state_in[55:48] ;
assign n9194 =  ( n9193 ) == ( bv_8_26_n53 )  ;
assign n9195 = state_in[55:48] ;
assign n9196 =  ( n9195 ) == ( bv_8_25_n399 )  ;
assign n9197 = state_in[55:48] ;
assign n9198 =  ( n9197 ) == ( bv_8_24_n448 )  ;
assign n9199 = state_in[55:48] ;
assign n9200 =  ( n9199 ) == ( bv_8_23_n144 )  ;
assign n9201 = state_in[55:48] ;
assign n9202 =  ( n9201 ) == ( bv_8_22_n357 )  ;
assign n9203 = state_in[55:48] ;
assign n9204 =  ( n9203 ) == ( bv_8_21_n89 )  ;
assign n9205 = state_in[55:48] ;
assign n9206 =  ( n9205 ) == ( bv_8_20_n341 )  ;
assign n9207 = state_in[55:48] ;
assign n9208 =  ( n9207 ) == ( bv_8_19_n588 )  ;
assign n9209 = state_in[55:48] ;
assign n9210 =  ( n9209 ) == ( bv_8_18_n628 )  ;
assign n9211 = state_in[55:48] ;
assign n9212 =  ( n9211 ) == ( bv_8_17_n525 )  ;
assign n9213 = state_in[55:48] ;
assign n9214 =  ( n9213 ) == ( bv_8_16_n248 )  ;
assign n9215 = state_in[55:48] ;
assign n9216 =  ( n9215 ) == ( bv_8_15_n190 )  ;
assign n9217 = state_in[55:48] ;
assign n9218 =  ( n9217 ) == ( bv_8_14_n648 )  ;
assign n9219 = state_in[55:48] ;
assign n9220 =  ( n9219 ) == ( bv_8_13_n194 )  ;
assign n9221 = state_in[55:48] ;
assign n9222 =  ( n9221 ) == ( bv_8_12_n333 )  ;
assign n9223 = state_in[55:48] ;
assign n9224 =  ( n9223 ) == ( bv_8_11_n379 )  ;
assign n9225 = state_in[55:48] ;
assign n9226 =  ( n9225 ) == ( bv_8_10_n655 )  ;
assign n9227 = state_in[55:48] ;
assign n9228 =  ( n9227 ) == ( bv_8_9_n57 )  ;
assign n9229 = state_in[55:48] ;
assign n9230 =  ( n9229 ) == ( bv_8_8_n669 )  ;
assign n9231 = state_in[55:48] ;
assign n9232 =  ( n9231 ) == ( bv_8_7_n105 )  ;
assign n9233 = state_in[55:48] ;
assign n9234 =  ( n9233 ) == ( bv_8_6_n169 )  ;
assign n9235 = state_in[55:48] ;
assign n9236 =  ( n9235 ) == ( bv_8_5_n492 )  ;
assign n9237 = state_in[55:48] ;
assign n9238 =  ( n9237 ) == ( bv_8_4_n516 )  ;
assign n9239 = state_in[55:48] ;
assign n9240 =  ( n9239 ) == ( bv_8_3_n65 )  ;
assign n9241 = state_in[55:48] ;
assign n9242 =  ( n9241 ) == ( bv_8_2_n751 )  ;
assign n9243 = state_in[55:48] ;
assign n9244 =  ( n9243 ) == ( bv_8_1_n287 )  ;
assign n9245 = state_in[55:48] ;
assign n9246 =  ( n9245 ) == ( bv_8_0_n580 )  ;
assign n9247 =  ( n9246 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n9248 =  ( n9244 ) ? ( bv_8_248_n31 ) : ( n9247 ) ;
assign n9249 =  ( n9242 ) ? ( bv_8_238_n71 ) : ( n9248 ) ;
assign n9250 =  ( n9240 ) ? ( bv_8_246_n39 ) : ( n9249 ) ;
assign n9251 =  ( n9238 ) ? ( bv_8_255_n3 ) : ( n9250 ) ;
assign n9252 =  ( n9236 ) ? ( bv_8_214_n164 ) : ( n9251 ) ;
assign n9253 =  ( n9234 ) ? ( bv_8_222_n134 ) : ( n9252 ) ;
assign n9254 =  ( n9232 ) ? ( bv_8_145_n397 ) : ( n9253 ) ;
assign n9255 =  ( n9230 ) ? ( bv_8_96_n542 ) : ( n9254 ) ;
assign n9256 =  ( n9228 ) ? ( bv_8_2_n751 ) : ( n9255 ) ;
assign n9257 =  ( n9226 ) ? ( bv_8_206_n192 ) : ( n9256 ) ;
assign n9258 =  ( n9224 ) ? ( bv_8_86_n567 ) : ( n9257 ) ;
assign n9259 =  ( n9222 ) ? ( bv_8_231_n99 ) : ( n9258 ) ;
assign n9260 =  ( n9220 ) ? ( bv_8_181_n281 ) : ( n9259 ) ;
assign n9261 =  ( n9218 ) ? ( bv_8_77_n593 ) : ( n9260 ) ;
assign n9262 =  ( n9216 ) ? ( bv_8_236_n79 ) : ( n9261 ) ;
assign n9263 =  ( n9214 ) ? ( bv_8_143_n403 ) : ( n9262 ) ;
assign n9264 =  ( n9212 ) ? ( bv_8_31_n705 ) : ( n9263 ) ;
assign n9265 =  ( n9210 ) ? ( bv_8_137_n421 ) : ( n9264 ) ;
assign n9266 =  ( n9208 ) ? ( bv_8_250_n23 ) : ( n9265 ) ;
assign n9267 =  ( n9206 ) ? ( bv_8_239_n67 ) : ( n9266 ) ;
assign n9268 =  ( n9204 ) ? ( bv_8_178_n292 ) : ( n9267 ) ;
assign n9269 =  ( n9202 ) ? ( bv_8_142_n406 ) : ( n9268 ) ;
assign n9270 =  ( n9200 ) ? ( bv_8_251_n19 ) : ( n9269 ) ;
assign n9271 =  ( n9198 ) ? ( bv_8_65_n623 ) : ( n9270 ) ;
assign n9272 =  ( n9196 ) ? ( bv_8_179_n289 ) : ( n9271 ) ;
assign n9273 =  ( n9194 ) ? ( bv_8_95_n545 ) : ( n9272 ) ;
assign n9274 =  ( n9192 ) ? ( bv_8_69_n612 ) : ( n9273 ) ;
assign n9275 =  ( n9190 ) ? ( bv_8_35_n696 ) : ( n9274 ) ;
assign n9276 =  ( n9188 ) ? ( bv_8_83_n575 ) : ( n9275 ) ;
assign n9277 =  ( n9186 ) ? ( bv_8_228_n111 ) : ( n9276 ) ;
assign n9278 =  ( n9184 ) ? ( bv_8_155_n364 ) : ( n9277 ) ;
assign n9279 =  ( n9182 ) ? ( bv_8_117_n484 ) : ( n9278 ) ;
assign n9280 =  ( n9180 ) ? ( bv_8_225_n123 ) : ( n9279 ) ;
assign n9281 =  ( n9178 ) ? ( bv_8_61_n634 ) : ( n9280 ) ;
assign n9282 =  ( n9176 ) ? ( bv_8_76_n596 ) : ( n9281 ) ;
assign n9283 =  ( n9174 ) ? ( bv_8_108_n510 ) : ( n9282 ) ;
assign n9284 =  ( n9172 ) ? ( bv_8_126_n456 ) : ( n9283 ) ;
assign n9285 =  ( n9170 ) ? ( bv_8_245_n43 ) : ( n9284 ) ;
assign n9286 =  ( n9168 ) ? ( bv_8_131_n440 ) : ( n9285 ) ;
assign n9287 =  ( n9166 ) ? ( bv_8_104_n520 ) : ( n9286 ) ;
assign n9288 =  ( n9164 ) ? ( bv_8_81_n582 ) : ( n9287 ) ;
assign n9289 =  ( n9162 ) ? ( bv_8_209_n182 ) : ( n9288 ) ;
assign n9290 =  ( n9160 ) ? ( bv_8_249_n27 ) : ( n9289 ) ;
assign n9291 =  ( n9158 ) ? ( bv_8_226_n119 ) : ( n9290 ) ;
assign n9292 =  ( n9156 ) ? ( bv_8_171_n314 ) : ( n9291 ) ;
assign n9293 =  ( n9154 ) ? ( bv_8_98_n536 ) : ( n9292 ) ;
assign n9294 =  ( n9152 ) ? ( bv_8_42_n672 ) : ( n9293 ) ;
assign n9295 =  ( n9150 ) ? ( bv_8_8_n669 ) : ( n9294 ) ;
assign n9296 =  ( n9148 ) ? ( bv_8_149_n384 ) : ( n9295 ) ;
assign n9297 =  ( n9146 ) ? ( bv_8_70_n609 ) : ( n9296 ) ;
assign n9298 =  ( n9144 ) ? ( bv_8_157_n359 ) : ( n9297 ) ;
assign n9299 =  ( n9142 ) ? ( bv_8_48_n660 ) : ( n9298 ) ;
assign n9300 =  ( n9140 ) ? ( bv_8_55_n650 ) : ( n9299 ) ;
assign n9301 =  ( n9138 ) ? ( bv_8_10_n655 ) : ( n9300 ) ;
assign n9302 =  ( n9136 ) ? ( bv_8_47_n652 ) : ( n9301 ) ;
assign n9303 =  ( n9134 ) ? ( bv_8_14_n648 ) : ( n9302 ) ;
assign n9304 =  ( n9132 ) ? ( bv_8_36_n645 ) : ( n9303 ) ;
assign n9305 =  ( n9130 ) ? ( bv_8_27_n642 ) : ( n9304 ) ;
assign n9306 =  ( n9128 ) ? ( bv_8_223_n130 ) : ( n9305 ) ;
assign n9307 =  ( n9126 ) ? ( bv_8_205_n196 ) : ( n9306 ) ;
assign n9308 =  ( n9124 ) ? ( bv_8_78_n590 ) : ( n9307 ) ;
assign n9309 =  ( n9122 ) ? ( bv_8_127_n453 ) : ( n9308 ) ;
assign n9310 =  ( n9120 ) ? ( bv_8_234_n87 ) : ( n9309 ) ;
assign n9311 =  ( n9118 ) ? ( bv_8_18_n628 ) : ( n9310 ) ;
assign n9312 =  ( n9116 ) ? ( bv_8_29_n625 ) : ( n9311 ) ;
assign n9313 =  ( n9114 ) ? ( bv_8_88_n562 ) : ( n9312 ) ;
assign n9314 =  ( n9112 ) ? ( bv_8_52_n619 ) : ( n9313 ) ;
assign n9315 =  ( n9110 ) ? ( bv_8_54_n616 ) : ( n9314 ) ;
assign n9316 =  ( n9108 ) ? ( bv_8_220_n142 ) : ( n9315 ) ;
assign n9317 =  ( n9106 ) ? ( bv_8_180_n285 ) : ( n9316 ) ;
assign n9318 =  ( n9104 ) ? ( bv_8_91_n555 ) : ( n9317 ) ;
assign n9319 =  ( n9102 ) ? ( bv_8_164_n335 ) : ( n9318 ) ;
assign n9320 =  ( n9100 ) ? ( bv_8_118_n480 ) : ( n9319 ) ;
assign n9321 =  ( n9098 ) ? ( bv_8_183_n273 ) : ( n9320 ) ;
assign n9322 =  ( n9096 ) ? ( bv_8_125_n459 ) : ( n9321 ) ;
assign n9323 =  ( n9094 ) ? ( bv_8_82_n578 ) : ( n9322 ) ;
assign n9324 =  ( n9092 ) ? ( bv_8_221_n138 ) : ( n9323 ) ;
assign n9325 =  ( n9090 ) ? ( bv_8_94_n548 ) : ( n9324 ) ;
assign n9326 =  ( n9088 ) ? ( bv_8_19_n588 ) : ( n9325 ) ;
assign n9327 =  ( n9086 ) ? ( bv_8_166_n328 ) : ( n9326 ) ;
assign n9328 =  ( n9084 ) ? ( bv_8_185_n266 ) : ( n9327 ) ;
assign n9329 =  ( n9082 ) ? ( bv_8_0_n580 ) : ( n9328 ) ;
assign n9330 =  ( n9080 ) ? ( bv_8_193_n239 ) : ( n9329 ) ;
assign n9331 =  ( n9078 ) ? ( bv_8_64_n573 ) : ( n9330 ) ;
assign n9332 =  ( n9076 ) ? ( bv_8_227_n115 ) : ( n9331 ) ;
assign n9333 =  ( n9074 ) ? ( bv_8_121_n470 ) : ( n9332 ) ;
assign n9334 =  ( n9072 ) ? ( bv_8_182_n277 ) : ( n9333 ) ;
assign n9335 =  ( n9070 ) ? ( bv_8_212_n171 ) : ( n9334 ) ;
assign n9336 =  ( n9068 ) ? ( bv_8_141_n410 ) : ( n9335 ) ;
assign n9337 =  ( n9066 ) ? ( bv_8_103_n523 ) : ( n9336 ) ;
assign n9338 =  ( n9064 ) ? ( bv_8_114_n494 ) : ( n9337 ) ;
assign n9339 =  ( n9062 ) ? ( bv_8_148_n388 ) : ( n9338 ) ;
assign n9340 =  ( n9060 ) ? ( bv_8_152_n374 ) : ( n9339 ) ;
assign n9341 =  ( n9058 ) ? ( bv_8_176_n299 ) : ( n9340 ) ;
assign n9342 =  ( n9056 ) ? ( bv_8_133_n434 ) : ( n9341 ) ;
assign n9343 =  ( n9054 ) ? ( bv_8_187_n260 ) : ( n9342 ) ;
assign n9344 =  ( n9052 ) ? ( bv_8_197_n224 ) : ( n9343 ) ;
assign n9345 =  ( n9050 ) ? ( bv_8_79_n538 ) : ( n9344 ) ;
assign n9346 =  ( n9048 ) ? ( bv_8_237_n75 ) : ( n9345 ) ;
assign n9347 =  ( n9046 ) ? ( bv_8_134_n431 ) : ( n9346 ) ;
assign n9348 =  ( n9044 ) ? ( bv_8_154_n368 ) : ( n9347 ) ;
assign n9349 =  ( n9042 ) ? ( bv_8_102_n527 ) : ( n9348 ) ;
assign n9350 =  ( n9040 ) ? ( bv_8_17_n525 ) : ( n9349 ) ;
assign n9351 =  ( n9038 ) ? ( bv_8_138_n418 ) : ( n9350 ) ;
assign n9352 =  ( n9036 ) ? ( bv_8_233_n91 ) : ( n9351 ) ;
assign n9353 =  ( n9034 ) ? ( bv_8_4_n516 ) : ( n9352 ) ;
assign n9354 =  ( n9032 ) ? ( bv_8_254_n7 ) : ( n9353 ) ;
assign n9355 =  ( n9030 ) ? ( bv_8_160_n350 ) : ( n9354 ) ;
assign n9356 =  ( n9028 ) ? ( bv_8_120_n474 ) : ( n9355 ) ;
assign n9357 =  ( n9026 ) ? ( bv_8_37_n506 ) : ( n9356 ) ;
assign n9358 =  ( n9024 ) ? ( bv_8_75_n503 ) : ( n9357 ) ;
assign n9359 =  ( n9022 ) ? ( bv_8_162_n343 ) : ( n9358 ) ;
assign n9360 =  ( n9020 ) ? ( bv_8_93_n498 ) : ( n9359 ) ;
assign n9361 =  ( n9018 ) ? ( bv_8_128_n450 ) : ( n9360 ) ;
assign n9362 =  ( n9016 ) ? ( bv_8_5_n492 ) : ( n9361 ) ;
assign n9363 =  ( n9014 ) ? ( bv_8_63_n489 ) : ( n9362 ) ;
assign n9364 =  ( n9012 ) ? ( bv_8_33_n486 ) : ( n9363 ) ;
assign n9365 =  ( n9010 ) ? ( bv_8_112_n482 ) : ( n9364 ) ;
assign n9366 =  ( n9008 ) ? ( bv_8_241_n59 ) : ( n9365 ) ;
assign n9367 =  ( n9006 ) ? ( bv_8_99_n476 ) : ( n9366 ) ;
assign n9368 =  ( n9004 ) ? ( bv_8_119_n472 ) : ( n9367 ) ;
assign n9369 =  ( n9002 ) ? ( bv_8_175_n302 ) : ( n9368 ) ;
assign n9370 =  ( n9000 ) ? ( bv_8_66_n466 ) : ( n9369 ) ;
assign n9371 =  ( n8998 ) ? ( bv_8_32_n463 ) : ( n9370 ) ;
assign n9372 =  ( n8996 ) ? ( bv_8_229_n107 ) : ( n9371 ) ;
assign n9373 =  ( n8994 ) ? ( bv_8_253_n11 ) : ( n9372 ) ;
assign n9374 =  ( n8992 ) ? ( bv_8_191_n246 ) : ( n9373 ) ;
assign n9375 =  ( n8990 ) ? ( bv_8_129_n446 ) : ( n9374 ) ;
assign n9376 =  ( n8988 ) ? ( bv_8_24_n448 ) : ( n9375 ) ;
assign n9377 =  ( n8986 ) ? ( bv_8_38_n444 ) : ( n9376 ) ;
assign n9378 =  ( n8984 ) ? ( bv_8_195_n232 ) : ( n9377 ) ;
assign n9379 =  ( n8982 ) ? ( bv_8_190_n250 ) : ( n9378 ) ;
assign n9380 =  ( n8980 ) ? ( bv_8_53_n436 ) : ( n9379 ) ;
assign n9381 =  ( n8978 ) ? ( bv_8_136_n425 ) : ( n9380 ) ;
assign n9382 =  ( n8976 ) ? ( bv_8_46_n429 ) : ( n9381 ) ;
assign n9383 =  ( n8974 ) ? ( bv_8_147_n392 ) : ( n9382 ) ;
assign n9384 =  ( n8972 ) ? ( bv_8_85_n423 ) : ( n9383 ) ;
assign n9385 =  ( n8970 ) ? ( bv_8_252_n15 ) : ( n9384 ) ;
assign n9386 =  ( n8968 ) ? ( bv_8_122_n416 ) : ( n9385 ) ;
assign n9387 =  ( n8966 ) ? ( bv_8_200_n213 ) : ( n9386 ) ;
assign n9388 =  ( n8964 ) ? ( bv_8_186_n263 ) : ( n9387 ) ;
assign n9389 =  ( n8962 ) ? ( bv_8_50_n408 ) : ( n9388 ) ;
assign n9390 =  ( n8960 ) ? ( bv_8_230_n103 ) : ( n9389 ) ;
assign n9391 =  ( n8958 ) ? ( bv_8_192_n242 ) : ( n9390 ) ;
assign n9392 =  ( n8956 ) ? ( bv_8_25_n399 ) : ( n9391 ) ;
assign n9393 =  ( n8954 ) ? ( bv_8_158_n355 ) : ( n9392 ) ;
assign n9394 =  ( n8952 ) ? ( bv_8_163_n339 ) : ( n9393 ) ;
assign n9395 =  ( n8950 ) ? ( bv_8_68_n390 ) : ( n9394 ) ;
assign n9396 =  ( n8948 ) ? ( bv_8_84_n386 ) : ( n9395 ) ;
assign n9397 =  ( n8946 ) ? ( bv_8_59_n382 ) : ( n9396 ) ;
assign n9398 =  ( n8944 ) ? ( bv_8_11_n379 ) : ( n9397 ) ;
assign n9399 =  ( n8942 ) ? ( bv_8_140_n376 ) : ( n9398 ) ;
assign n9400 =  ( n8940 ) ? ( bv_8_199_n216 ) : ( n9399 ) ;
assign n9401 =  ( n8938 ) ? ( bv_8_107_n370 ) : ( n9400 ) ;
assign n9402 =  ( n8936 ) ? ( bv_8_40_n366 ) : ( n9401 ) ;
assign n9403 =  ( n8934 ) ? ( bv_8_167_n325 ) : ( n9402 ) ;
assign n9404 =  ( n8932 ) ? ( bv_8_188_n257 ) : ( n9403 ) ;
assign n9405 =  ( n8930 ) ? ( bv_8_22_n357 ) : ( n9404 ) ;
assign n9406 =  ( n8928 ) ? ( bv_8_173_n307 ) : ( n9405 ) ;
assign n9407 =  ( n8926 ) ? ( bv_8_219_n146 ) : ( n9406 ) ;
assign n9408 =  ( n8924 ) ? ( bv_8_100_n348 ) : ( n9407 ) ;
assign n9409 =  ( n8922 ) ? ( bv_8_116_n345 ) : ( n9408 ) ;
assign n9410 =  ( n8920 ) ? ( bv_8_20_n341 ) : ( n9409 ) ;
assign n9411 =  ( n8918 ) ? ( bv_8_146_n337 ) : ( n9410 ) ;
assign n9412 =  ( n8916 ) ? ( bv_8_12_n333 ) : ( n9411 ) ;
assign n9413 =  ( n8914 ) ? ( bv_8_72_n330 ) : ( n9412 ) ;
assign n9414 =  ( n8912 ) ? ( bv_8_184_n270 ) : ( n9413 ) ;
assign n9415 =  ( n8910 ) ? ( bv_8_159_n323 ) : ( n9414 ) ;
assign n9416 =  ( n8908 ) ? ( bv_8_189_n254 ) : ( n9415 ) ;
assign n9417 =  ( n8906 ) ? ( bv_8_67_n318 ) : ( n9416 ) ;
assign n9418 =  ( n8904 ) ? ( bv_8_196_n228 ) : ( n9417 ) ;
assign n9419 =  ( n8902 ) ? ( bv_8_57_n312 ) : ( n9418 ) ;
assign n9420 =  ( n8900 ) ? ( bv_8_49_n309 ) : ( n9419 ) ;
assign n9421 =  ( n8898 ) ? ( bv_8_211_n175 ) : ( n9420 ) ;
assign n9422 =  ( n8896 ) ? ( bv_8_242_n55 ) : ( n9421 ) ;
assign n9423 =  ( n8894 ) ? ( bv_8_213_n167 ) : ( n9422 ) ;
assign n9424 =  ( n8892 ) ? ( bv_8_139_n297 ) : ( n9423 ) ;
assign n9425 =  ( n8890 ) ? ( bv_8_110_n294 ) : ( n9424 ) ;
assign n9426 =  ( n8888 ) ? ( bv_8_218_n150 ) : ( n9425 ) ;
assign n9427 =  ( n8886 ) ? ( bv_8_1_n287 ) : ( n9426 ) ;
assign n9428 =  ( n8884 ) ? ( bv_8_177_n283 ) : ( n9427 ) ;
assign n9429 =  ( n8882 ) ? ( bv_8_156_n279 ) : ( n9428 ) ;
assign n9430 =  ( n8880 ) ? ( bv_8_73_n275 ) : ( n9429 ) ;
assign n9431 =  ( n8878 ) ? ( bv_8_216_n157 ) : ( n9430 ) ;
assign n9432 =  ( n8876 ) ? ( bv_8_172_n268 ) : ( n9431 ) ;
assign n9433 =  ( n8874 ) ? ( bv_8_243_n51 ) : ( n9432 ) ;
assign n9434 =  ( n8872 ) ? ( bv_8_207_n188 ) : ( n9433 ) ;
assign n9435 =  ( n8870 ) ? ( bv_8_202_n207 ) : ( n9434 ) ;
assign n9436 =  ( n8868 ) ? ( bv_8_244_n47 ) : ( n9435 ) ;
assign n9437 =  ( n8866 ) ? ( bv_8_71_n252 ) : ( n9436 ) ;
assign n9438 =  ( n8864 ) ? ( bv_8_16_n248 ) : ( n9437 ) ;
assign n9439 =  ( n8862 ) ? ( bv_8_111_n244 ) : ( n9438 ) ;
assign n9440 =  ( n8860 ) ? ( bv_8_240_n63 ) : ( n9439 ) ;
assign n9441 =  ( n8858 ) ? ( bv_8_74_n237 ) : ( n9440 ) ;
assign n9442 =  ( n8856 ) ? ( bv_8_92_n234 ) : ( n9441 ) ;
assign n9443 =  ( n8854 ) ? ( bv_8_56_n230 ) : ( n9442 ) ;
assign n9444 =  ( n8852 ) ? ( bv_8_87_n226 ) : ( n9443 ) ;
assign n9445 =  ( n8850 ) ? ( bv_8_115_n222 ) : ( n9444 ) ;
assign n9446 =  ( n8848 ) ? ( bv_8_151_n218 ) : ( n9445 ) ;
assign n9447 =  ( n8846 ) ? ( bv_8_203_n203 ) : ( n9446 ) ;
assign n9448 =  ( n8844 ) ? ( bv_8_161_n211 ) : ( n9447 ) ;
assign n9449 =  ( n8842 ) ? ( bv_8_232_n95 ) : ( n9448 ) ;
assign n9450 =  ( n8840 ) ? ( bv_8_62_n205 ) : ( n9449 ) ;
assign n9451 =  ( n8838 ) ? ( bv_8_150_n201 ) : ( n9450 ) ;
assign n9452 =  ( n8836 ) ? ( bv_8_97_n198 ) : ( n9451 ) ;
assign n9453 =  ( n8834 ) ? ( bv_8_13_n194 ) : ( n9452 ) ;
assign n9454 =  ( n8832 ) ? ( bv_8_15_n190 ) : ( n9453 ) ;
assign n9455 =  ( n8830 ) ? ( bv_8_224_n126 ) : ( n9454 ) ;
assign n9456 =  ( n8828 ) ? ( bv_8_124_n184 ) : ( n9455 ) ;
assign n9457 =  ( n8826 ) ? ( bv_8_113_n180 ) : ( n9456 ) ;
assign n9458 =  ( n8824 ) ? ( bv_8_204_n177 ) : ( n9457 ) ;
assign n9459 =  ( n8822 ) ? ( bv_8_144_n173 ) : ( n9458 ) ;
assign n9460 =  ( n8820 ) ? ( bv_8_6_n169 ) : ( n9459 ) ;
assign n9461 =  ( n8818 ) ? ( bv_8_247_n35 ) : ( n9460 ) ;
assign n9462 =  ( n8816 ) ? ( bv_8_28_n162 ) : ( n9461 ) ;
assign n9463 =  ( n8814 ) ? ( bv_8_194_n159 ) : ( n9462 ) ;
assign n9464 =  ( n8812 ) ? ( bv_8_106_n155 ) : ( n9463 ) ;
assign n9465 =  ( n8810 ) ? ( bv_8_174_n152 ) : ( n9464 ) ;
assign n9466 =  ( n8808 ) ? ( bv_8_105_n148 ) : ( n9465 ) ;
assign n9467 =  ( n8806 ) ? ( bv_8_23_n144 ) : ( n9466 ) ;
assign n9468 =  ( n8804 ) ? ( bv_8_153_n140 ) : ( n9467 ) ;
assign n9469 =  ( n8802 ) ? ( bv_8_58_n136 ) : ( n9468 ) ;
assign n9470 =  ( n8800 ) ? ( bv_8_39_n132 ) : ( n9469 ) ;
assign n9471 =  ( n8798 ) ? ( bv_8_217_n128 ) : ( n9470 ) ;
assign n9472 =  ( n8796 ) ? ( bv_8_235_n83 ) : ( n9471 ) ;
assign n9473 =  ( n8794 ) ? ( bv_8_43_n121 ) : ( n9472 ) ;
assign n9474 =  ( n8792 ) ? ( bv_8_34_n117 ) : ( n9473 ) ;
assign n9475 =  ( n8790 ) ? ( bv_8_210_n113 ) : ( n9474 ) ;
assign n9476 =  ( n8788 ) ? ( bv_8_169_n109 ) : ( n9475 ) ;
assign n9477 =  ( n8786 ) ? ( bv_8_7_n105 ) : ( n9476 ) ;
assign n9478 =  ( n8784 ) ? ( bv_8_51_n101 ) : ( n9477 ) ;
assign n9479 =  ( n8782 ) ? ( bv_8_45_n97 ) : ( n9478 ) ;
assign n9480 =  ( n8780 ) ? ( bv_8_60_n93 ) : ( n9479 ) ;
assign n9481 =  ( n8778 ) ? ( bv_8_21_n89 ) : ( n9480 ) ;
assign n9482 =  ( n8776 ) ? ( bv_8_201_n85 ) : ( n9481 ) ;
assign n9483 =  ( n8774 ) ? ( bv_8_135_n81 ) : ( n9482 ) ;
assign n9484 =  ( n8772 ) ? ( bv_8_170_n77 ) : ( n9483 ) ;
assign n9485 =  ( n8770 ) ? ( bv_8_80_n73 ) : ( n9484 ) ;
assign n9486 =  ( n8768 ) ? ( bv_8_165_n69 ) : ( n9485 ) ;
assign n9487 =  ( n8766 ) ? ( bv_8_3_n65 ) : ( n9486 ) ;
assign n9488 =  ( n8764 ) ? ( bv_8_89_n61 ) : ( n9487 ) ;
assign n9489 =  ( n8762 ) ? ( bv_8_9_n57 ) : ( n9488 ) ;
assign n9490 =  ( n8760 ) ? ( bv_8_26_n53 ) : ( n9489 ) ;
assign n9491 =  ( n8758 ) ? ( bv_8_101_n49 ) : ( n9490 ) ;
assign n9492 =  ( n8756 ) ? ( bv_8_215_n45 ) : ( n9491 ) ;
assign n9493 =  ( n8754 ) ? ( bv_8_132_n41 ) : ( n9492 ) ;
assign n9494 =  ( n8752 ) ? ( bv_8_208_n37 ) : ( n9493 ) ;
assign n9495 =  ( n8750 ) ? ( bv_8_130_n33 ) : ( n9494 ) ;
assign n9496 =  ( n8748 ) ? ( bv_8_41_n29 ) : ( n9495 ) ;
assign n9497 =  ( n8746 ) ? ( bv_8_90_n25 ) : ( n9496 ) ;
assign n9498 =  ( n8744 ) ? ( bv_8_30_n21 ) : ( n9497 ) ;
assign n9499 =  ( n8742 ) ? ( bv_8_123_n17 ) : ( n9498 ) ;
assign n9500 =  ( n8740 ) ? ( bv_8_168_n13 ) : ( n9499 ) ;
assign n9501 =  ( n8738 ) ? ( bv_8_109_n9 ) : ( n9500 ) ;
assign n9502 =  ( n8736 ) ? ( bv_8_44_n5 ) : ( n9501 ) ;
assign n9503 =  ( n8734 ) ^ ( n9502 )  ;
assign n9504 = state_in[15:8] ;
assign n9505 =  ( n9504 ) == ( bv_8_255_n3 )  ;
assign n9506 = state_in[15:8] ;
assign n9507 =  ( n9506 ) == ( bv_8_254_n7 )  ;
assign n9508 = state_in[15:8] ;
assign n9509 =  ( n9508 ) == ( bv_8_253_n11 )  ;
assign n9510 = state_in[15:8] ;
assign n9511 =  ( n9510 ) == ( bv_8_252_n15 )  ;
assign n9512 = state_in[15:8] ;
assign n9513 =  ( n9512 ) == ( bv_8_251_n19 )  ;
assign n9514 = state_in[15:8] ;
assign n9515 =  ( n9514 ) == ( bv_8_250_n23 )  ;
assign n9516 = state_in[15:8] ;
assign n9517 =  ( n9516 ) == ( bv_8_249_n27 )  ;
assign n9518 = state_in[15:8] ;
assign n9519 =  ( n9518 ) == ( bv_8_248_n31 )  ;
assign n9520 = state_in[15:8] ;
assign n9521 =  ( n9520 ) == ( bv_8_247_n35 )  ;
assign n9522 = state_in[15:8] ;
assign n9523 =  ( n9522 ) == ( bv_8_246_n39 )  ;
assign n9524 = state_in[15:8] ;
assign n9525 =  ( n9524 ) == ( bv_8_245_n43 )  ;
assign n9526 = state_in[15:8] ;
assign n9527 =  ( n9526 ) == ( bv_8_244_n47 )  ;
assign n9528 = state_in[15:8] ;
assign n9529 =  ( n9528 ) == ( bv_8_243_n51 )  ;
assign n9530 = state_in[15:8] ;
assign n9531 =  ( n9530 ) == ( bv_8_242_n55 )  ;
assign n9532 = state_in[15:8] ;
assign n9533 =  ( n9532 ) == ( bv_8_241_n59 )  ;
assign n9534 = state_in[15:8] ;
assign n9535 =  ( n9534 ) == ( bv_8_240_n63 )  ;
assign n9536 = state_in[15:8] ;
assign n9537 =  ( n9536 ) == ( bv_8_239_n67 )  ;
assign n9538 = state_in[15:8] ;
assign n9539 =  ( n9538 ) == ( bv_8_238_n71 )  ;
assign n9540 = state_in[15:8] ;
assign n9541 =  ( n9540 ) == ( bv_8_237_n75 )  ;
assign n9542 = state_in[15:8] ;
assign n9543 =  ( n9542 ) == ( bv_8_236_n79 )  ;
assign n9544 = state_in[15:8] ;
assign n9545 =  ( n9544 ) == ( bv_8_235_n83 )  ;
assign n9546 = state_in[15:8] ;
assign n9547 =  ( n9546 ) == ( bv_8_234_n87 )  ;
assign n9548 = state_in[15:8] ;
assign n9549 =  ( n9548 ) == ( bv_8_233_n91 )  ;
assign n9550 = state_in[15:8] ;
assign n9551 =  ( n9550 ) == ( bv_8_232_n95 )  ;
assign n9552 = state_in[15:8] ;
assign n9553 =  ( n9552 ) == ( bv_8_231_n99 )  ;
assign n9554 = state_in[15:8] ;
assign n9555 =  ( n9554 ) == ( bv_8_230_n103 )  ;
assign n9556 = state_in[15:8] ;
assign n9557 =  ( n9556 ) == ( bv_8_229_n107 )  ;
assign n9558 = state_in[15:8] ;
assign n9559 =  ( n9558 ) == ( bv_8_228_n111 )  ;
assign n9560 = state_in[15:8] ;
assign n9561 =  ( n9560 ) == ( bv_8_227_n115 )  ;
assign n9562 = state_in[15:8] ;
assign n9563 =  ( n9562 ) == ( bv_8_226_n119 )  ;
assign n9564 = state_in[15:8] ;
assign n9565 =  ( n9564 ) == ( bv_8_225_n123 )  ;
assign n9566 = state_in[15:8] ;
assign n9567 =  ( n9566 ) == ( bv_8_224_n126 )  ;
assign n9568 = state_in[15:8] ;
assign n9569 =  ( n9568 ) == ( bv_8_223_n130 )  ;
assign n9570 = state_in[15:8] ;
assign n9571 =  ( n9570 ) == ( bv_8_222_n134 )  ;
assign n9572 = state_in[15:8] ;
assign n9573 =  ( n9572 ) == ( bv_8_221_n138 )  ;
assign n9574 = state_in[15:8] ;
assign n9575 =  ( n9574 ) == ( bv_8_220_n142 )  ;
assign n9576 = state_in[15:8] ;
assign n9577 =  ( n9576 ) == ( bv_8_219_n146 )  ;
assign n9578 = state_in[15:8] ;
assign n9579 =  ( n9578 ) == ( bv_8_218_n150 )  ;
assign n9580 = state_in[15:8] ;
assign n9581 =  ( n9580 ) == ( bv_8_217_n128 )  ;
assign n9582 = state_in[15:8] ;
assign n9583 =  ( n9582 ) == ( bv_8_216_n157 )  ;
assign n9584 = state_in[15:8] ;
assign n9585 =  ( n9584 ) == ( bv_8_215_n45 )  ;
assign n9586 = state_in[15:8] ;
assign n9587 =  ( n9586 ) == ( bv_8_214_n164 )  ;
assign n9588 = state_in[15:8] ;
assign n9589 =  ( n9588 ) == ( bv_8_213_n167 )  ;
assign n9590 = state_in[15:8] ;
assign n9591 =  ( n9590 ) == ( bv_8_212_n171 )  ;
assign n9592 = state_in[15:8] ;
assign n9593 =  ( n9592 ) == ( bv_8_211_n175 )  ;
assign n9594 = state_in[15:8] ;
assign n9595 =  ( n9594 ) == ( bv_8_210_n113 )  ;
assign n9596 = state_in[15:8] ;
assign n9597 =  ( n9596 ) == ( bv_8_209_n182 )  ;
assign n9598 = state_in[15:8] ;
assign n9599 =  ( n9598 ) == ( bv_8_208_n37 )  ;
assign n9600 = state_in[15:8] ;
assign n9601 =  ( n9600 ) == ( bv_8_207_n188 )  ;
assign n9602 = state_in[15:8] ;
assign n9603 =  ( n9602 ) == ( bv_8_206_n192 )  ;
assign n9604 = state_in[15:8] ;
assign n9605 =  ( n9604 ) == ( bv_8_205_n196 )  ;
assign n9606 = state_in[15:8] ;
assign n9607 =  ( n9606 ) == ( bv_8_204_n177 )  ;
assign n9608 = state_in[15:8] ;
assign n9609 =  ( n9608 ) == ( bv_8_203_n203 )  ;
assign n9610 = state_in[15:8] ;
assign n9611 =  ( n9610 ) == ( bv_8_202_n207 )  ;
assign n9612 = state_in[15:8] ;
assign n9613 =  ( n9612 ) == ( bv_8_201_n85 )  ;
assign n9614 = state_in[15:8] ;
assign n9615 =  ( n9614 ) == ( bv_8_200_n213 )  ;
assign n9616 = state_in[15:8] ;
assign n9617 =  ( n9616 ) == ( bv_8_199_n216 )  ;
assign n9618 = state_in[15:8] ;
assign n9619 =  ( n9618 ) == ( bv_8_198_n220 )  ;
assign n9620 = state_in[15:8] ;
assign n9621 =  ( n9620 ) == ( bv_8_197_n224 )  ;
assign n9622 = state_in[15:8] ;
assign n9623 =  ( n9622 ) == ( bv_8_196_n228 )  ;
assign n9624 = state_in[15:8] ;
assign n9625 =  ( n9624 ) == ( bv_8_195_n232 )  ;
assign n9626 = state_in[15:8] ;
assign n9627 =  ( n9626 ) == ( bv_8_194_n159 )  ;
assign n9628 = state_in[15:8] ;
assign n9629 =  ( n9628 ) == ( bv_8_193_n239 )  ;
assign n9630 = state_in[15:8] ;
assign n9631 =  ( n9630 ) == ( bv_8_192_n242 )  ;
assign n9632 = state_in[15:8] ;
assign n9633 =  ( n9632 ) == ( bv_8_191_n246 )  ;
assign n9634 = state_in[15:8] ;
assign n9635 =  ( n9634 ) == ( bv_8_190_n250 )  ;
assign n9636 = state_in[15:8] ;
assign n9637 =  ( n9636 ) == ( bv_8_189_n254 )  ;
assign n9638 = state_in[15:8] ;
assign n9639 =  ( n9638 ) == ( bv_8_188_n257 )  ;
assign n9640 = state_in[15:8] ;
assign n9641 =  ( n9640 ) == ( bv_8_187_n260 )  ;
assign n9642 = state_in[15:8] ;
assign n9643 =  ( n9642 ) == ( bv_8_186_n263 )  ;
assign n9644 = state_in[15:8] ;
assign n9645 =  ( n9644 ) == ( bv_8_185_n266 )  ;
assign n9646 = state_in[15:8] ;
assign n9647 =  ( n9646 ) == ( bv_8_184_n270 )  ;
assign n9648 = state_in[15:8] ;
assign n9649 =  ( n9648 ) == ( bv_8_183_n273 )  ;
assign n9650 = state_in[15:8] ;
assign n9651 =  ( n9650 ) == ( bv_8_182_n277 )  ;
assign n9652 = state_in[15:8] ;
assign n9653 =  ( n9652 ) == ( bv_8_181_n281 )  ;
assign n9654 = state_in[15:8] ;
assign n9655 =  ( n9654 ) == ( bv_8_180_n285 )  ;
assign n9656 = state_in[15:8] ;
assign n9657 =  ( n9656 ) == ( bv_8_179_n289 )  ;
assign n9658 = state_in[15:8] ;
assign n9659 =  ( n9658 ) == ( bv_8_178_n292 )  ;
assign n9660 = state_in[15:8] ;
assign n9661 =  ( n9660 ) == ( bv_8_177_n283 )  ;
assign n9662 = state_in[15:8] ;
assign n9663 =  ( n9662 ) == ( bv_8_176_n299 )  ;
assign n9664 = state_in[15:8] ;
assign n9665 =  ( n9664 ) == ( bv_8_175_n302 )  ;
assign n9666 = state_in[15:8] ;
assign n9667 =  ( n9666 ) == ( bv_8_174_n152 )  ;
assign n9668 = state_in[15:8] ;
assign n9669 =  ( n9668 ) == ( bv_8_173_n307 )  ;
assign n9670 = state_in[15:8] ;
assign n9671 =  ( n9670 ) == ( bv_8_172_n268 )  ;
assign n9672 = state_in[15:8] ;
assign n9673 =  ( n9672 ) == ( bv_8_171_n314 )  ;
assign n9674 = state_in[15:8] ;
assign n9675 =  ( n9674 ) == ( bv_8_170_n77 )  ;
assign n9676 = state_in[15:8] ;
assign n9677 =  ( n9676 ) == ( bv_8_169_n109 )  ;
assign n9678 = state_in[15:8] ;
assign n9679 =  ( n9678 ) == ( bv_8_168_n13 )  ;
assign n9680 = state_in[15:8] ;
assign n9681 =  ( n9680 ) == ( bv_8_167_n325 )  ;
assign n9682 = state_in[15:8] ;
assign n9683 =  ( n9682 ) == ( bv_8_166_n328 )  ;
assign n9684 = state_in[15:8] ;
assign n9685 =  ( n9684 ) == ( bv_8_165_n69 )  ;
assign n9686 = state_in[15:8] ;
assign n9687 =  ( n9686 ) == ( bv_8_164_n335 )  ;
assign n9688 = state_in[15:8] ;
assign n9689 =  ( n9688 ) == ( bv_8_163_n339 )  ;
assign n9690 = state_in[15:8] ;
assign n9691 =  ( n9690 ) == ( bv_8_162_n343 )  ;
assign n9692 = state_in[15:8] ;
assign n9693 =  ( n9692 ) == ( bv_8_161_n211 )  ;
assign n9694 = state_in[15:8] ;
assign n9695 =  ( n9694 ) == ( bv_8_160_n350 )  ;
assign n9696 = state_in[15:8] ;
assign n9697 =  ( n9696 ) == ( bv_8_159_n323 )  ;
assign n9698 = state_in[15:8] ;
assign n9699 =  ( n9698 ) == ( bv_8_158_n355 )  ;
assign n9700 = state_in[15:8] ;
assign n9701 =  ( n9700 ) == ( bv_8_157_n359 )  ;
assign n9702 = state_in[15:8] ;
assign n9703 =  ( n9702 ) == ( bv_8_156_n279 )  ;
assign n9704 = state_in[15:8] ;
assign n9705 =  ( n9704 ) == ( bv_8_155_n364 )  ;
assign n9706 = state_in[15:8] ;
assign n9707 =  ( n9706 ) == ( bv_8_154_n368 )  ;
assign n9708 = state_in[15:8] ;
assign n9709 =  ( n9708 ) == ( bv_8_153_n140 )  ;
assign n9710 = state_in[15:8] ;
assign n9711 =  ( n9710 ) == ( bv_8_152_n374 )  ;
assign n9712 = state_in[15:8] ;
assign n9713 =  ( n9712 ) == ( bv_8_151_n218 )  ;
assign n9714 = state_in[15:8] ;
assign n9715 =  ( n9714 ) == ( bv_8_150_n201 )  ;
assign n9716 = state_in[15:8] ;
assign n9717 =  ( n9716 ) == ( bv_8_149_n384 )  ;
assign n9718 = state_in[15:8] ;
assign n9719 =  ( n9718 ) == ( bv_8_148_n388 )  ;
assign n9720 = state_in[15:8] ;
assign n9721 =  ( n9720 ) == ( bv_8_147_n392 )  ;
assign n9722 = state_in[15:8] ;
assign n9723 =  ( n9722 ) == ( bv_8_146_n337 )  ;
assign n9724 = state_in[15:8] ;
assign n9725 =  ( n9724 ) == ( bv_8_145_n397 )  ;
assign n9726 = state_in[15:8] ;
assign n9727 =  ( n9726 ) == ( bv_8_144_n173 )  ;
assign n9728 = state_in[15:8] ;
assign n9729 =  ( n9728 ) == ( bv_8_143_n403 )  ;
assign n9730 = state_in[15:8] ;
assign n9731 =  ( n9730 ) == ( bv_8_142_n406 )  ;
assign n9732 = state_in[15:8] ;
assign n9733 =  ( n9732 ) == ( bv_8_141_n410 )  ;
assign n9734 = state_in[15:8] ;
assign n9735 =  ( n9734 ) == ( bv_8_140_n376 )  ;
assign n9736 = state_in[15:8] ;
assign n9737 =  ( n9736 ) == ( bv_8_139_n297 )  ;
assign n9738 = state_in[15:8] ;
assign n9739 =  ( n9738 ) == ( bv_8_138_n418 )  ;
assign n9740 = state_in[15:8] ;
assign n9741 =  ( n9740 ) == ( bv_8_137_n421 )  ;
assign n9742 = state_in[15:8] ;
assign n9743 =  ( n9742 ) == ( bv_8_136_n425 )  ;
assign n9744 = state_in[15:8] ;
assign n9745 =  ( n9744 ) == ( bv_8_135_n81 )  ;
assign n9746 = state_in[15:8] ;
assign n9747 =  ( n9746 ) == ( bv_8_134_n431 )  ;
assign n9748 = state_in[15:8] ;
assign n9749 =  ( n9748 ) == ( bv_8_133_n434 )  ;
assign n9750 = state_in[15:8] ;
assign n9751 =  ( n9750 ) == ( bv_8_132_n41 )  ;
assign n9752 = state_in[15:8] ;
assign n9753 =  ( n9752 ) == ( bv_8_131_n440 )  ;
assign n9754 = state_in[15:8] ;
assign n9755 =  ( n9754 ) == ( bv_8_130_n33 )  ;
assign n9756 = state_in[15:8] ;
assign n9757 =  ( n9756 ) == ( bv_8_129_n446 )  ;
assign n9758 = state_in[15:8] ;
assign n9759 =  ( n9758 ) == ( bv_8_128_n450 )  ;
assign n9760 = state_in[15:8] ;
assign n9761 =  ( n9760 ) == ( bv_8_127_n453 )  ;
assign n9762 = state_in[15:8] ;
assign n9763 =  ( n9762 ) == ( bv_8_126_n456 )  ;
assign n9764 = state_in[15:8] ;
assign n9765 =  ( n9764 ) == ( bv_8_125_n459 )  ;
assign n9766 = state_in[15:8] ;
assign n9767 =  ( n9766 ) == ( bv_8_124_n184 )  ;
assign n9768 = state_in[15:8] ;
assign n9769 =  ( n9768 ) == ( bv_8_123_n17 )  ;
assign n9770 = state_in[15:8] ;
assign n9771 =  ( n9770 ) == ( bv_8_122_n416 )  ;
assign n9772 = state_in[15:8] ;
assign n9773 =  ( n9772 ) == ( bv_8_121_n470 )  ;
assign n9774 = state_in[15:8] ;
assign n9775 =  ( n9774 ) == ( bv_8_120_n474 )  ;
assign n9776 = state_in[15:8] ;
assign n9777 =  ( n9776 ) == ( bv_8_119_n472 )  ;
assign n9778 = state_in[15:8] ;
assign n9779 =  ( n9778 ) == ( bv_8_118_n480 )  ;
assign n9780 = state_in[15:8] ;
assign n9781 =  ( n9780 ) == ( bv_8_117_n484 )  ;
assign n9782 = state_in[15:8] ;
assign n9783 =  ( n9782 ) == ( bv_8_116_n345 )  ;
assign n9784 = state_in[15:8] ;
assign n9785 =  ( n9784 ) == ( bv_8_115_n222 )  ;
assign n9786 = state_in[15:8] ;
assign n9787 =  ( n9786 ) == ( bv_8_114_n494 )  ;
assign n9788 = state_in[15:8] ;
assign n9789 =  ( n9788 ) == ( bv_8_113_n180 )  ;
assign n9790 = state_in[15:8] ;
assign n9791 =  ( n9790 ) == ( bv_8_112_n482 )  ;
assign n9792 = state_in[15:8] ;
assign n9793 =  ( n9792 ) == ( bv_8_111_n244 )  ;
assign n9794 = state_in[15:8] ;
assign n9795 =  ( n9794 ) == ( bv_8_110_n294 )  ;
assign n9796 = state_in[15:8] ;
assign n9797 =  ( n9796 ) == ( bv_8_109_n9 )  ;
assign n9798 = state_in[15:8] ;
assign n9799 =  ( n9798 ) == ( bv_8_108_n510 )  ;
assign n9800 = state_in[15:8] ;
assign n9801 =  ( n9800 ) == ( bv_8_107_n370 )  ;
assign n9802 = state_in[15:8] ;
assign n9803 =  ( n9802 ) == ( bv_8_106_n155 )  ;
assign n9804 = state_in[15:8] ;
assign n9805 =  ( n9804 ) == ( bv_8_105_n148 )  ;
assign n9806 = state_in[15:8] ;
assign n9807 =  ( n9806 ) == ( bv_8_104_n520 )  ;
assign n9808 = state_in[15:8] ;
assign n9809 =  ( n9808 ) == ( bv_8_103_n523 )  ;
assign n9810 = state_in[15:8] ;
assign n9811 =  ( n9810 ) == ( bv_8_102_n527 )  ;
assign n9812 = state_in[15:8] ;
assign n9813 =  ( n9812 ) == ( bv_8_101_n49 )  ;
assign n9814 = state_in[15:8] ;
assign n9815 =  ( n9814 ) == ( bv_8_100_n348 )  ;
assign n9816 = state_in[15:8] ;
assign n9817 =  ( n9816 ) == ( bv_8_99_n476 )  ;
assign n9818 = state_in[15:8] ;
assign n9819 =  ( n9818 ) == ( bv_8_98_n536 )  ;
assign n9820 = state_in[15:8] ;
assign n9821 =  ( n9820 ) == ( bv_8_97_n198 )  ;
assign n9822 = state_in[15:8] ;
assign n9823 =  ( n9822 ) == ( bv_8_96_n542 )  ;
assign n9824 = state_in[15:8] ;
assign n9825 =  ( n9824 ) == ( bv_8_95_n545 )  ;
assign n9826 = state_in[15:8] ;
assign n9827 =  ( n9826 ) == ( bv_8_94_n548 )  ;
assign n9828 = state_in[15:8] ;
assign n9829 =  ( n9828 ) == ( bv_8_93_n498 )  ;
assign n9830 = state_in[15:8] ;
assign n9831 =  ( n9830 ) == ( bv_8_92_n234 )  ;
assign n9832 = state_in[15:8] ;
assign n9833 =  ( n9832 ) == ( bv_8_91_n555 )  ;
assign n9834 = state_in[15:8] ;
assign n9835 =  ( n9834 ) == ( bv_8_90_n25 )  ;
assign n9836 = state_in[15:8] ;
assign n9837 =  ( n9836 ) == ( bv_8_89_n61 )  ;
assign n9838 = state_in[15:8] ;
assign n9839 =  ( n9838 ) == ( bv_8_88_n562 )  ;
assign n9840 = state_in[15:8] ;
assign n9841 =  ( n9840 ) == ( bv_8_87_n226 )  ;
assign n9842 = state_in[15:8] ;
assign n9843 =  ( n9842 ) == ( bv_8_86_n567 )  ;
assign n9844 = state_in[15:8] ;
assign n9845 =  ( n9844 ) == ( bv_8_85_n423 )  ;
assign n9846 = state_in[15:8] ;
assign n9847 =  ( n9846 ) == ( bv_8_84_n386 )  ;
assign n9848 = state_in[15:8] ;
assign n9849 =  ( n9848 ) == ( bv_8_83_n575 )  ;
assign n9850 = state_in[15:8] ;
assign n9851 =  ( n9850 ) == ( bv_8_82_n578 )  ;
assign n9852 = state_in[15:8] ;
assign n9853 =  ( n9852 ) == ( bv_8_81_n582 )  ;
assign n9854 = state_in[15:8] ;
assign n9855 =  ( n9854 ) == ( bv_8_80_n73 )  ;
assign n9856 = state_in[15:8] ;
assign n9857 =  ( n9856 ) == ( bv_8_79_n538 )  ;
assign n9858 = state_in[15:8] ;
assign n9859 =  ( n9858 ) == ( bv_8_78_n590 )  ;
assign n9860 = state_in[15:8] ;
assign n9861 =  ( n9860 ) == ( bv_8_77_n593 )  ;
assign n9862 = state_in[15:8] ;
assign n9863 =  ( n9862 ) == ( bv_8_76_n596 )  ;
assign n9864 = state_in[15:8] ;
assign n9865 =  ( n9864 ) == ( bv_8_75_n503 )  ;
assign n9866 = state_in[15:8] ;
assign n9867 =  ( n9866 ) == ( bv_8_74_n237 )  ;
assign n9868 = state_in[15:8] ;
assign n9869 =  ( n9868 ) == ( bv_8_73_n275 )  ;
assign n9870 = state_in[15:8] ;
assign n9871 =  ( n9870 ) == ( bv_8_72_n330 )  ;
assign n9872 = state_in[15:8] ;
assign n9873 =  ( n9872 ) == ( bv_8_71_n252 )  ;
assign n9874 = state_in[15:8] ;
assign n9875 =  ( n9874 ) == ( bv_8_70_n609 )  ;
assign n9876 = state_in[15:8] ;
assign n9877 =  ( n9876 ) == ( bv_8_69_n612 )  ;
assign n9878 = state_in[15:8] ;
assign n9879 =  ( n9878 ) == ( bv_8_68_n390 )  ;
assign n9880 = state_in[15:8] ;
assign n9881 =  ( n9880 ) == ( bv_8_67_n318 )  ;
assign n9882 = state_in[15:8] ;
assign n9883 =  ( n9882 ) == ( bv_8_66_n466 )  ;
assign n9884 = state_in[15:8] ;
assign n9885 =  ( n9884 ) == ( bv_8_65_n623 )  ;
assign n9886 = state_in[15:8] ;
assign n9887 =  ( n9886 ) == ( bv_8_64_n573 )  ;
assign n9888 = state_in[15:8] ;
assign n9889 =  ( n9888 ) == ( bv_8_63_n489 )  ;
assign n9890 = state_in[15:8] ;
assign n9891 =  ( n9890 ) == ( bv_8_62_n205 )  ;
assign n9892 = state_in[15:8] ;
assign n9893 =  ( n9892 ) == ( bv_8_61_n634 )  ;
assign n9894 = state_in[15:8] ;
assign n9895 =  ( n9894 ) == ( bv_8_60_n93 )  ;
assign n9896 = state_in[15:8] ;
assign n9897 =  ( n9896 ) == ( bv_8_59_n382 )  ;
assign n9898 = state_in[15:8] ;
assign n9899 =  ( n9898 ) == ( bv_8_58_n136 )  ;
assign n9900 = state_in[15:8] ;
assign n9901 =  ( n9900 ) == ( bv_8_57_n312 )  ;
assign n9902 = state_in[15:8] ;
assign n9903 =  ( n9902 ) == ( bv_8_56_n230 )  ;
assign n9904 = state_in[15:8] ;
assign n9905 =  ( n9904 ) == ( bv_8_55_n650 )  ;
assign n9906 = state_in[15:8] ;
assign n9907 =  ( n9906 ) == ( bv_8_54_n616 )  ;
assign n9908 = state_in[15:8] ;
assign n9909 =  ( n9908 ) == ( bv_8_53_n436 )  ;
assign n9910 = state_in[15:8] ;
assign n9911 =  ( n9910 ) == ( bv_8_52_n619 )  ;
assign n9912 = state_in[15:8] ;
assign n9913 =  ( n9912 ) == ( bv_8_51_n101 )  ;
assign n9914 = state_in[15:8] ;
assign n9915 =  ( n9914 ) == ( bv_8_50_n408 )  ;
assign n9916 = state_in[15:8] ;
assign n9917 =  ( n9916 ) == ( bv_8_49_n309 )  ;
assign n9918 = state_in[15:8] ;
assign n9919 =  ( n9918 ) == ( bv_8_48_n660 )  ;
assign n9920 = state_in[15:8] ;
assign n9921 =  ( n9920 ) == ( bv_8_47_n652 )  ;
assign n9922 = state_in[15:8] ;
assign n9923 =  ( n9922 ) == ( bv_8_46_n429 )  ;
assign n9924 = state_in[15:8] ;
assign n9925 =  ( n9924 ) == ( bv_8_45_n97 )  ;
assign n9926 = state_in[15:8] ;
assign n9927 =  ( n9926 ) == ( bv_8_44_n5 )  ;
assign n9928 = state_in[15:8] ;
assign n9929 =  ( n9928 ) == ( bv_8_43_n121 )  ;
assign n9930 = state_in[15:8] ;
assign n9931 =  ( n9930 ) == ( bv_8_42_n672 )  ;
assign n9932 = state_in[15:8] ;
assign n9933 =  ( n9932 ) == ( bv_8_41_n29 )  ;
assign n9934 = state_in[15:8] ;
assign n9935 =  ( n9934 ) == ( bv_8_40_n366 )  ;
assign n9936 = state_in[15:8] ;
assign n9937 =  ( n9936 ) == ( bv_8_39_n132 )  ;
assign n9938 = state_in[15:8] ;
assign n9939 =  ( n9938 ) == ( bv_8_38_n444 )  ;
assign n9940 = state_in[15:8] ;
assign n9941 =  ( n9940 ) == ( bv_8_37_n506 )  ;
assign n9942 = state_in[15:8] ;
assign n9943 =  ( n9942 ) == ( bv_8_36_n645 )  ;
assign n9944 = state_in[15:8] ;
assign n9945 =  ( n9944 ) == ( bv_8_35_n696 )  ;
assign n9946 = state_in[15:8] ;
assign n9947 =  ( n9946 ) == ( bv_8_34_n117 )  ;
assign n9948 = state_in[15:8] ;
assign n9949 =  ( n9948 ) == ( bv_8_33_n486 )  ;
assign n9950 = state_in[15:8] ;
assign n9951 =  ( n9950 ) == ( bv_8_32_n463 )  ;
assign n9952 = state_in[15:8] ;
assign n9953 =  ( n9952 ) == ( bv_8_31_n705 )  ;
assign n9954 = state_in[15:8] ;
assign n9955 =  ( n9954 ) == ( bv_8_30_n21 )  ;
assign n9956 = state_in[15:8] ;
assign n9957 =  ( n9956 ) == ( bv_8_29_n625 )  ;
assign n9958 = state_in[15:8] ;
assign n9959 =  ( n9958 ) == ( bv_8_28_n162 )  ;
assign n9960 = state_in[15:8] ;
assign n9961 =  ( n9960 ) == ( bv_8_27_n642 )  ;
assign n9962 = state_in[15:8] ;
assign n9963 =  ( n9962 ) == ( bv_8_26_n53 )  ;
assign n9964 = state_in[15:8] ;
assign n9965 =  ( n9964 ) == ( bv_8_25_n399 )  ;
assign n9966 = state_in[15:8] ;
assign n9967 =  ( n9966 ) == ( bv_8_24_n448 )  ;
assign n9968 = state_in[15:8] ;
assign n9969 =  ( n9968 ) == ( bv_8_23_n144 )  ;
assign n9970 = state_in[15:8] ;
assign n9971 =  ( n9970 ) == ( bv_8_22_n357 )  ;
assign n9972 = state_in[15:8] ;
assign n9973 =  ( n9972 ) == ( bv_8_21_n89 )  ;
assign n9974 = state_in[15:8] ;
assign n9975 =  ( n9974 ) == ( bv_8_20_n341 )  ;
assign n9976 = state_in[15:8] ;
assign n9977 =  ( n9976 ) == ( bv_8_19_n588 )  ;
assign n9978 = state_in[15:8] ;
assign n9979 =  ( n9978 ) == ( bv_8_18_n628 )  ;
assign n9980 = state_in[15:8] ;
assign n9981 =  ( n9980 ) == ( bv_8_17_n525 )  ;
assign n9982 = state_in[15:8] ;
assign n9983 =  ( n9982 ) == ( bv_8_16_n248 )  ;
assign n9984 = state_in[15:8] ;
assign n9985 =  ( n9984 ) == ( bv_8_15_n190 )  ;
assign n9986 = state_in[15:8] ;
assign n9987 =  ( n9986 ) == ( bv_8_14_n648 )  ;
assign n9988 = state_in[15:8] ;
assign n9989 =  ( n9988 ) == ( bv_8_13_n194 )  ;
assign n9990 = state_in[15:8] ;
assign n9991 =  ( n9990 ) == ( bv_8_12_n333 )  ;
assign n9992 = state_in[15:8] ;
assign n9993 =  ( n9992 ) == ( bv_8_11_n379 )  ;
assign n9994 = state_in[15:8] ;
assign n9995 =  ( n9994 ) == ( bv_8_10_n655 )  ;
assign n9996 = state_in[15:8] ;
assign n9997 =  ( n9996 ) == ( bv_8_9_n57 )  ;
assign n9998 = state_in[15:8] ;
assign n9999 =  ( n9998 ) == ( bv_8_8_n669 )  ;
assign n10000 = state_in[15:8] ;
assign n10001 =  ( n10000 ) == ( bv_8_7_n105 )  ;
assign n10002 = state_in[15:8] ;
assign n10003 =  ( n10002 ) == ( bv_8_6_n169 )  ;
assign n10004 = state_in[15:8] ;
assign n10005 =  ( n10004 ) == ( bv_8_5_n492 )  ;
assign n10006 = state_in[15:8] ;
assign n10007 =  ( n10006 ) == ( bv_8_4_n516 )  ;
assign n10008 = state_in[15:8] ;
assign n10009 =  ( n10008 ) == ( bv_8_3_n65 )  ;
assign n10010 = state_in[15:8] ;
assign n10011 =  ( n10010 ) == ( bv_8_2_n751 )  ;
assign n10012 = state_in[15:8] ;
assign n10013 =  ( n10012 ) == ( bv_8_1_n287 )  ;
assign n10014 = state_in[15:8] ;
assign n10015 =  ( n10014 ) == ( bv_8_0_n580 )  ;
assign n10016 =  ( n10015 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n10017 =  ( n10013 ) ? ( bv_8_124_n184 ) : ( n10016 ) ;
assign n10018 =  ( n10011 ) ? ( bv_8_119_n472 ) : ( n10017 ) ;
assign n10019 =  ( n10009 ) ? ( bv_8_123_n17 ) : ( n10018 ) ;
assign n10020 =  ( n10007 ) ? ( bv_8_242_n55 ) : ( n10019 ) ;
assign n10021 =  ( n10005 ) ? ( bv_8_107_n370 ) : ( n10020 ) ;
assign n10022 =  ( n10003 ) ? ( bv_8_111_n244 ) : ( n10021 ) ;
assign n10023 =  ( n10001 ) ? ( bv_8_197_n224 ) : ( n10022 ) ;
assign n10024 =  ( n9999 ) ? ( bv_8_48_n660 ) : ( n10023 ) ;
assign n10025 =  ( n9997 ) ? ( bv_8_1_n287 ) : ( n10024 ) ;
assign n10026 =  ( n9995 ) ? ( bv_8_103_n523 ) : ( n10025 ) ;
assign n10027 =  ( n9993 ) ? ( bv_8_43_n121 ) : ( n10026 ) ;
assign n10028 =  ( n9991 ) ? ( bv_8_254_n7 ) : ( n10027 ) ;
assign n10029 =  ( n9989 ) ? ( bv_8_215_n45 ) : ( n10028 ) ;
assign n10030 =  ( n9987 ) ? ( bv_8_171_n314 ) : ( n10029 ) ;
assign n10031 =  ( n9985 ) ? ( bv_8_118_n480 ) : ( n10030 ) ;
assign n10032 =  ( n9983 ) ? ( bv_8_202_n207 ) : ( n10031 ) ;
assign n10033 =  ( n9981 ) ? ( bv_8_130_n33 ) : ( n10032 ) ;
assign n10034 =  ( n9979 ) ? ( bv_8_201_n85 ) : ( n10033 ) ;
assign n10035 =  ( n9977 ) ? ( bv_8_125_n459 ) : ( n10034 ) ;
assign n10036 =  ( n9975 ) ? ( bv_8_250_n23 ) : ( n10035 ) ;
assign n10037 =  ( n9973 ) ? ( bv_8_89_n61 ) : ( n10036 ) ;
assign n10038 =  ( n9971 ) ? ( bv_8_71_n252 ) : ( n10037 ) ;
assign n10039 =  ( n9969 ) ? ( bv_8_240_n63 ) : ( n10038 ) ;
assign n10040 =  ( n9967 ) ? ( bv_8_173_n307 ) : ( n10039 ) ;
assign n10041 =  ( n9965 ) ? ( bv_8_212_n171 ) : ( n10040 ) ;
assign n10042 =  ( n9963 ) ? ( bv_8_162_n343 ) : ( n10041 ) ;
assign n10043 =  ( n9961 ) ? ( bv_8_175_n302 ) : ( n10042 ) ;
assign n10044 =  ( n9959 ) ? ( bv_8_156_n279 ) : ( n10043 ) ;
assign n10045 =  ( n9957 ) ? ( bv_8_164_n335 ) : ( n10044 ) ;
assign n10046 =  ( n9955 ) ? ( bv_8_114_n494 ) : ( n10045 ) ;
assign n10047 =  ( n9953 ) ? ( bv_8_192_n242 ) : ( n10046 ) ;
assign n10048 =  ( n9951 ) ? ( bv_8_183_n273 ) : ( n10047 ) ;
assign n10049 =  ( n9949 ) ? ( bv_8_253_n11 ) : ( n10048 ) ;
assign n10050 =  ( n9947 ) ? ( bv_8_147_n392 ) : ( n10049 ) ;
assign n10051 =  ( n9945 ) ? ( bv_8_38_n444 ) : ( n10050 ) ;
assign n10052 =  ( n9943 ) ? ( bv_8_54_n616 ) : ( n10051 ) ;
assign n10053 =  ( n9941 ) ? ( bv_8_63_n489 ) : ( n10052 ) ;
assign n10054 =  ( n9939 ) ? ( bv_8_247_n35 ) : ( n10053 ) ;
assign n10055 =  ( n9937 ) ? ( bv_8_204_n177 ) : ( n10054 ) ;
assign n10056 =  ( n9935 ) ? ( bv_8_52_n619 ) : ( n10055 ) ;
assign n10057 =  ( n9933 ) ? ( bv_8_165_n69 ) : ( n10056 ) ;
assign n10058 =  ( n9931 ) ? ( bv_8_229_n107 ) : ( n10057 ) ;
assign n10059 =  ( n9929 ) ? ( bv_8_241_n59 ) : ( n10058 ) ;
assign n10060 =  ( n9927 ) ? ( bv_8_113_n180 ) : ( n10059 ) ;
assign n10061 =  ( n9925 ) ? ( bv_8_216_n157 ) : ( n10060 ) ;
assign n10062 =  ( n9923 ) ? ( bv_8_49_n309 ) : ( n10061 ) ;
assign n10063 =  ( n9921 ) ? ( bv_8_21_n89 ) : ( n10062 ) ;
assign n10064 =  ( n9919 ) ? ( bv_8_4_n516 ) : ( n10063 ) ;
assign n10065 =  ( n9917 ) ? ( bv_8_199_n216 ) : ( n10064 ) ;
assign n10066 =  ( n9915 ) ? ( bv_8_35_n696 ) : ( n10065 ) ;
assign n10067 =  ( n9913 ) ? ( bv_8_195_n232 ) : ( n10066 ) ;
assign n10068 =  ( n9911 ) ? ( bv_8_24_n448 ) : ( n10067 ) ;
assign n10069 =  ( n9909 ) ? ( bv_8_150_n201 ) : ( n10068 ) ;
assign n10070 =  ( n9907 ) ? ( bv_8_5_n492 ) : ( n10069 ) ;
assign n10071 =  ( n9905 ) ? ( bv_8_154_n368 ) : ( n10070 ) ;
assign n10072 =  ( n9903 ) ? ( bv_8_7_n105 ) : ( n10071 ) ;
assign n10073 =  ( n9901 ) ? ( bv_8_18_n628 ) : ( n10072 ) ;
assign n10074 =  ( n9899 ) ? ( bv_8_128_n450 ) : ( n10073 ) ;
assign n10075 =  ( n9897 ) ? ( bv_8_226_n119 ) : ( n10074 ) ;
assign n10076 =  ( n9895 ) ? ( bv_8_235_n83 ) : ( n10075 ) ;
assign n10077 =  ( n9893 ) ? ( bv_8_39_n132 ) : ( n10076 ) ;
assign n10078 =  ( n9891 ) ? ( bv_8_178_n292 ) : ( n10077 ) ;
assign n10079 =  ( n9889 ) ? ( bv_8_117_n484 ) : ( n10078 ) ;
assign n10080 =  ( n9887 ) ? ( bv_8_9_n57 ) : ( n10079 ) ;
assign n10081 =  ( n9885 ) ? ( bv_8_131_n440 ) : ( n10080 ) ;
assign n10082 =  ( n9883 ) ? ( bv_8_44_n5 ) : ( n10081 ) ;
assign n10083 =  ( n9881 ) ? ( bv_8_26_n53 ) : ( n10082 ) ;
assign n10084 =  ( n9879 ) ? ( bv_8_27_n642 ) : ( n10083 ) ;
assign n10085 =  ( n9877 ) ? ( bv_8_110_n294 ) : ( n10084 ) ;
assign n10086 =  ( n9875 ) ? ( bv_8_90_n25 ) : ( n10085 ) ;
assign n10087 =  ( n9873 ) ? ( bv_8_160_n350 ) : ( n10086 ) ;
assign n10088 =  ( n9871 ) ? ( bv_8_82_n578 ) : ( n10087 ) ;
assign n10089 =  ( n9869 ) ? ( bv_8_59_n382 ) : ( n10088 ) ;
assign n10090 =  ( n9867 ) ? ( bv_8_214_n164 ) : ( n10089 ) ;
assign n10091 =  ( n9865 ) ? ( bv_8_179_n289 ) : ( n10090 ) ;
assign n10092 =  ( n9863 ) ? ( bv_8_41_n29 ) : ( n10091 ) ;
assign n10093 =  ( n9861 ) ? ( bv_8_227_n115 ) : ( n10092 ) ;
assign n10094 =  ( n9859 ) ? ( bv_8_47_n652 ) : ( n10093 ) ;
assign n10095 =  ( n9857 ) ? ( bv_8_132_n41 ) : ( n10094 ) ;
assign n10096 =  ( n9855 ) ? ( bv_8_83_n575 ) : ( n10095 ) ;
assign n10097 =  ( n9853 ) ? ( bv_8_209_n182 ) : ( n10096 ) ;
assign n10098 =  ( n9851 ) ? ( bv_8_0_n580 ) : ( n10097 ) ;
assign n10099 =  ( n9849 ) ? ( bv_8_237_n75 ) : ( n10098 ) ;
assign n10100 =  ( n9847 ) ? ( bv_8_32_n463 ) : ( n10099 ) ;
assign n10101 =  ( n9845 ) ? ( bv_8_252_n15 ) : ( n10100 ) ;
assign n10102 =  ( n9843 ) ? ( bv_8_177_n283 ) : ( n10101 ) ;
assign n10103 =  ( n9841 ) ? ( bv_8_91_n555 ) : ( n10102 ) ;
assign n10104 =  ( n9839 ) ? ( bv_8_106_n155 ) : ( n10103 ) ;
assign n10105 =  ( n9837 ) ? ( bv_8_203_n203 ) : ( n10104 ) ;
assign n10106 =  ( n9835 ) ? ( bv_8_190_n250 ) : ( n10105 ) ;
assign n10107 =  ( n9833 ) ? ( bv_8_57_n312 ) : ( n10106 ) ;
assign n10108 =  ( n9831 ) ? ( bv_8_74_n237 ) : ( n10107 ) ;
assign n10109 =  ( n9829 ) ? ( bv_8_76_n596 ) : ( n10108 ) ;
assign n10110 =  ( n9827 ) ? ( bv_8_88_n562 ) : ( n10109 ) ;
assign n10111 =  ( n9825 ) ? ( bv_8_207_n188 ) : ( n10110 ) ;
assign n10112 =  ( n9823 ) ? ( bv_8_208_n37 ) : ( n10111 ) ;
assign n10113 =  ( n9821 ) ? ( bv_8_239_n67 ) : ( n10112 ) ;
assign n10114 =  ( n9819 ) ? ( bv_8_170_n77 ) : ( n10113 ) ;
assign n10115 =  ( n9817 ) ? ( bv_8_251_n19 ) : ( n10114 ) ;
assign n10116 =  ( n9815 ) ? ( bv_8_67_n318 ) : ( n10115 ) ;
assign n10117 =  ( n9813 ) ? ( bv_8_77_n593 ) : ( n10116 ) ;
assign n10118 =  ( n9811 ) ? ( bv_8_51_n101 ) : ( n10117 ) ;
assign n10119 =  ( n9809 ) ? ( bv_8_133_n434 ) : ( n10118 ) ;
assign n10120 =  ( n9807 ) ? ( bv_8_69_n612 ) : ( n10119 ) ;
assign n10121 =  ( n9805 ) ? ( bv_8_249_n27 ) : ( n10120 ) ;
assign n10122 =  ( n9803 ) ? ( bv_8_2_n751 ) : ( n10121 ) ;
assign n10123 =  ( n9801 ) ? ( bv_8_127_n453 ) : ( n10122 ) ;
assign n10124 =  ( n9799 ) ? ( bv_8_80_n73 ) : ( n10123 ) ;
assign n10125 =  ( n9797 ) ? ( bv_8_60_n93 ) : ( n10124 ) ;
assign n10126 =  ( n9795 ) ? ( bv_8_159_n323 ) : ( n10125 ) ;
assign n10127 =  ( n9793 ) ? ( bv_8_168_n13 ) : ( n10126 ) ;
assign n10128 =  ( n9791 ) ? ( bv_8_81_n582 ) : ( n10127 ) ;
assign n10129 =  ( n9789 ) ? ( bv_8_163_n339 ) : ( n10128 ) ;
assign n10130 =  ( n9787 ) ? ( bv_8_64_n573 ) : ( n10129 ) ;
assign n10131 =  ( n9785 ) ? ( bv_8_143_n403 ) : ( n10130 ) ;
assign n10132 =  ( n9783 ) ? ( bv_8_146_n337 ) : ( n10131 ) ;
assign n10133 =  ( n9781 ) ? ( bv_8_157_n359 ) : ( n10132 ) ;
assign n10134 =  ( n9779 ) ? ( bv_8_56_n230 ) : ( n10133 ) ;
assign n10135 =  ( n9777 ) ? ( bv_8_245_n43 ) : ( n10134 ) ;
assign n10136 =  ( n9775 ) ? ( bv_8_188_n257 ) : ( n10135 ) ;
assign n10137 =  ( n9773 ) ? ( bv_8_182_n277 ) : ( n10136 ) ;
assign n10138 =  ( n9771 ) ? ( bv_8_218_n150 ) : ( n10137 ) ;
assign n10139 =  ( n9769 ) ? ( bv_8_33_n486 ) : ( n10138 ) ;
assign n10140 =  ( n9767 ) ? ( bv_8_16_n248 ) : ( n10139 ) ;
assign n10141 =  ( n9765 ) ? ( bv_8_255_n3 ) : ( n10140 ) ;
assign n10142 =  ( n9763 ) ? ( bv_8_243_n51 ) : ( n10141 ) ;
assign n10143 =  ( n9761 ) ? ( bv_8_210_n113 ) : ( n10142 ) ;
assign n10144 =  ( n9759 ) ? ( bv_8_205_n196 ) : ( n10143 ) ;
assign n10145 =  ( n9757 ) ? ( bv_8_12_n333 ) : ( n10144 ) ;
assign n10146 =  ( n9755 ) ? ( bv_8_19_n588 ) : ( n10145 ) ;
assign n10147 =  ( n9753 ) ? ( bv_8_236_n79 ) : ( n10146 ) ;
assign n10148 =  ( n9751 ) ? ( bv_8_95_n545 ) : ( n10147 ) ;
assign n10149 =  ( n9749 ) ? ( bv_8_151_n218 ) : ( n10148 ) ;
assign n10150 =  ( n9747 ) ? ( bv_8_68_n390 ) : ( n10149 ) ;
assign n10151 =  ( n9745 ) ? ( bv_8_23_n144 ) : ( n10150 ) ;
assign n10152 =  ( n9743 ) ? ( bv_8_196_n228 ) : ( n10151 ) ;
assign n10153 =  ( n9741 ) ? ( bv_8_167_n325 ) : ( n10152 ) ;
assign n10154 =  ( n9739 ) ? ( bv_8_126_n456 ) : ( n10153 ) ;
assign n10155 =  ( n9737 ) ? ( bv_8_61_n634 ) : ( n10154 ) ;
assign n10156 =  ( n9735 ) ? ( bv_8_100_n348 ) : ( n10155 ) ;
assign n10157 =  ( n9733 ) ? ( bv_8_93_n498 ) : ( n10156 ) ;
assign n10158 =  ( n9731 ) ? ( bv_8_25_n399 ) : ( n10157 ) ;
assign n10159 =  ( n9729 ) ? ( bv_8_115_n222 ) : ( n10158 ) ;
assign n10160 =  ( n9727 ) ? ( bv_8_96_n542 ) : ( n10159 ) ;
assign n10161 =  ( n9725 ) ? ( bv_8_129_n446 ) : ( n10160 ) ;
assign n10162 =  ( n9723 ) ? ( bv_8_79_n538 ) : ( n10161 ) ;
assign n10163 =  ( n9721 ) ? ( bv_8_220_n142 ) : ( n10162 ) ;
assign n10164 =  ( n9719 ) ? ( bv_8_34_n117 ) : ( n10163 ) ;
assign n10165 =  ( n9717 ) ? ( bv_8_42_n672 ) : ( n10164 ) ;
assign n10166 =  ( n9715 ) ? ( bv_8_144_n173 ) : ( n10165 ) ;
assign n10167 =  ( n9713 ) ? ( bv_8_136_n425 ) : ( n10166 ) ;
assign n10168 =  ( n9711 ) ? ( bv_8_70_n609 ) : ( n10167 ) ;
assign n10169 =  ( n9709 ) ? ( bv_8_238_n71 ) : ( n10168 ) ;
assign n10170 =  ( n9707 ) ? ( bv_8_184_n270 ) : ( n10169 ) ;
assign n10171 =  ( n9705 ) ? ( bv_8_20_n341 ) : ( n10170 ) ;
assign n10172 =  ( n9703 ) ? ( bv_8_222_n134 ) : ( n10171 ) ;
assign n10173 =  ( n9701 ) ? ( bv_8_94_n548 ) : ( n10172 ) ;
assign n10174 =  ( n9699 ) ? ( bv_8_11_n379 ) : ( n10173 ) ;
assign n10175 =  ( n9697 ) ? ( bv_8_219_n146 ) : ( n10174 ) ;
assign n10176 =  ( n9695 ) ? ( bv_8_224_n126 ) : ( n10175 ) ;
assign n10177 =  ( n9693 ) ? ( bv_8_50_n408 ) : ( n10176 ) ;
assign n10178 =  ( n9691 ) ? ( bv_8_58_n136 ) : ( n10177 ) ;
assign n10179 =  ( n9689 ) ? ( bv_8_10_n655 ) : ( n10178 ) ;
assign n10180 =  ( n9687 ) ? ( bv_8_73_n275 ) : ( n10179 ) ;
assign n10181 =  ( n9685 ) ? ( bv_8_6_n169 ) : ( n10180 ) ;
assign n10182 =  ( n9683 ) ? ( bv_8_36_n645 ) : ( n10181 ) ;
assign n10183 =  ( n9681 ) ? ( bv_8_92_n234 ) : ( n10182 ) ;
assign n10184 =  ( n9679 ) ? ( bv_8_194_n159 ) : ( n10183 ) ;
assign n10185 =  ( n9677 ) ? ( bv_8_211_n175 ) : ( n10184 ) ;
assign n10186 =  ( n9675 ) ? ( bv_8_172_n268 ) : ( n10185 ) ;
assign n10187 =  ( n9673 ) ? ( bv_8_98_n536 ) : ( n10186 ) ;
assign n10188 =  ( n9671 ) ? ( bv_8_145_n397 ) : ( n10187 ) ;
assign n10189 =  ( n9669 ) ? ( bv_8_149_n384 ) : ( n10188 ) ;
assign n10190 =  ( n9667 ) ? ( bv_8_228_n111 ) : ( n10189 ) ;
assign n10191 =  ( n9665 ) ? ( bv_8_121_n470 ) : ( n10190 ) ;
assign n10192 =  ( n9663 ) ? ( bv_8_231_n99 ) : ( n10191 ) ;
assign n10193 =  ( n9661 ) ? ( bv_8_200_n213 ) : ( n10192 ) ;
assign n10194 =  ( n9659 ) ? ( bv_8_55_n650 ) : ( n10193 ) ;
assign n10195 =  ( n9657 ) ? ( bv_8_109_n9 ) : ( n10194 ) ;
assign n10196 =  ( n9655 ) ? ( bv_8_141_n410 ) : ( n10195 ) ;
assign n10197 =  ( n9653 ) ? ( bv_8_213_n167 ) : ( n10196 ) ;
assign n10198 =  ( n9651 ) ? ( bv_8_78_n590 ) : ( n10197 ) ;
assign n10199 =  ( n9649 ) ? ( bv_8_169_n109 ) : ( n10198 ) ;
assign n10200 =  ( n9647 ) ? ( bv_8_108_n510 ) : ( n10199 ) ;
assign n10201 =  ( n9645 ) ? ( bv_8_86_n567 ) : ( n10200 ) ;
assign n10202 =  ( n9643 ) ? ( bv_8_244_n47 ) : ( n10201 ) ;
assign n10203 =  ( n9641 ) ? ( bv_8_234_n87 ) : ( n10202 ) ;
assign n10204 =  ( n9639 ) ? ( bv_8_101_n49 ) : ( n10203 ) ;
assign n10205 =  ( n9637 ) ? ( bv_8_122_n416 ) : ( n10204 ) ;
assign n10206 =  ( n9635 ) ? ( bv_8_174_n152 ) : ( n10205 ) ;
assign n10207 =  ( n9633 ) ? ( bv_8_8_n669 ) : ( n10206 ) ;
assign n10208 =  ( n9631 ) ? ( bv_8_186_n263 ) : ( n10207 ) ;
assign n10209 =  ( n9629 ) ? ( bv_8_120_n474 ) : ( n10208 ) ;
assign n10210 =  ( n9627 ) ? ( bv_8_37_n506 ) : ( n10209 ) ;
assign n10211 =  ( n9625 ) ? ( bv_8_46_n429 ) : ( n10210 ) ;
assign n10212 =  ( n9623 ) ? ( bv_8_28_n162 ) : ( n10211 ) ;
assign n10213 =  ( n9621 ) ? ( bv_8_166_n328 ) : ( n10212 ) ;
assign n10214 =  ( n9619 ) ? ( bv_8_180_n285 ) : ( n10213 ) ;
assign n10215 =  ( n9617 ) ? ( bv_8_198_n220 ) : ( n10214 ) ;
assign n10216 =  ( n9615 ) ? ( bv_8_232_n95 ) : ( n10215 ) ;
assign n10217 =  ( n9613 ) ? ( bv_8_221_n138 ) : ( n10216 ) ;
assign n10218 =  ( n9611 ) ? ( bv_8_116_n345 ) : ( n10217 ) ;
assign n10219 =  ( n9609 ) ? ( bv_8_31_n705 ) : ( n10218 ) ;
assign n10220 =  ( n9607 ) ? ( bv_8_75_n503 ) : ( n10219 ) ;
assign n10221 =  ( n9605 ) ? ( bv_8_189_n254 ) : ( n10220 ) ;
assign n10222 =  ( n9603 ) ? ( bv_8_139_n297 ) : ( n10221 ) ;
assign n10223 =  ( n9601 ) ? ( bv_8_138_n418 ) : ( n10222 ) ;
assign n10224 =  ( n9599 ) ? ( bv_8_112_n482 ) : ( n10223 ) ;
assign n10225 =  ( n9597 ) ? ( bv_8_62_n205 ) : ( n10224 ) ;
assign n10226 =  ( n9595 ) ? ( bv_8_181_n281 ) : ( n10225 ) ;
assign n10227 =  ( n9593 ) ? ( bv_8_102_n527 ) : ( n10226 ) ;
assign n10228 =  ( n9591 ) ? ( bv_8_72_n330 ) : ( n10227 ) ;
assign n10229 =  ( n9589 ) ? ( bv_8_3_n65 ) : ( n10228 ) ;
assign n10230 =  ( n9587 ) ? ( bv_8_246_n39 ) : ( n10229 ) ;
assign n10231 =  ( n9585 ) ? ( bv_8_14_n648 ) : ( n10230 ) ;
assign n10232 =  ( n9583 ) ? ( bv_8_97_n198 ) : ( n10231 ) ;
assign n10233 =  ( n9581 ) ? ( bv_8_53_n436 ) : ( n10232 ) ;
assign n10234 =  ( n9579 ) ? ( bv_8_87_n226 ) : ( n10233 ) ;
assign n10235 =  ( n9577 ) ? ( bv_8_185_n266 ) : ( n10234 ) ;
assign n10236 =  ( n9575 ) ? ( bv_8_134_n431 ) : ( n10235 ) ;
assign n10237 =  ( n9573 ) ? ( bv_8_193_n239 ) : ( n10236 ) ;
assign n10238 =  ( n9571 ) ? ( bv_8_29_n625 ) : ( n10237 ) ;
assign n10239 =  ( n9569 ) ? ( bv_8_158_n355 ) : ( n10238 ) ;
assign n10240 =  ( n9567 ) ? ( bv_8_225_n123 ) : ( n10239 ) ;
assign n10241 =  ( n9565 ) ? ( bv_8_248_n31 ) : ( n10240 ) ;
assign n10242 =  ( n9563 ) ? ( bv_8_152_n374 ) : ( n10241 ) ;
assign n10243 =  ( n9561 ) ? ( bv_8_17_n525 ) : ( n10242 ) ;
assign n10244 =  ( n9559 ) ? ( bv_8_105_n148 ) : ( n10243 ) ;
assign n10245 =  ( n9557 ) ? ( bv_8_217_n128 ) : ( n10244 ) ;
assign n10246 =  ( n9555 ) ? ( bv_8_142_n406 ) : ( n10245 ) ;
assign n10247 =  ( n9553 ) ? ( bv_8_148_n388 ) : ( n10246 ) ;
assign n10248 =  ( n9551 ) ? ( bv_8_155_n364 ) : ( n10247 ) ;
assign n10249 =  ( n9549 ) ? ( bv_8_30_n21 ) : ( n10248 ) ;
assign n10250 =  ( n9547 ) ? ( bv_8_135_n81 ) : ( n10249 ) ;
assign n10251 =  ( n9545 ) ? ( bv_8_233_n91 ) : ( n10250 ) ;
assign n10252 =  ( n9543 ) ? ( bv_8_206_n192 ) : ( n10251 ) ;
assign n10253 =  ( n9541 ) ? ( bv_8_85_n423 ) : ( n10252 ) ;
assign n10254 =  ( n9539 ) ? ( bv_8_40_n366 ) : ( n10253 ) ;
assign n10255 =  ( n9537 ) ? ( bv_8_223_n130 ) : ( n10254 ) ;
assign n10256 =  ( n9535 ) ? ( bv_8_140_n376 ) : ( n10255 ) ;
assign n10257 =  ( n9533 ) ? ( bv_8_161_n211 ) : ( n10256 ) ;
assign n10258 =  ( n9531 ) ? ( bv_8_137_n421 ) : ( n10257 ) ;
assign n10259 =  ( n9529 ) ? ( bv_8_13_n194 ) : ( n10258 ) ;
assign n10260 =  ( n9527 ) ? ( bv_8_191_n246 ) : ( n10259 ) ;
assign n10261 =  ( n9525 ) ? ( bv_8_230_n103 ) : ( n10260 ) ;
assign n10262 =  ( n9523 ) ? ( bv_8_66_n466 ) : ( n10261 ) ;
assign n10263 =  ( n9521 ) ? ( bv_8_104_n520 ) : ( n10262 ) ;
assign n10264 =  ( n9519 ) ? ( bv_8_65_n623 ) : ( n10263 ) ;
assign n10265 =  ( n9517 ) ? ( bv_8_153_n140 ) : ( n10264 ) ;
assign n10266 =  ( n9515 ) ? ( bv_8_45_n97 ) : ( n10265 ) ;
assign n10267 =  ( n9513 ) ? ( bv_8_15_n190 ) : ( n10266 ) ;
assign n10268 =  ( n9511 ) ? ( bv_8_176_n299 ) : ( n10267 ) ;
assign n10269 =  ( n9509 ) ? ( bv_8_84_n386 ) : ( n10268 ) ;
assign n10270 =  ( n9507 ) ? ( bv_8_187_n260 ) : ( n10269 ) ;
assign n10271 =  ( n9505 ) ? ( bv_8_22_n357 ) : ( n10270 ) ;
assign n10272 =  ( n9503 ) ^ ( n10271 )  ;
assign n10273 = key[95:88] ;
assign n10274 =  ( n10272 ) ^ ( n10273 )  ;
assign n10275 =  { ( n6428 ) , ( n10274 ) }  ;
assign n10276 = state_in[95:88] ;
assign n10277 =  ( n10276 ) == ( bv_8_255_n3 )  ;
assign n10278 = state_in[95:88] ;
assign n10279 =  ( n10278 ) == ( bv_8_254_n7 )  ;
assign n10280 = state_in[95:88] ;
assign n10281 =  ( n10280 ) == ( bv_8_253_n11 )  ;
assign n10282 = state_in[95:88] ;
assign n10283 =  ( n10282 ) == ( bv_8_252_n15 )  ;
assign n10284 = state_in[95:88] ;
assign n10285 =  ( n10284 ) == ( bv_8_251_n19 )  ;
assign n10286 = state_in[95:88] ;
assign n10287 =  ( n10286 ) == ( bv_8_250_n23 )  ;
assign n10288 = state_in[95:88] ;
assign n10289 =  ( n10288 ) == ( bv_8_249_n27 )  ;
assign n10290 = state_in[95:88] ;
assign n10291 =  ( n10290 ) == ( bv_8_248_n31 )  ;
assign n10292 = state_in[95:88] ;
assign n10293 =  ( n10292 ) == ( bv_8_247_n35 )  ;
assign n10294 = state_in[95:88] ;
assign n10295 =  ( n10294 ) == ( bv_8_246_n39 )  ;
assign n10296 = state_in[95:88] ;
assign n10297 =  ( n10296 ) == ( bv_8_245_n43 )  ;
assign n10298 = state_in[95:88] ;
assign n10299 =  ( n10298 ) == ( bv_8_244_n47 )  ;
assign n10300 = state_in[95:88] ;
assign n10301 =  ( n10300 ) == ( bv_8_243_n51 )  ;
assign n10302 = state_in[95:88] ;
assign n10303 =  ( n10302 ) == ( bv_8_242_n55 )  ;
assign n10304 = state_in[95:88] ;
assign n10305 =  ( n10304 ) == ( bv_8_241_n59 )  ;
assign n10306 = state_in[95:88] ;
assign n10307 =  ( n10306 ) == ( bv_8_240_n63 )  ;
assign n10308 = state_in[95:88] ;
assign n10309 =  ( n10308 ) == ( bv_8_239_n67 )  ;
assign n10310 = state_in[95:88] ;
assign n10311 =  ( n10310 ) == ( bv_8_238_n71 )  ;
assign n10312 = state_in[95:88] ;
assign n10313 =  ( n10312 ) == ( bv_8_237_n75 )  ;
assign n10314 = state_in[95:88] ;
assign n10315 =  ( n10314 ) == ( bv_8_236_n79 )  ;
assign n10316 = state_in[95:88] ;
assign n10317 =  ( n10316 ) == ( bv_8_235_n83 )  ;
assign n10318 = state_in[95:88] ;
assign n10319 =  ( n10318 ) == ( bv_8_234_n87 )  ;
assign n10320 = state_in[95:88] ;
assign n10321 =  ( n10320 ) == ( bv_8_233_n91 )  ;
assign n10322 = state_in[95:88] ;
assign n10323 =  ( n10322 ) == ( bv_8_232_n95 )  ;
assign n10324 = state_in[95:88] ;
assign n10325 =  ( n10324 ) == ( bv_8_231_n99 )  ;
assign n10326 = state_in[95:88] ;
assign n10327 =  ( n10326 ) == ( bv_8_230_n103 )  ;
assign n10328 = state_in[95:88] ;
assign n10329 =  ( n10328 ) == ( bv_8_229_n107 )  ;
assign n10330 = state_in[95:88] ;
assign n10331 =  ( n10330 ) == ( bv_8_228_n111 )  ;
assign n10332 = state_in[95:88] ;
assign n10333 =  ( n10332 ) == ( bv_8_227_n115 )  ;
assign n10334 = state_in[95:88] ;
assign n10335 =  ( n10334 ) == ( bv_8_226_n119 )  ;
assign n10336 = state_in[95:88] ;
assign n10337 =  ( n10336 ) == ( bv_8_225_n123 )  ;
assign n10338 = state_in[95:88] ;
assign n10339 =  ( n10338 ) == ( bv_8_224_n126 )  ;
assign n10340 = state_in[95:88] ;
assign n10341 =  ( n10340 ) == ( bv_8_223_n130 )  ;
assign n10342 = state_in[95:88] ;
assign n10343 =  ( n10342 ) == ( bv_8_222_n134 )  ;
assign n10344 = state_in[95:88] ;
assign n10345 =  ( n10344 ) == ( bv_8_221_n138 )  ;
assign n10346 = state_in[95:88] ;
assign n10347 =  ( n10346 ) == ( bv_8_220_n142 )  ;
assign n10348 = state_in[95:88] ;
assign n10349 =  ( n10348 ) == ( bv_8_219_n146 )  ;
assign n10350 = state_in[95:88] ;
assign n10351 =  ( n10350 ) == ( bv_8_218_n150 )  ;
assign n10352 = state_in[95:88] ;
assign n10353 =  ( n10352 ) == ( bv_8_217_n128 )  ;
assign n10354 = state_in[95:88] ;
assign n10355 =  ( n10354 ) == ( bv_8_216_n157 )  ;
assign n10356 = state_in[95:88] ;
assign n10357 =  ( n10356 ) == ( bv_8_215_n45 )  ;
assign n10358 = state_in[95:88] ;
assign n10359 =  ( n10358 ) == ( bv_8_214_n164 )  ;
assign n10360 = state_in[95:88] ;
assign n10361 =  ( n10360 ) == ( bv_8_213_n167 )  ;
assign n10362 = state_in[95:88] ;
assign n10363 =  ( n10362 ) == ( bv_8_212_n171 )  ;
assign n10364 = state_in[95:88] ;
assign n10365 =  ( n10364 ) == ( bv_8_211_n175 )  ;
assign n10366 = state_in[95:88] ;
assign n10367 =  ( n10366 ) == ( bv_8_210_n113 )  ;
assign n10368 = state_in[95:88] ;
assign n10369 =  ( n10368 ) == ( bv_8_209_n182 )  ;
assign n10370 = state_in[95:88] ;
assign n10371 =  ( n10370 ) == ( bv_8_208_n37 )  ;
assign n10372 = state_in[95:88] ;
assign n10373 =  ( n10372 ) == ( bv_8_207_n188 )  ;
assign n10374 = state_in[95:88] ;
assign n10375 =  ( n10374 ) == ( bv_8_206_n192 )  ;
assign n10376 = state_in[95:88] ;
assign n10377 =  ( n10376 ) == ( bv_8_205_n196 )  ;
assign n10378 = state_in[95:88] ;
assign n10379 =  ( n10378 ) == ( bv_8_204_n177 )  ;
assign n10380 = state_in[95:88] ;
assign n10381 =  ( n10380 ) == ( bv_8_203_n203 )  ;
assign n10382 = state_in[95:88] ;
assign n10383 =  ( n10382 ) == ( bv_8_202_n207 )  ;
assign n10384 = state_in[95:88] ;
assign n10385 =  ( n10384 ) == ( bv_8_201_n85 )  ;
assign n10386 = state_in[95:88] ;
assign n10387 =  ( n10386 ) == ( bv_8_200_n213 )  ;
assign n10388 = state_in[95:88] ;
assign n10389 =  ( n10388 ) == ( bv_8_199_n216 )  ;
assign n10390 = state_in[95:88] ;
assign n10391 =  ( n10390 ) == ( bv_8_198_n220 )  ;
assign n10392 = state_in[95:88] ;
assign n10393 =  ( n10392 ) == ( bv_8_197_n224 )  ;
assign n10394 = state_in[95:88] ;
assign n10395 =  ( n10394 ) == ( bv_8_196_n228 )  ;
assign n10396 = state_in[95:88] ;
assign n10397 =  ( n10396 ) == ( bv_8_195_n232 )  ;
assign n10398 = state_in[95:88] ;
assign n10399 =  ( n10398 ) == ( bv_8_194_n159 )  ;
assign n10400 = state_in[95:88] ;
assign n10401 =  ( n10400 ) == ( bv_8_193_n239 )  ;
assign n10402 = state_in[95:88] ;
assign n10403 =  ( n10402 ) == ( bv_8_192_n242 )  ;
assign n10404 = state_in[95:88] ;
assign n10405 =  ( n10404 ) == ( bv_8_191_n246 )  ;
assign n10406 = state_in[95:88] ;
assign n10407 =  ( n10406 ) == ( bv_8_190_n250 )  ;
assign n10408 = state_in[95:88] ;
assign n10409 =  ( n10408 ) == ( bv_8_189_n254 )  ;
assign n10410 = state_in[95:88] ;
assign n10411 =  ( n10410 ) == ( bv_8_188_n257 )  ;
assign n10412 = state_in[95:88] ;
assign n10413 =  ( n10412 ) == ( bv_8_187_n260 )  ;
assign n10414 = state_in[95:88] ;
assign n10415 =  ( n10414 ) == ( bv_8_186_n263 )  ;
assign n10416 = state_in[95:88] ;
assign n10417 =  ( n10416 ) == ( bv_8_185_n266 )  ;
assign n10418 = state_in[95:88] ;
assign n10419 =  ( n10418 ) == ( bv_8_184_n270 )  ;
assign n10420 = state_in[95:88] ;
assign n10421 =  ( n10420 ) == ( bv_8_183_n273 )  ;
assign n10422 = state_in[95:88] ;
assign n10423 =  ( n10422 ) == ( bv_8_182_n277 )  ;
assign n10424 = state_in[95:88] ;
assign n10425 =  ( n10424 ) == ( bv_8_181_n281 )  ;
assign n10426 = state_in[95:88] ;
assign n10427 =  ( n10426 ) == ( bv_8_180_n285 )  ;
assign n10428 = state_in[95:88] ;
assign n10429 =  ( n10428 ) == ( bv_8_179_n289 )  ;
assign n10430 = state_in[95:88] ;
assign n10431 =  ( n10430 ) == ( bv_8_178_n292 )  ;
assign n10432 = state_in[95:88] ;
assign n10433 =  ( n10432 ) == ( bv_8_177_n283 )  ;
assign n10434 = state_in[95:88] ;
assign n10435 =  ( n10434 ) == ( bv_8_176_n299 )  ;
assign n10436 = state_in[95:88] ;
assign n10437 =  ( n10436 ) == ( bv_8_175_n302 )  ;
assign n10438 = state_in[95:88] ;
assign n10439 =  ( n10438 ) == ( bv_8_174_n152 )  ;
assign n10440 = state_in[95:88] ;
assign n10441 =  ( n10440 ) == ( bv_8_173_n307 )  ;
assign n10442 = state_in[95:88] ;
assign n10443 =  ( n10442 ) == ( bv_8_172_n268 )  ;
assign n10444 = state_in[95:88] ;
assign n10445 =  ( n10444 ) == ( bv_8_171_n314 )  ;
assign n10446 = state_in[95:88] ;
assign n10447 =  ( n10446 ) == ( bv_8_170_n77 )  ;
assign n10448 = state_in[95:88] ;
assign n10449 =  ( n10448 ) == ( bv_8_169_n109 )  ;
assign n10450 = state_in[95:88] ;
assign n10451 =  ( n10450 ) == ( bv_8_168_n13 )  ;
assign n10452 = state_in[95:88] ;
assign n10453 =  ( n10452 ) == ( bv_8_167_n325 )  ;
assign n10454 = state_in[95:88] ;
assign n10455 =  ( n10454 ) == ( bv_8_166_n328 )  ;
assign n10456 = state_in[95:88] ;
assign n10457 =  ( n10456 ) == ( bv_8_165_n69 )  ;
assign n10458 = state_in[95:88] ;
assign n10459 =  ( n10458 ) == ( bv_8_164_n335 )  ;
assign n10460 = state_in[95:88] ;
assign n10461 =  ( n10460 ) == ( bv_8_163_n339 )  ;
assign n10462 = state_in[95:88] ;
assign n10463 =  ( n10462 ) == ( bv_8_162_n343 )  ;
assign n10464 = state_in[95:88] ;
assign n10465 =  ( n10464 ) == ( bv_8_161_n211 )  ;
assign n10466 = state_in[95:88] ;
assign n10467 =  ( n10466 ) == ( bv_8_160_n350 )  ;
assign n10468 = state_in[95:88] ;
assign n10469 =  ( n10468 ) == ( bv_8_159_n323 )  ;
assign n10470 = state_in[95:88] ;
assign n10471 =  ( n10470 ) == ( bv_8_158_n355 )  ;
assign n10472 = state_in[95:88] ;
assign n10473 =  ( n10472 ) == ( bv_8_157_n359 )  ;
assign n10474 = state_in[95:88] ;
assign n10475 =  ( n10474 ) == ( bv_8_156_n279 )  ;
assign n10476 = state_in[95:88] ;
assign n10477 =  ( n10476 ) == ( bv_8_155_n364 )  ;
assign n10478 = state_in[95:88] ;
assign n10479 =  ( n10478 ) == ( bv_8_154_n368 )  ;
assign n10480 = state_in[95:88] ;
assign n10481 =  ( n10480 ) == ( bv_8_153_n140 )  ;
assign n10482 = state_in[95:88] ;
assign n10483 =  ( n10482 ) == ( bv_8_152_n374 )  ;
assign n10484 = state_in[95:88] ;
assign n10485 =  ( n10484 ) == ( bv_8_151_n218 )  ;
assign n10486 = state_in[95:88] ;
assign n10487 =  ( n10486 ) == ( bv_8_150_n201 )  ;
assign n10488 = state_in[95:88] ;
assign n10489 =  ( n10488 ) == ( bv_8_149_n384 )  ;
assign n10490 = state_in[95:88] ;
assign n10491 =  ( n10490 ) == ( bv_8_148_n388 )  ;
assign n10492 = state_in[95:88] ;
assign n10493 =  ( n10492 ) == ( bv_8_147_n392 )  ;
assign n10494 = state_in[95:88] ;
assign n10495 =  ( n10494 ) == ( bv_8_146_n337 )  ;
assign n10496 = state_in[95:88] ;
assign n10497 =  ( n10496 ) == ( bv_8_145_n397 )  ;
assign n10498 = state_in[95:88] ;
assign n10499 =  ( n10498 ) == ( bv_8_144_n173 )  ;
assign n10500 = state_in[95:88] ;
assign n10501 =  ( n10500 ) == ( bv_8_143_n403 )  ;
assign n10502 = state_in[95:88] ;
assign n10503 =  ( n10502 ) == ( bv_8_142_n406 )  ;
assign n10504 = state_in[95:88] ;
assign n10505 =  ( n10504 ) == ( bv_8_141_n410 )  ;
assign n10506 = state_in[95:88] ;
assign n10507 =  ( n10506 ) == ( bv_8_140_n376 )  ;
assign n10508 = state_in[95:88] ;
assign n10509 =  ( n10508 ) == ( bv_8_139_n297 )  ;
assign n10510 = state_in[95:88] ;
assign n10511 =  ( n10510 ) == ( bv_8_138_n418 )  ;
assign n10512 = state_in[95:88] ;
assign n10513 =  ( n10512 ) == ( bv_8_137_n421 )  ;
assign n10514 = state_in[95:88] ;
assign n10515 =  ( n10514 ) == ( bv_8_136_n425 )  ;
assign n10516 = state_in[95:88] ;
assign n10517 =  ( n10516 ) == ( bv_8_135_n81 )  ;
assign n10518 = state_in[95:88] ;
assign n10519 =  ( n10518 ) == ( bv_8_134_n431 )  ;
assign n10520 = state_in[95:88] ;
assign n10521 =  ( n10520 ) == ( bv_8_133_n434 )  ;
assign n10522 = state_in[95:88] ;
assign n10523 =  ( n10522 ) == ( bv_8_132_n41 )  ;
assign n10524 = state_in[95:88] ;
assign n10525 =  ( n10524 ) == ( bv_8_131_n440 )  ;
assign n10526 = state_in[95:88] ;
assign n10527 =  ( n10526 ) == ( bv_8_130_n33 )  ;
assign n10528 = state_in[95:88] ;
assign n10529 =  ( n10528 ) == ( bv_8_129_n446 )  ;
assign n10530 = state_in[95:88] ;
assign n10531 =  ( n10530 ) == ( bv_8_128_n450 )  ;
assign n10532 = state_in[95:88] ;
assign n10533 =  ( n10532 ) == ( bv_8_127_n453 )  ;
assign n10534 = state_in[95:88] ;
assign n10535 =  ( n10534 ) == ( bv_8_126_n456 )  ;
assign n10536 = state_in[95:88] ;
assign n10537 =  ( n10536 ) == ( bv_8_125_n459 )  ;
assign n10538 = state_in[95:88] ;
assign n10539 =  ( n10538 ) == ( bv_8_124_n184 )  ;
assign n10540 = state_in[95:88] ;
assign n10541 =  ( n10540 ) == ( bv_8_123_n17 )  ;
assign n10542 = state_in[95:88] ;
assign n10543 =  ( n10542 ) == ( bv_8_122_n416 )  ;
assign n10544 = state_in[95:88] ;
assign n10545 =  ( n10544 ) == ( bv_8_121_n470 )  ;
assign n10546 = state_in[95:88] ;
assign n10547 =  ( n10546 ) == ( bv_8_120_n474 )  ;
assign n10548 = state_in[95:88] ;
assign n10549 =  ( n10548 ) == ( bv_8_119_n472 )  ;
assign n10550 = state_in[95:88] ;
assign n10551 =  ( n10550 ) == ( bv_8_118_n480 )  ;
assign n10552 = state_in[95:88] ;
assign n10553 =  ( n10552 ) == ( bv_8_117_n484 )  ;
assign n10554 = state_in[95:88] ;
assign n10555 =  ( n10554 ) == ( bv_8_116_n345 )  ;
assign n10556 = state_in[95:88] ;
assign n10557 =  ( n10556 ) == ( bv_8_115_n222 )  ;
assign n10558 = state_in[95:88] ;
assign n10559 =  ( n10558 ) == ( bv_8_114_n494 )  ;
assign n10560 = state_in[95:88] ;
assign n10561 =  ( n10560 ) == ( bv_8_113_n180 )  ;
assign n10562 = state_in[95:88] ;
assign n10563 =  ( n10562 ) == ( bv_8_112_n482 )  ;
assign n10564 = state_in[95:88] ;
assign n10565 =  ( n10564 ) == ( bv_8_111_n244 )  ;
assign n10566 = state_in[95:88] ;
assign n10567 =  ( n10566 ) == ( bv_8_110_n294 )  ;
assign n10568 = state_in[95:88] ;
assign n10569 =  ( n10568 ) == ( bv_8_109_n9 )  ;
assign n10570 = state_in[95:88] ;
assign n10571 =  ( n10570 ) == ( bv_8_108_n510 )  ;
assign n10572 = state_in[95:88] ;
assign n10573 =  ( n10572 ) == ( bv_8_107_n370 )  ;
assign n10574 = state_in[95:88] ;
assign n10575 =  ( n10574 ) == ( bv_8_106_n155 )  ;
assign n10576 = state_in[95:88] ;
assign n10577 =  ( n10576 ) == ( bv_8_105_n148 )  ;
assign n10578 = state_in[95:88] ;
assign n10579 =  ( n10578 ) == ( bv_8_104_n520 )  ;
assign n10580 = state_in[95:88] ;
assign n10581 =  ( n10580 ) == ( bv_8_103_n523 )  ;
assign n10582 = state_in[95:88] ;
assign n10583 =  ( n10582 ) == ( bv_8_102_n527 )  ;
assign n10584 = state_in[95:88] ;
assign n10585 =  ( n10584 ) == ( bv_8_101_n49 )  ;
assign n10586 = state_in[95:88] ;
assign n10587 =  ( n10586 ) == ( bv_8_100_n348 )  ;
assign n10588 = state_in[95:88] ;
assign n10589 =  ( n10588 ) == ( bv_8_99_n476 )  ;
assign n10590 = state_in[95:88] ;
assign n10591 =  ( n10590 ) == ( bv_8_98_n536 )  ;
assign n10592 = state_in[95:88] ;
assign n10593 =  ( n10592 ) == ( bv_8_97_n198 )  ;
assign n10594 = state_in[95:88] ;
assign n10595 =  ( n10594 ) == ( bv_8_96_n542 )  ;
assign n10596 = state_in[95:88] ;
assign n10597 =  ( n10596 ) == ( bv_8_95_n545 )  ;
assign n10598 = state_in[95:88] ;
assign n10599 =  ( n10598 ) == ( bv_8_94_n548 )  ;
assign n10600 = state_in[95:88] ;
assign n10601 =  ( n10600 ) == ( bv_8_93_n498 )  ;
assign n10602 = state_in[95:88] ;
assign n10603 =  ( n10602 ) == ( bv_8_92_n234 )  ;
assign n10604 = state_in[95:88] ;
assign n10605 =  ( n10604 ) == ( bv_8_91_n555 )  ;
assign n10606 = state_in[95:88] ;
assign n10607 =  ( n10606 ) == ( bv_8_90_n25 )  ;
assign n10608 = state_in[95:88] ;
assign n10609 =  ( n10608 ) == ( bv_8_89_n61 )  ;
assign n10610 = state_in[95:88] ;
assign n10611 =  ( n10610 ) == ( bv_8_88_n562 )  ;
assign n10612 = state_in[95:88] ;
assign n10613 =  ( n10612 ) == ( bv_8_87_n226 )  ;
assign n10614 = state_in[95:88] ;
assign n10615 =  ( n10614 ) == ( bv_8_86_n567 )  ;
assign n10616 = state_in[95:88] ;
assign n10617 =  ( n10616 ) == ( bv_8_85_n423 )  ;
assign n10618 = state_in[95:88] ;
assign n10619 =  ( n10618 ) == ( bv_8_84_n386 )  ;
assign n10620 = state_in[95:88] ;
assign n10621 =  ( n10620 ) == ( bv_8_83_n575 )  ;
assign n10622 = state_in[95:88] ;
assign n10623 =  ( n10622 ) == ( bv_8_82_n578 )  ;
assign n10624 = state_in[95:88] ;
assign n10625 =  ( n10624 ) == ( bv_8_81_n582 )  ;
assign n10626 = state_in[95:88] ;
assign n10627 =  ( n10626 ) == ( bv_8_80_n73 )  ;
assign n10628 = state_in[95:88] ;
assign n10629 =  ( n10628 ) == ( bv_8_79_n538 )  ;
assign n10630 = state_in[95:88] ;
assign n10631 =  ( n10630 ) == ( bv_8_78_n590 )  ;
assign n10632 = state_in[95:88] ;
assign n10633 =  ( n10632 ) == ( bv_8_77_n593 )  ;
assign n10634 = state_in[95:88] ;
assign n10635 =  ( n10634 ) == ( bv_8_76_n596 )  ;
assign n10636 = state_in[95:88] ;
assign n10637 =  ( n10636 ) == ( bv_8_75_n503 )  ;
assign n10638 = state_in[95:88] ;
assign n10639 =  ( n10638 ) == ( bv_8_74_n237 )  ;
assign n10640 = state_in[95:88] ;
assign n10641 =  ( n10640 ) == ( bv_8_73_n275 )  ;
assign n10642 = state_in[95:88] ;
assign n10643 =  ( n10642 ) == ( bv_8_72_n330 )  ;
assign n10644 = state_in[95:88] ;
assign n10645 =  ( n10644 ) == ( bv_8_71_n252 )  ;
assign n10646 = state_in[95:88] ;
assign n10647 =  ( n10646 ) == ( bv_8_70_n609 )  ;
assign n10648 = state_in[95:88] ;
assign n10649 =  ( n10648 ) == ( bv_8_69_n612 )  ;
assign n10650 = state_in[95:88] ;
assign n10651 =  ( n10650 ) == ( bv_8_68_n390 )  ;
assign n10652 = state_in[95:88] ;
assign n10653 =  ( n10652 ) == ( bv_8_67_n318 )  ;
assign n10654 = state_in[95:88] ;
assign n10655 =  ( n10654 ) == ( bv_8_66_n466 )  ;
assign n10656 = state_in[95:88] ;
assign n10657 =  ( n10656 ) == ( bv_8_65_n623 )  ;
assign n10658 = state_in[95:88] ;
assign n10659 =  ( n10658 ) == ( bv_8_64_n573 )  ;
assign n10660 = state_in[95:88] ;
assign n10661 =  ( n10660 ) == ( bv_8_63_n489 )  ;
assign n10662 = state_in[95:88] ;
assign n10663 =  ( n10662 ) == ( bv_8_62_n205 )  ;
assign n10664 = state_in[95:88] ;
assign n10665 =  ( n10664 ) == ( bv_8_61_n634 )  ;
assign n10666 = state_in[95:88] ;
assign n10667 =  ( n10666 ) == ( bv_8_60_n93 )  ;
assign n10668 = state_in[95:88] ;
assign n10669 =  ( n10668 ) == ( bv_8_59_n382 )  ;
assign n10670 = state_in[95:88] ;
assign n10671 =  ( n10670 ) == ( bv_8_58_n136 )  ;
assign n10672 = state_in[95:88] ;
assign n10673 =  ( n10672 ) == ( bv_8_57_n312 )  ;
assign n10674 = state_in[95:88] ;
assign n10675 =  ( n10674 ) == ( bv_8_56_n230 )  ;
assign n10676 = state_in[95:88] ;
assign n10677 =  ( n10676 ) == ( bv_8_55_n650 )  ;
assign n10678 = state_in[95:88] ;
assign n10679 =  ( n10678 ) == ( bv_8_54_n616 )  ;
assign n10680 = state_in[95:88] ;
assign n10681 =  ( n10680 ) == ( bv_8_53_n436 )  ;
assign n10682 = state_in[95:88] ;
assign n10683 =  ( n10682 ) == ( bv_8_52_n619 )  ;
assign n10684 = state_in[95:88] ;
assign n10685 =  ( n10684 ) == ( bv_8_51_n101 )  ;
assign n10686 = state_in[95:88] ;
assign n10687 =  ( n10686 ) == ( bv_8_50_n408 )  ;
assign n10688 = state_in[95:88] ;
assign n10689 =  ( n10688 ) == ( bv_8_49_n309 )  ;
assign n10690 = state_in[95:88] ;
assign n10691 =  ( n10690 ) == ( bv_8_48_n660 )  ;
assign n10692 = state_in[95:88] ;
assign n10693 =  ( n10692 ) == ( bv_8_47_n652 )  ;
assign n10694 = state_in[95:88] ;
assign n10695 =  ( n10694 ) == ( bv_8_46_n429 )  ;
assign n10696 = state_in[95:88] ;
assign n10697 =  ( n10696 ) == ( bv_8_45_n97 )  ;
assign n10698 = state_in[95:88] ;
assign n10699 =  ( n10698 ) == ( bv_8_44_n5 )  ;
assign n10700 = state_in[95:88] ;
assign n10701 =  ( n10700 ) == ( bv_8_43_n121 )  ;
assign n10702 = state_in[95:88] ;
assign n10703 =  ( n10702 ) == ( bv_8_42_n672 )  ;
assign n10704 = state_in[95:88] ;
assign n10705 =  ( n10704 ) == ( bv_8_41_n29 )  ;
assign n10706 = state_in[95:88] ;
assign n10707 =  ( n10706 ) == ( bv_8_40_n366 )  ;
assign n10708 = state_in[95:88] ;
assign n10709 =  ( n10708 ) == ( bv_8_39_n132 )  ;
assign n10710 = state_in[95:88] ;
assign n10711 =  ( n10710 ) == ( bv_8_38_n444 )  ;
assign n10712 = state_in[95:88] ;
assign n10713 =  ( n10712 ) == ( bv_8_37_n506 )  ;
assign n10714 = state_in[95:88] ;
assign n10715 =  ( n10714 ) == ( bv_8_36_n645 )  ;
assign n10716 = state_in[95:88] ;
assign n10717 =  ( n10716 ) == ( bv_8_35_n696 )  ;
assign n10718 = state_in[95:88] ;
assign n10719 =  ( n10718 ) == ( bv_8_34_n117 )  ;
assign n10720 = state_in[95:88] ;
assign n10721 =  ( n10720 ) == ( bv_8_33_n486 )  ;
assign n10722 = state_in[95:88] ;
assign n10723 =  ( n10722 ) == ( bv_8_32_n463 )  ;
assign n10724 = state_in[95:88] ;
assign n10725 =  ( n10724 ) == ( bv_8_31_n705 )  ;
assign n10726 = state_in[95:88] ;
assign n10727 =  ( n10726 ) == ( bv_8_30_n21 )  ;
assign n10728 = state_in[95:88] ;
assign n10729 =  ( n10728 ) == ( bv_8_29_n625 )  ;
assign n10730 = state_in[95:88] ;
assign n10731 =  ( n10730 ) == ( bv_8_28_n162 )  ;
assign n10732 = state_in[95:88] ;
assign n10733 =  ( n10732 ) == ( bv_8_27_n642 )  ;
assign n10734 = state_in[95:88] ;
assign n10735 =  ( n10734 ) == ( bv_8_26_n53 )  ;
assign n10736 = state_in[95:88] ;
assign n10737 =  ( n10736 ) == ( bv_8_25_n399 )  ;
assign n10738 = state_in[95:88] ;
assign n10739 =  ( n10738 ) == ( bv_8_24_n448 )  ;
assign n10740 = state_in[95:88] ;
assign n10741 =  ( n10740 ) == ( bv_8_23_n144 )  ;
assign n10742 = state_in[95:88] ;
assign n10743 =  ( n10742 ) == ( bv_8_22_n357 )  ;
assign n10744 = state_in[95:88] ;
assign n10745 =  ( n10744 ) == ( bv_8_21_n89 )  ;
assign n10746 = state_in[95:88] ;
assign n10747 =  ( n10746 ) == ( bv_8_20_n341 )  ;
assign n10748 = state_in[95:88] ;
assign n10749 =  ( n10748 ) == ( bv_8_19_n588 )  ;
assign n10750 = state_in[95:88] ;
assign n10751 =  ( n10750 ) == ( bv_8_18_n628 )  ;
assign n10752 = state_in[95:88] ;
assign n10753 =  ( n10752 ) == ( bv_8_17_n525 )  ;
assign n10754 = state_in[95:88] ;
assign n10755 =  ( n10754 ) == ( bv_8_16_n248 )  ;
assign n10756 = state_in[95:88] ;
assign n10757 =  ( n10756 ) == ( bv_8_15_n190 )  ;
assign n10758 = state_in[95:88] ;
assign n10759 =  ( n10758 ) == ( bv_8_14_n648 )  ;
assign n10760 = state_in[95:88] ;
assign n10761 =  ( n10760 ) == ( bv_8_13_n194 )  ;
assign n10762 = state_in[95:88] ;
assign n10763 =  ( n10762 ) == ( bv_8_12_n333 )  ;
assign n10764 = state_in[95:88] ;
assign n10765 =  ( n10764 ) == ( bv_8_11_n379 )  ;
assign n10766 = state_in[95:88] ;
assign n10767 =  ( n10766 ) == ( bv_8_10_n655 )  ;
assign n10768 = state_in[95:88] ;
assign n10769 =  ( n10768 ) == ( bv_8_9_n57 )  ;
assign n10770 = state_in[95:88] ;
assign n10771 =  ( n10770 ) == ( bv_8_8_n669 )  ;
assign n10772 = state_in[95:88] ;
assign n10773 =  ( n10772 ) == ( bv_8_7_n105 )  ;
assign n10774 = state_in[95:88] ;
assign n10775 =  ( n10774 ) == ( bv_8_6_n169 )  ;
assign n10776 = state_in[95:88] ;
assign n10777 =  ( n10776 ) == ( bv_8_5_n492 )  ;
assign n10778 = state_in[95:88] ;
assign n10779 =  ( n10778 ) == ( bv_8_4_n516 )  ;
assign n10780 = state_in[95:88] ;
assign n10781 =  ( n10780 ) == ( bv_8_3_n65 )  ;
assign n10782 = state_in[95:88] ;
assign n10783 =  ( n10782 ) == ( bv_8_2_n751 )  ;
assign n10784 = state_in[95:88] ;
assign n10785 =  ( n10784 ) == ( bv_8_1_n287 )  ;
assign n10786 = state_in[95:88] ;
assign n10787 =  ( n10786 ) == ( bv_8_0_n580 )  ;
assign n10788 =  ( n10787 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n10789 =  ( n10785 ) ? ( bv_8_124_n184 ) : ( n10788 ) ;
assign n10790 =  ( n10783 ) ? ( bv_8_119_n472 ) : ( n10789 ) ;
assign n10791 =  ( n10781 ) ? ( bv_8_123_n17 ) : ( n10790 ) ;
assign n10792 =  ( n10779 ) ? ( bv_8_242_n55 ) : ( n10791 ) ;
assign n10793 =  ( n10777 ) ? ( bv_8_107_n370 ) : ( n10792 ) ;
assign n10794 =  ( n10775 ) ? ( bv_8_111_n244 ) : ( n10793 ) ;
assign n10795 =  ( n10773 ) ? ( bv_8_197_n224 ) : ( n10794 ) ;
assign n10796 =  ( n10771 ) ? ( bv_8_48_n660 ) : ( n10795 ) ;
assign n10797 =  ( n10769 ) ? ( bv_8_1_n287 ) : ( n10796 ) ;
assign n10798 =  ( n10767 ) ? ( bv_8_103_n523 ) : ( n10797 ) ;
assign n10799 =  ( n10765 ) ? ( bv_8_43_n121 ) : ( n10798 ) ;
assign n10800 =  ( n10763 ) ? ( bv_8_254_n7 ) : ( n10799 ) ;
assign n10801 =  ( n10761 ) ? ( bv_8_215_n45 ) : ( n10800 ) ;
assign n10802 =  ( n10759 ) ? ( bv_8_171_n314 ) : ( n10801 ) ;
assign n10803 =  ( n10757 ) ? ( bv_8_118_n480 ) : ( n10802 ) ;
assign n10804 =  ( n10755 ) ? ( bv_8_202_n207 ) : ( n10803 ) ;
assign n10805 =  ( n10753 ) ? ( bv_8_130_n33 ) : ( n10804 ) ;
assign n10806 =  ( n10751 ) ? ( bv_8_201_n85 ) : ( n10805 ) ;
assign n10807 =  ( n10749 ) ? ( bv_8_125_n459 ) : ( n10806 ) ;
assign n10808 =  ( n10747 ) ? ( bv_8_250_n23 ) : ( n10807 ) ;
assign n10809 =  ( n10745 ) ? ( bv_8_89_n61 ) : ( n10808 ) ;
assign n10810 =  ( n10743 ) ? ( bv_8_71_n252 ) : ( n10809 ) ;
assign n10811 =  ( n10741 ) ? ( bv_8_240_n63 ) : ( n10810 ) ;
assign n10812 =  ( n10739 ) ? ( bv_8_173_n307 ) : ( n10811 ) ;
assign n10813 =  ( n10737 ) ? ( bv_8_212_n171 ) : ( n10812 ) ;
assign n10814 =  ( n10735 ) ? ( bv_8_162_n343 ) : ( n10813 ) ;
assign n10815 =  ( n10733 ) ? ( bv_8_175_n302 ) : ( n10814 ) ;
assign n10816 =  ( n10731 ) ? ( bv_8_156_n279 ) : ( n10815 ) ;
assign n10817 =  ( n10729 ) ? ( bv_8_164_n335 ) : ( n10816 ) ;
assign n10818 =  ( n10727 ) ? ( bv_8_114_n494 ) : ( n10817 ) ;
assign n10819 =  ( n10725 ) ? ( bv_8_192_n242 ) : ( n10818 ) ;
assign n10820 =  ( n10723 ) ? ( bv_8_183_n273 ) : ( n10819 ) ;
assign n10821 =  ( n10721 ) ? ( bv_8_253_n11 ) : ( n10820 ) ;
assign n10822 =  ( n10719 ) ? ( bv_8_147_n392 ) : ( n10821 ) ;
assign n10823 =  ( n10717 ) ? ( bv_8_38_n444 ) : ( n10822 ) ;
assign n10824 =  ( n10715 ) ? ( bv_8_54_n616 ) : ( n10823 ) ;
assign n10825 =  ( n10713 ) ? ( bv_8_63_n489 ) : ( n10824 ) ;
assign n10826 =  ( n10711 ) ? ( bv_8_247_n35 ) : ( n10825 ) ;
assign n10827 =  ( n10709 ) ? ( bv_8_204_n177 ) : ( n10826 ) ;
assign n10828 =  ( n10707 ) ? ( bv_8_52_n619 ) : ( n10827 ) ;
assign n10829 =  ( n10705 ) ? ( bv_8_165_n69 ) : ( n10828 ) ;
assign n10830 =  ( n10703 ) ? ( bv_8_229_n107 ) : ( n10829 ) ;
assign n10831 =  ( n10701 ) ? ( bv_8_241_n59 ) : ( n10830 ) ;
assign n10832 =  ( n10699 ) ? ( bv_8_113_n180 ) : ( n10831 ) ;
assign n10833 =  ( n10697 ) ? ( bv_8_216_n157 ) : ( n10832 ) ;
assign n10834 =  ( n10695 ) ? ( bv_8_49_n309 ) : ( n10833 ) ;
assign n10835 =  ( n10693 ) ? ( bv_8_21_n89 ) : ( n10834 ) ;
assign n10836 =  ( n10691 ) ? ( bv_8_4_n516 ) : ( n10835 ) ;
assign n10837 =  ( n10689 ) ? ( bv_8_199_n216 ) : ( n10836 ) ;
assign n10838 =  ( n10687 ) ? ( bv_8_35_n696 ) : ( n10837 ) ;
assign n10839 =  ( n10685 ) ? ( bv_8_195_n232 ) : ( n10838 ) ;
assign n10840 =  ( n10683 ) ? ( bv_8_24_n448 ) : ( n10839 ) ;
assign n10841 =  ( n10681 ) ? ( bv_8_150_n201 ) : ( n10840 ) ;
assign n10842 =  ( n10679 ) ? ( bv_8_5_n492 ) : ( n10841 ) ;
assign n10843 =  ( n10677 ) ? ( bv_8_154_n368 ) : ( n10842 ) ;
assign n10844 =  ( n10675 ) ? ( bv_8_7_n105 ) : ( n10843 ) ;
assign n10845 =  ( n10673 ) ? ( bv_8_18_n628 ) : ( n10844 ) ;
assign n10846 =  ( n10671 ) ? ( bv_8_128_n450 ) : ( n10845 ) ;
assign n10847 =  ( n10669 ) ? ( bv_8_226_n119 ) : ( n10846 ) ;
assign n10848 =  ( n10667 ) ? ( bv_8_235_n83 ) : ( n10847 ) ;
assign n10849 =  ( n10665 ) ? ( bv_8_39_n132 ) : ( n10848 ) ;
assign n10850 =  ( n10663 ) ? ( bv_8_178_n292 ) : ( n10849 ) ;
assign n10851 =  ( n10661 ) ? ( bv_8_117_n484 ) : ( n10850 ) ;
assign n10852 =  ( n10659 ) ? ( bv_8_9_n57 ) : ( n10851 ) ;
assign n10853 =  ( n10657 ) ? ( bv_8_131_n440 ) : ( n10852 ) ;
assign n10854 =  ( n10655 ) ? ( bv_8_44_n5 ) : ( n10853 ) ;
assign n10855 =  ( n10653 ) ? ( bv_8_26_n53 ) : ( n10854 ) ;
assign n10856 =  ( n10651 ) ? ( bv_8_27_n642 ) : ( n10855 ) ;
assign n10857 =  ( n10649 ) ? ( bv_8_110_n294 ) : ( n10856 ) ;
assign n10858 =  ( n10647 ) ? ( bv_8_90_n25 ) : ( n10857 ) ;
assign n10859 =  ( n10645 ) ? ( bv_8_160_n350 ) : ( n10858 ) ;
assign n10860 =  ( n10643 ) ? ( bv_8_82_n578 ) : ( n10859 ) ;
assign n10861 =  ( n10641 ) ? ( bv_8_59_n382 ) : ( n10860 ) ;
assign n10862 =  ( n10639 ) ? ( bv_8_214_n164 ) : ( n10861 ) ;
assign n10863 =  ( n10637 ) ? ( bv_8_179_n289 ) : ( n10862 ) ;
assign n10864 =  ( n10635 ) ? ( bv_8_41_n29 ) : ( n10863 ) ;
assign n10865 =  ( n10633 ) ? ( bv_8_227_n115 ) : ( n10864 ) ;
assign n10866 =  ( n10631 ) ? ( bv_8_47_n652 ) : ( n10865 ) ;
assign n10867 =  ( n10629 ) ? ( bv_8_132_n41 ) : ( n10866 ) ;
assign n10868 =  ( n10627 ) ? ( bv_8_83_n575 ) : ( n10867 ) ;
assign n10869 =  ( n10625 ) ? ( bv_8_209_n182 ) : ( n10868 ) ;
assign n10870 =  ( n10623 ) ? ( bv_8_0_n580 ) : ( n10869 ) ;
assign n10871 =  ( n10621 ) ? ( bv_8_237_n75 ) : ( n10870 ) ;
assign n10872 =  ( n10619 ) ? ( bv_8_32_n463 ) : ( n10871 ) ;
assign n10873 =  ( n10617 ) ? ( bv_8_252_n15 ) : ( n10872 ) ;
assign n10874 =  ( n10615 ) ? ( bv_8_177_n283 ) : ( n10873 ) ;
assign n10875 =  ( n10613 ) ? ( bv_8_91_n555 ) : ( n10874 ) ;
assign n10876 =  ( n10611 ) ? ( bv_8_106_n155 ) : ( n10875 ) ;
assign n10877 =  ( n10609 ) ? ( bv_8_203_n203 ) : ( n10876 ) ;
assign n10878 =  ( n10607 ) ? ( bv_8_190_n250 ) : ( n10877 ) ;
assign n10879 =  ( n10605 ) ? ( bv_8_57_n312 ) : ( n10878 ) ;
assign n10880 =  ( n10603 ) ? ( bv_8_74_n237 ) : ( n10879 ) ;
assign n10881 =  ( n10601 ) ? ( bv_8_76_n596 ) : ( n10880 ) ;
assign n10882 =  ( n10599 ) ? ( bv_8_88_n562 ) : ( n10881 ) ;
assign n10883 =  ( n10597 ) ? ( bv_8_207_n188 ) : ( n10882 ) ;
assign n10884 =  ( n10595 ) ? ( bv_8_208_n37 ) : ( n10883 ) ;
assign n10885 =  ( n10593 ) ? ( bv_8_239_n67 ) : ( n10884 ) ;
assign n10886 =  ( n10591 ) ? ( bv_8_170_n77 ) : ( n10885 ) ;
assign n10887 =  ( n10589 ) ? ( bv_8_251_n19 ) : ( n10886 ) ;
assign n10888 =  ( n10587 ) ? ( bv_8_67_n318 ) : ( n10887 ) ;
assign n10889 =  ( n10585 ) ? ( bv_8_77_n593 ) : ( n10888 ) ;
assign n10890 =  ( n10583 ) ? ( bv_8_51_n101 ) : ( n10889 ) ;
assign n10891 =  ( n10581 ) ? ( bv_8_133_n434 ) : ( n10890 ) ;
assign n10892 =  ( n10579 ) ? ( bv_8_69_n612 ) : ( n10891 ) ;
assign n10893 =  ( n10577 ) ? ( bv_8_249_n27 ) : ( n10892 ) ;
assign n10894 =  ( n10575 ) ? ( bv_8_2_n751 ) : ( n10893 ) ;
assign n10895 =  ( n10573 ) ? ( bv_8_127_n453 ) : ( n10894 ) ;
assign n10896 =  ( n10571 ) ? ( bv_8_80_n73 ) : ( n10895 ) ;
assign n10897 =  ( n10569 ) ? ( bv_8_60_n93 ) : ( n10896 ) ;
assign n10898 =  ( n10567 ) ? ( bv_8_159_n323 ) : ( n10897 ) ;
assign n10899 =  ( n10565 ) ? ( bv_8_168_n13 ) : ( n10898 ) ;
assign n10900 =  ( n10563 ) ? ( bv_8_81_n582 ) : ( n10899 ) ;
assign n10901 =  ( n10561 ) ? ( bv_8_163_n339 ) : ( n10900 ) ;
assign n10902 =  ( n10559 ) ? ( bv_8_64_n573 ) : ( n10901 ) ;
assign n10903 =  ( n10557 ) ? ( bv_8_143_n403 ) : ( n10902 ) ;
assign n10904 =  ( n10555 ) ? ( bv_8_146_n337 ) : ( n10903 ) ;
assign n10905 =  ( n10553 ) ? ( bv_8_157_n359 ) : ( n10904 ) ;
assign n10906 =  ( n10551 ) ? ( bv_8_56_n230 ) : ( n10905 ) ;
assign n10907 =  ( n10549 ) ? ( bv_8_245_n43 ) : ( n10906 ) ;
assign n10908 =  ( n10547 ) ? ( bv_8_188_n257 ) : ( n10907 ) ;
assign n10909 =  ( n10545 ) ? ( bv_8_182_n277 ) : ( n10908 ) ;
assign n10910 =  ( n10543 ) ? ( bv_8_218_n150 ) : ( n10909 ) ;
assign n10911 =  ( n10541 ) ? ( bv_8_33_n486 ) : ( n10910 ) ;
assign n10912 =  ( n10539 ) ? ( bv_8_16_n248 ) : ( n10911 ) ;
assign n10913 =  ( n10537 ) ? ( bv_8_255_n3 ) : ( n10912 ) ;
assign n10914 =  ( n10535 ) ? ( bv_8_243_n51 ) : ( n10913 ) ;
assign n10915 =  ( n10533 ) ? ( bv_8_210_n113 ) : ( n10914 ) ;
assign n10916 =  ( n10531 ) ? ( bv_8_205_n196 ) : ( n10915 ) ;
assign n10917 =  ( n10529 ) ? ( bv_8_12_n333 ) : ( n10916 ) ;
assign n10918 =  ( n10527 ) ? ( bv_8_19_n588 ) : ( n10917 ) ;
assign n10919 =  ( n10525 ) ? ( bv_8_236_n79 ) : ( n10918 ) ;
assign n10920 =  ( n10523 ) ? ( bv_8_95_n545 ) : ( n10919 ) ;
assign n10921 =  ( n10521 ) ? ( bv_8_151_n218 ) : ( n10920 ) ;
assign n10922 =  ( n10519 ) ? ( bv_8_68_n390 ) : ( n10921 ) ;
assign n10923 =  ( n10517 ) ? ( bv_8_23_n144 ) : ( n10922 ) ;
assign n10924 =  ( n10515 ) ? ( bv_8_196_n228 ) : ( n10923 ) ;
assign n10925 =  ( n10513 ) ? ( bv_8_167_n325 ) : ( n10924 ) ;
assign n10926 =  ( n10511 ) ? ( bv_8_126_n456 ) : ( n10925 ) ;
assign n10927 =  ( n10509 ) ? ( bv_8_61_n634 ) : ( n10926 ) ;
assign n10928 =  ( n10507 ) ? ( bv_8_100_n348 ) : ( n10927 ) ;
assign n10929 =  ( n10505 ) ? ( bv_8_93_n498 ) : ( n10928 ) ;
assign n10930 =  ( n10503 ) ? ( bv_8_25_n399 ) : ( n10929 ) ;
assign n10931 =  ( n10501 ) ? ( bv_8_115_n222 ) : ( n10930 ) ;
assign n10932 =  ( n10499 ) ? ( bv_8_96_n542 ) : ( n10931 ) ;
assign n10933 =  ( n10497 ) ? ( bv_8_129_n446 ) : ( n10932 ) ;
assign n10934 =  ( n10495 ) ? ( bv_8_79_n538 ) : ( n10933 ) ;
assign n10935 =  ( n10493 ) ? ( bv_8_220_n142 ) : ( n10934 ) ;
assign n10936 =  ( n10491 ) ? ( bv_8_34_n117 ) : ( n10935 ) ;
assign n10937 =  ( n10489 ) ? ( bv_8_42_n672 ) : ( n10936 ) ;
assign n10938 =  ( n10487 ) ? ( bv_8_144_n173 ) : ( n10937 ) ;
assign n10939 =  ( n10485 ) ? ( bv_8_136_n425 ) : ( n10938 ) ;
assign n10940 =  ( n10483 ) ? ( bv_8_70_n609 ) : ( n10939 ) ;
assign n10941 =  ( n10481 ) ? ( bv_8_238_n71 ) : ( n10940 ) ;
assign n10942 =  ( n10479 ) ? ( bv_8_184_n270 ) : ( n10941 ) ;
assign n10943 =  ( n10477 ) ? ( bv_8_20_n341 ) : ( n10942 ) ;
assign n10944 =  ( n10475 ) ? ( bv_8_222_n134 ) : ( n10943 ) ;
assign n10945 =  ( n10473 ) ? ( bv_8_94_n548 ) : ( n10944 ) ;
assign n10946 =  ( n10471 ) ? ( bv_8_11_n379 ) : ( n10945 ) ;
assign n10947 =  ( n10469 ) ? ( bv_8_219_n146 ) : ( n10946 ) ;
assign n10948 =  ( n10467 ) ? ( bv_8_224_n126 ) : ( n10947 ) ;
assign n10949 =  ( n10465 ) ? ( bv_8_50_n408 ) : ( n10948 ) ;
assign n10950 =  ( n10463 ) ? ( bv_8_58_n136 ) : ( n10949 ) ;
assign n10951 =  ( n10461 ) ? ( bv_8_10_n655 ) : ( n10950 ) ;
assign n10952 =  ( n10459 ) ? ( bv_8_73_n275 ) : ( n10951 ) ;
assign n10953 =  ( n10457 ) ? ( bv_8_6_n169 ) : ( n10952 ) ;
assign n10954 =  ( n10455 ) ? ( bv_8_36_n645 ) : ( n10953 ) ;
assign n10955 =  ( n10453 ) ? ( bv_8_92_n234 ) : ( n10954 ) ;
assign n10956 =  ( n10451 ) ? ( bv_8_194_n159 ) : ( n10955 ) ;
assign n10957 =  ( n10449 ) ? ( bv_8_211_n175 ) : ( n10956 ) ;
assign n10958 =  ( n10447 ) ? ( bv_8_172_n268 ) : ( n10957 ) ;
assign n10959 =  ( n10445 ) ? ( bv_8_98_n536 ) : ( n10958 ) ;
assign n10960 =  ( n10443 ) ? ( bv_8_145_n397 ) : ( n10959 ) ;
assign n10961 =  ( n10441 ) ? ( bv_8_149_n384 ) : ( n10960 ) ;
assign n10962 =  ( n10439 ) ? ( bv_8_228_n111 ) : ( n10961 ) ;
assign n10963 =  ( n10437 ) ? ( bv_8_121_n470 ) : ( n10962 ) ;
assign n10964 =  ( n10435 ) ? ( bv_8_231_n99 ) : ( n10963 ) ;
assign n10965 =  ( n10433 ) ? ( bv_8_200_n213 ) : ( n10964 ) ;
assign n10966 =  ( n10431 ) ? ( bv_8_55_n650 ) : ( n10965 ) ;
assign n10967 =  ( n10429 ) ? ( bv_8_109_n9 ) : ( n10966 ) ;
assign n10968 =  ( n10427 ) ? ( bv_8_141_n410 ) : ( n10967 ) ;
assign n10969 =  ( n10425 ) ? ( bv_8_213_n167 ) : ( n10968 ) ;
assign n10970 =  ( n10423 ) ? ( bv_8_78_n590 ) : ( n10969 ) ;
assign n10971 =  ( n10421 ) ? ( bv_8_169_n109 ) : ( n10970 ) ;
assign n10972 =  ( n10419 ) ? ( bv_8_108_n510 ) : ( n10971 ) ;
assign n10973 =  ( n10417 ) ? ( bv_8_86_n567 ) : ( n10972 ) ;
assign n10974 =  ( n10415 ) ? ( bv_8_244_n47 ) : ( n10973 ) ;
assign n10975 =  ( n10413 ) ? ( bv_8_234_n87 ) : ( n10974 ) ;
assign n10976 =  ( n10411 ) ? ( bv_8_101_n49 ) : ( n10975 ) ;
assign n10977 =  ( n10409 ) ? ( bv_8_122_n416 ) : ( n10976 ) ;
assign n10978 =  ( n10407 ) ? ( bv_8_174_n152 ) : ( n10977 ) ;
assign n10979 =  ( n10405 ) ? ( bv_8_8_n669 ) : ( n10978 ) ;
assign n10980 =  ( n10403 ) ? ( bv_8_186_n263 ) : ( n10979 ) ;
assign n10981 =  ( n10401 ) ? ( bv_8_120_n474 ) : ( n10980 ) ;
assign n10982 =  ( n10399 ) ? ( bv_8_37_n506 ) : ( n10981 ) ;
assign n10983 =  ( n10397 ) ? ( bv_8_46_n429 ) : ( n10982 ) ;
assign n10984 =  ( n10395 ) ? ( bv_8_28_n162 ) : ( n10983 ) ;
assign n10985 =  ( n10393 ) ? ( bv_8_166_n328 ) : ( n10984 ) ;
assign n10986 =  ( n10391 ) ? ( bv_8_180_n285 ) : ( n10985 ) ;
assign n10987 =  ( n10389 ) ? ( bv_8_198_n220 ) : ( n10986 ) ;
assign n10988 =  ( n10387 ) ? ( bv_8_232_n95 ) : ( n10987 ) ;
assign n10989 =  ( n10385 ) ? ( bv_8_221_n138 ) : ( n10988 ) ;
assign n10990 =  ( n10383 ) ? ( bv_8_116_n345 ) : ( n10989 ) ;
assign n10991 =  ( n10381 ) ? ( bv_8_31_n705 ) : ( n10990 ) ;
assign n10992 =  ( n10379 ) ? ( bv_8_75_n503 ) : ( n10991 ) ;
assign n10993 =  ( n10377 ) ? ( bv_8_189_n254 ) : ( n10992 ) ;
assign n10994 =  ( n10375 ) ? ( bv_8_139_n297 ) : ( n10993 ) ;
assign n10995 =  ( n10373 ) ? ( bv_8_138_n418 ) : ( n10994 ) ;
assign n10996 =  ( n10371 ) ? ( bv_8_112_n482 ) : ( n10995 ) ;
assign n10997 =  ( n10369 ) ? ( bv_8_62_n205 ) : ( n10996 ) ;
assign n10998 =  ( n10367 ) ? ( bv_8_181_n281 ) : ( n10997 ) ;
assign n10999 =  ( n10365 ) ? ( bv_8_102_n527 ) : ( n10998 ) ;
assign n11000 =  ( n10363 ) ? ( bv_8_72_n330 ) : ( n10999 ) ;
assign n11001 =  ( n10361 ) ? ( bv_8_3_n65 ) : ( n11000 ) ;
assign n11002 =  ( n10359 ) ? ( bv_8_246_n39 ) : ( n11001 ) ;
assign n11003 =  ( n10357 ) ? ( bv_8_14_n648 ) : ( n11002 ) ;
assign n11004 =  ( n10355 ) ? ( bv_8_97_n198 ) : ( n11003 ) ;
assign n11005 =  ( n10353 ) ? ( bv_8_53_n436 ) : ( n11004 ) ;
assign n11006 =  ( n10351 ) ? ( bv_8_87_n226 ) : ( n11005 ) ;
assign n11007 =  ( n10349 ) ? ( bv_8_185_n266 ) : ( n11006 ) ;
assign n11008 =  ( n10347 ) ? ( bv_8_134_n431 ) : ( n11007 ) ;
assign n11009 =  ( n10345 ) ? ( bv_8_193_n239 ) : ( n11008 ) ;
assign n11010 =  ( n10343 ) ? ( bv_8_29_n625 ) : ( n11009 ) ;
assign n11011 =  ( n10341 ) ? ( bv_8_158_n355 ) : ( n11010 ) ;
assign n11012 =  ( n10339 ) ? ( bv_8_225_n123 ) : ( n11011 ) ;
assign n11013 =  ( n10337 ) ? ( bv_8_248_n31 ) : ( n11012 ) ;
assign n11014 =  ( n10335 ) ? ( bv_8_152_n374 ) : ( n11013 ) ;
assign n11015 =  ( n10333 ) ? ( bv_8_17_n525 ) : ( n11014 ) ;
assign n11016 =  ( n10331 ) ? ( bv_8_105_n148 ) : ( n11015 ) ;
assign n11017 =  ( n10329 ) ? ( bv_8_217_n128 ) : ( n11016 ) ;
assign n11018 =  ( n10327 ) ? ( bv_8_142_n406 ) : ( n11017 ) ;
assign n11019 =  ( n10325 ) ? ( bv_8_148_n388 ) : ( n11018 ) ;
assign n11020 =  ( n10323 ) ? ( bv_8_155_n364 ) : ( n11019 ) ;
assign n11021 =  ( n10321 ) ? ( bv_8_30_n21 ) : ( n11020 ) ;
assign n11022 =  ( n10319 ) ? ( bv_8_135_n81 ) : ( n11021 ) ;
assign n11023 =  ( n10317 ) ? ( bv_8_233_n91 ) : ( n11022 ) ;
assign n11024 =  ( n10315 ) ? ( bv_8_206_n192 ) : ( n11023 ) ;
assign n11025 =  ( n10313 ) ? ( bv_8_85_n423 ) : ( n11024 ) ;
assign n11026 =  ( n10311 ) ? ( bv_8_40_n366 ) : ( n11025 ) ;
assign n11027 =  ( n10309 ) ? ( bv_8_223_n130 ) : ( n11026 ) ;
assign n11028 =  ( n10307 ) ? ( bv_8_140_n376 ) : ( n11027 ) ;
assign n11029 =  ( n10305 ) ? ( bv_8_161_n211 ) : ( n11028 ) ;
assign n11030 =  ( n10303 ) ? ( bv_8_137_n421 ) : ( n11029 ) ;
assign n11031 =  ( n10301 ) ? ( bv_8_13_n194 ) : ( n11030 ) ;
assign n11032 =  ( n10299 ) ? ( bv_8_191_n246 ) : ( n11031 ) ;
assign n11033 =  ( n10297 ) ? ( bv_8_230_n103 ) : ( n11032 ) ;
assign n11034 =  ( n10295 ) ? ( bv_8_66_n466 ) : ( n11033 ) ;
assign n11035 =  ( n10293 ) ? ( bv_8_104_n520 ) : ( n11034 ) ;
assign n11036 =  ( n10291 ) ? ( bv_8_65_n623 ) : ( n11035 ) ;
assign n11037 =  ( n10289 ) ? ( bv_8_153_n140 ) : ( n11036 ) ;
assign n11038 =  ( n10287 ) ? ( bv_8_45_n97 ) : ( n11037 ) ;
assign n11039 =  ( n10285 ) ? ( bv_8_15_n190 ) : ( n11038 ) ;
assign n11040 =  ( n10283 ) ? ( bv_8_176_n299 ) : ( n11039 ) ;
assign n11041 =  ( n10281 ) ? ( bv_8_84_n386 ) : ( n11040 ) ;
assign n11042 =  ( n10279 ) ? ( bv_8_187_n260 ) : ( n11041 ) ;
assign n11043 =  ( n10277 ) ? ( bv_8_22_n357 ) : ( n11042 ) ;
assign n11044 =  ( n7196 ) ^ ( n11043 )  ;
assign n11045 =  ( n11044 ) ^ ( n9502 )  ;
assign n11046 =  ( n11045 ) ^ ( n10271 )  ;
assign n11047 = state_in[15:8] ;
assign n11048 =  ( n11047 ) == ( bv_8_255_n3 )  ;
assign n11049 = state_in[15:8] ;
assign n11050 =  ( n11049 ) == ( bv_8_254_n7 )  ;
assign n11051 = state_in[15:8] ;
assign n11052 =  ( n11051 ) == ( bv_8_253_n11 )  ;
assign n11053 = state_in[15:8] ;
assign n11054 =  ( n11053 ) == ( bv_8_252_n15 )  ;
assign n11055 = state_in[15:8] ;
assign n11056 =  ( n11055 ) == ( bv_8_251_n19 )  ;
assign n11057 = state_in[15:8] ;
assign n11058 =  ( n11057 ) == ( bv_8_250_n23 )  ;
assign n11059 = state_in[15:8] ;
assign n11060 =  ( n11059 ) == ( bv_8_249_n27 )  ;
assign n11061 = state_in[15:8] ;
assign n11062 =  ( n11061 ) == ( bv_8_248_n31 )  ;
assign n11063 = state_in[15:8] ;
assign n11064 =  ( n11063 ) == ( bv_8_247_n35 )  ;
assign n11065 = state_in[15:8] ;
assign n11066 =  ( n11065 ) == ( bv_8_246_n39 )  ;
assign n11067 = state_in[15:8] ;
assign n11068 =  ( n11067 ) == ( bv_8_245_n43 )  ;
assign n11069 = state_in[15:8] ;
assign n11070 =  ( n11069 ) == ( bv_8_244_n47 )  ;
assign n11071 = state_in[15:8] ;
assign n11072 =  ( n11071 ) == ( bv_8_243_n51 )  ;
assign n11073 = state_in[15:8] ;
assign n11074 =  ( n11073 ) == ( bv_8_242_n55 )  ;
assign n11075 = state_in[15:8] ;
assign n11076 =  ( n11075 ) == ( bv_8_241_n59 )  ;
assign n11077 = state_in[15:8] ;
assign n11078 =  ( n11077 ) == ( bv_8_240_n63 )  ;
assign n11079 = state_in[15:8] ;
assign n11080 =  ( n11079 ) == ( bv_8_239_n67 )  ;
assign n11081 = state_in[15:8] ;
assign n11082 =  ( n11081 ) == ( bv_8_238_n71 )  ;
assign n11083 = state_in[15:8] ;
assign n11084 =  ( n11083 ) == ( bv_8_237_n75 )  ;
assign n11085 = state_in[15:8] ;
assign n11086 =  ( n11085 ) == ( bv_8_236_n79 )  ;
assign n11087 = state_in[15:8] ;
assign n11088 =  ( n11087 ) == ( bv_8_235_n83 )  ;
assign n11089 = state_in[15:8] ;
assign n11090 =  ( n11089 ) == ( bv_8_234_n87 )  ;
assign n11091 = state_in[15:8] ;
assign n11092 =  ( n11091 ) == ( bv_8_233_n91 )  ;
assign n11093 = state_in[15:8] ;
assign n11094 =  ( n11093 ) == ( bv_8_232_n95 )  ;
assign n11095 = state_in[15:8] ;
assign n11096 =  ( n11095 ) == ( bv_8_231_n99 )  ;
assign n11097 = state_in[15:8] ;
assign n11098 =  ( n11097 ) == ( bv_8_230_n103 )  ;
assign n11099 = state_in[15:8] ;
assign n11100 =  ( n11099 ) == ( bv_8_229_n107 )  ;
assign n11101 = state_in[15:8] ;
assign n11102 =  ( n11101 ) == ( bv_8_228_n111 )  ;
assign n11103 = state_in[15:8] ;
assign n11104 =  ( n11103 ) == ( bv_8_227_n115 )  ;
assign n11105 = state_in[15:8] ;
assign n11106 =  ( n11105 ) == ( bv_8_226_n119 )  ;
assign n11107 = state_in[15:8] ;
assign n11108 =  ( n11107 ) == ( bv_8_225_n123 )  ;
assign n11109 = state_in[15:8] ;
assign n11110 =  ( n11109 ) == ( bv_8_224_n126 )  ;
assign n11111 = state_in[15:8] ;
assign n11112 =  ( n11111 ) == ( bv_8_223_n130 )  ;
assign n11113 = state_in[15:8] ;
assign n11114 =  ( n11113 ) == ( bv_8_222_n134 )  ;
assign n11115 = state_in[15:8] ;
assign n11116 =  ( n11115 ) == ( bv_8_221_n138 )  ;
assign n11117 = state_in[15:8] ;
assign n11118 =  ( n11117 ) == ( bv_8_220_n142 )  ;
assign n11119 = state_in[15:8] ;
assign n11120 =  ( n11119 ) == ( bv_8_219_n146 )  ;
assign n11121 = state_in[15:8] ;
assign n11122 =  ( n11121 ) == ( bv_8_218_n150 )  ;
assign n11123 = state_in[15:8] ;
assign n11124 =  ( n11123 ) == ( bv_8_217_n128 )  ;
assign n11125 = state_in[15:8] ;
assign n11126 =  ( n11125 ) == ( bv_8_216_n157 )  ;
assign n11127 = state_in[15:8] ;
assign n11128 =  ( n11127 ) == ( bv_8_215_n45 )  ;
assign n11129 = state_in[15:8] ;
assign n11130 =  ( n11129 ) == ( bv_8_214_n164 )  ;
assign n11131 = state_in[15:8] ;
assign n11132 =  ( n11131 ) == ( bv_8_213_n167 )  ;
assign n11133 = state_in[15:8] ;
assign n11134 =  ( n11133 ) == ( bv_8_212_n171 )  ;
assign n11135 = state_in[15:8] ;
assign n11136 =  ( n11135 ) == ( bv_8_211_n175 )  ;
assign n11137 = state_in[15:8] ;
assign n11138 =  ( n11137 ) == ( bv_8_210_n113 )  ;
assign n11139 = state_in[15:8] ;
assign n11140 =  ( n11139 ) == ( bv_8_209_n182 )  ;
assign n11141 = state_in[15:8] ;
assign n11142 =  ( n11141 ) == ( bv_8_208_n37 )  ;
assign n11143 = state_in[15:8] ;
assign n11144 =  ( n11143 ) == ( bv_8_207_n188 )  ;
assign n11145 = state_in[15:8] ;
assign n11146 =  ( n11145 ) == ( bv_8_206_n192 )  ;
assign n11147 = state_in[15:8] ;
assign n11148 =  ( n11147 ) == ( bv_8_205_n196 )  ;
assign n11149 = state_in[15:8] ;
assign n11150 =  ( n11149 ) == ( bv_8_204_n177 )  ;
assign n11151 = state_in[15:8] ;
assign n11152 =  ( n11151 ) == ( bv_8_203_n203 )  ;
assign n11153 = state_in[15:8] ;
assign n11154 =  ( n11153 ) == ( bv_8_202_n207 )  ;
assign n11155 = state_in[15:8] ;
assign n11156 =  ( n11155 ) == ( bv_8_201_n85 )  ;
assign n11157 = state_in[15:8] ;
assign n11158 =  ( n11157 ) == ( bv_8_200_n213 )  ;
assign n11159 = state_in[15:8] ;
assign n11160 =  ( n11159 ) == ( bv_8_199_n216 )  ;
assign n11161 = state_in[15:8] ;
assign n11162 =  ( n11161 ) == ( bv_8_198_n220 )  ;
assign n11163 = state_in[15:8] ;
assign n11164 =  ( n11163 ) == ( bv_8_197_n224 )  ;
assign n11165 = state_in[15:8] ;
assign n11166 =  ( n11165 ) == ( bv_8_196_n228 )  ;
assign n11167 = state_in[15:8] ;
assign n11168 =  ( n11167 ) == ( bv_8_195_n232 )  ;
assign n11169 = state_in[15:8] ;
assign n11170 =  ( n11169 ) == ( bv_8_194_n159 )  ;
assign n11171 = state_in[15:8] ;
assign n11172 =  ( n11171 ) == ( bv_8_193_n239 )  ;
assign n11173 = state_in[15:8] ;
assign n11174 =  ( n11173 ) == ( bv_8_192_n242 )  ;
assign n11175 = state_in[15:8] ;
assign n11176 =  ( n11175 ) == ( bv_8_191_n246 )  ;
assign n11177 = state_in[15:8] ;
assign n11178 =  ( n11177 ) == ( bv_8_190_n250 )  ;
assign n11179 = state_in[15:8] ;
assign n11180 =  ( n11179 ) == ( bv_8_189_n254 )  ;
assign n11181 = state_in[15:8] ;
assign n11182 =  ( n11181 ) == ( bv_8_188_n257 )  ;
assign n11183 = state_in[15:8] ;
assign n11184 =  ( n11183 ) == ( bv_8_187_n260 )  ;
assign n11185 = state_in[15:8] ;
assign n11186 =  ( n11185 ) == ( bv_8_186_n263 )  ;
assign n11187 = state_in[15:8] ;
assign n11188 =  ( n11187 ) == ( bv_8_185_n266 )  ;
assign n11189 = state_in[15:8] ;
assign n11190 =  ( n11189 ) == ( bv_8_184_n270 )  ;
assign n11191 = state_in[15:8] ;
assign n11192 =  ( n11191 ) == ( bv_8_183_n273 )  ;
assign n11193 = state_in[15:8] ;
assign n11194 =  ( n11193 ) == ( bv_8_182_n277 )  ;
assign n11195 = state_in[15:8] ;
assign n11196 =  ( n11195 ) == ( bv_8_181_n281 )  ;
assign n11197 = state_in[15:8] ;
assign n11198 =  ( n11197 ) == ( bv_8_180_n285 )  ;
assign n11199 = state_in[15:8] ;
assign n11200 =  ( n11199 ) == ( bv_8_179_n289 )  ;
assign n11201 = state_in[15:8] ;
assign n11202 =  ( n11201 ) == ( bv_8_178_n292 )  ;
assign n11203 = state_in[15:8] ;
assign n11204 =  ( n11203 ) == ( bv_8_177_n283 )  ;
assign n11205 = state_in[15:8] ;
assign n11206 =  ( n11205 ) == ( bv_8_176_n299 )  ;
assign n11207 = state_in[15:8] ;
assign n11208 =  ( n11207 ) == ( bv_8_175_n302 )  ;
assign n11209 = state_in[15:8] ;
assign n11210 =  ( n11209 ) == ( bv_8_174_n152 )  ;
assign n11211 = state_in[15:8] ;
assign n11212 =  ( n11211 ) == ( bv_8_173_n307 )  ;
assign n11213 = state_in[15:8] ;
assign n11214 =  ( n11213 ) == ( bv_8_172_n268 )  ;
assign n11215 = state_in[15:8] ;
assign n11216 =  ( n11215 ) == ( bv_8_171_n314 )  ;
assign n11217 = state_in[15:8] ;
assign n11218 =  ( n11217 ) == ( bv_8_170_n77 )  ;
assign n11219 = state_in[15:8] ;
assign n11220 =  ( n11219 ) == ( bv_8_169_n109 )  ;
assign n11221 = state_in[15:8] ;
assign n11222 =  ( n11221 ) == ( bv_8_168_n13 )  ;
assign n11223 = state_in[15:8] ;
assign n11224 =  ( n11223 ) == ( bv_8_167_n325 )  ;
assign n11225 = state_in[15:8] ;
assign n11226 =  ( n11225 ) == ( bv_8_166_n328 )  ;
assign n11227 = state_in[15:8] ;
assign n11228 =  ( n11227 ) == ( bv_8_165_n69 )  ;
assign n11229 = state_in[15:8] ;
assign n11230 =  ( n11229 ) == ( bv_8_164_n335 )  ;
assign n11231 = state_in[15:8] ;
assign n11232 =  ( n11231 ) == ( bv_8_163_n339 )  ;
assign n11233 = state_in[15:8] ;
assign n11234 =  ( n11233 ) == ( bv_8_162_n343 )  ;
assign n11235 = state_in[15:8] ;
assign n11236 =  ( n11235 ) == ( bv_8_161_n211 )  ;
assign n11237 = state_in[15:8] ;
assign n11238 =  ( n11237 ) == ( bv_8_160_n350 )  ;
assign n11239 = state_in[15:8] ;
assign n11240 =  ( n11239 ) == ( bv_8_159_n323 )  ;
assign n11241 = state_in[15:8] ;
assign n11242 =  ( n11241 ) == ( bv_8_158_n355 )  ;
assign n11243 = state_in[15:8] ;
assign n11244 =  ( n11243 ) == ( bv_8_157_n359 )  ;
assign n11245 = state_in[15:8] ;
assign n11246 =  ( n11245 ) == ( bv_8_156_n279 )  ;
assign n11247 = state_in[15:8] ;
assign n11248 =  ( n11247 ) == ( bv_8_155_n364 )  ;
assign n11249 = state_in[15:8] ;
assign n11250 =  ( n11249 ) == ( bv_8_154_n368 )  ;
assign n11251 = state_in[15:8] ;
assign n11252 =  ( n11251 ) == ( bv_8_153_n140 )  ;
assign n11253 = state_in[15:8] ;
assign n11254 =  ( n11253 ) == ( bv_8_152_n374 )  ;
assign n11255 = state_in[15:8] ;
assign n11256 =  ( n11255 ) == ( bv_8_151_n218 )  ;
assign n11257 = state_in[15:8] ;
assign n11258 =  ( n11257 ) == ( bv_8_150_n201 )  ;
assign n11259 = state_in[15:8] ;
assign n11260 =  ( n11259 ) == ( bv_8_149_n384 )  ;
assign n11261 = state_in[15:8] ;
assign n11262 =  ( n11261 ) == ( bv_8_148_n388 )  ;
assign n11263 = state_in[15:8] ;
assign n11264 =  ( n11263 ) == ( bv_8_147_n392 )  ;
assign n11265 = state_in[15:8] ;
assign n11266 =  ( n11265 ) == ( bv_8_146_n337 )  ;
assign n11267 = state_in[15:8] ;
assign n11268 =  ( n11267 ) == ( bv_8_145_n397 )  ;
assign n11269 = state_in[15:8] ;
assign n11270 =  ( n11269 ) == ( bv_8_144_n173 )  ;
assign n11271 = state_in[15:8] ;
assign n11272 =  ( n11271 ) == ( bv_8_143_n403 )  ;
assign n11273 = state_in[15:8] ;
assign n11274 =  ( n11273 ) == ( bv_8_142_n406 )  ;
assign n11275 = state_in[15:8] ;
assign n11276 =  ( n11275 ) == ( bv_8_141_n410 )  ;
assign n11277 = state_in[15:8] ;
assign n11278 =  ( n11277 ) == ( bv_8_140_n376 )  ;
assign n11279 = state_in[15:8] ;
assign n11280 =  ( n11279 ) == ( bv_8_139_n297 )  ;
assign n11281 = state_in[15:8] ;
assign n11282 =  ( n11281 ) == ( bv_8_138_n418 )  ;
assign n11283 = state_in[15:8] ;
assign n11284 =  ( n11283 ) == ( bv_8_137_n421 )  ;
assign n11285 = state_in[15:8] ;
assign n11286 =  ( n11285 ) == ( bv_8_136_n425 )  ;
assign n11287 = state_in[15:8] ;
assign n11288 =  ( n11287 ) == ( bv_8_135_n81 )  ;
assign n11289 = state_in[15:8] ;
assign n11290 =  ( n11289 ) == ( bv_8_134_n431 )  ;
assign n11291 = state_in[15:8] ;
assign n11292 =  ( n11291 ) == ( bv_8_133_n434 )  ;
assign n11293 = state_in[15:8] ;
assign n11294 =  ( n11293 ) == ( bv_8_132_n41 )  ;
assign n11295 = state_in[15:8] ;
assign n11296 =  ( n11295 ) == ( bv_8_131_n440 )  ;
assign n11297 = state_in[15:8] ;
assign n11298 =  ( n11297 ) == ( bv_8_130_n33 )  ;
assign n11299 = state_in[15:8] ;
assign n11300 =  ( n11299 ) == ( bv_8_129_n446 )  ;
assign n11301 = state_in[15:8] ;
assign n11302 =  ( n11301 ) == ( bv_8_128_n450 )  ;
assign n11303 = state_in[15:8] ;
assign n11304 =  ( n11303 ) == ( bv_8_127_n453 )  ;
assign n11305 = state_in[15:8] ;
assign n11306 =  ( n11305 ) == ( bv_8_126_n456 )  ;
assign n11307 = state_in[15:8] ;
assign n11308 =  ( n11307 ) == ( bv_8_125_n459 )  ;
assign n11309 = state_in[15:8] ;
assign n11310 =  ( n11309 ) == ( bv_8_124_n184 )  ;
assign n11311 = state_in[15:8] ;
assign n11312 =  ( n11311 ) == ( bv_8_123_n17 )  ;
assign n11313 = state_in[15:8] ;
assign n11314 =  ( n11313 ) == ( bv_8_122_n416 )  ;
assign n11315 = state_in[15:8] ;
assign n11316 =  ( n11315 ) == ( bv_8_121_n470 )  ;
assign n11317 = state_in[15:8] ;
assign n11318 =  ( n11317 ) == ( bv_8_120_n474 )  ;
assign n11319 = state_in[15:8] ;
assign n11320 =  ( n11319 ) == ( bv_8_119_n472 )  ;
assign n11321 = state_in[15:8] ;
assign n11322 =  ( n11321 ) == ( bv_8_118_n480 )  ;
assign n11323 = state_in[15:8] ;
assign n11324 =  ( n11323 ) == ( bv_8_117_n484 )  ;
assign n11325 = state_in[15:8] ;
assign n11326 =  ( n11325 ) == ( bv_8_116_n345 )  ;
assign n11327 = state_in[15:8] ;
assign n11328 =  ( n11327 ) == ( bv_8_115_n222 )  ;
assign n11329 = state_in[15:8] ;
assign n11330 =  ( n11329 ) == ( bv_8_114_n494 )  ;
assign n11331 = state_in[15:8] ;
assign n11332 =  ( n11331 ) == ( bv_8_113_n180 )  ;
assign n11333 = state_in[15:8] ;
assign n11334 =  ( n11333 ) == ( bv_8_112_n482 )  ;
assign n11335 = state_in[15:8] ;
assign n11336 =  ( n11335 ) == ( bv_8_111_n244 )  ;
assign n11337 = state_in[15:8] ;
assign n11338 =  ( n11337 ) == ( bv_8_110_n294 )  ;
assign n11339 = state_in[15:8] ;
assign n11340 =  ( n11339 ) == ( bv_8_109_n9 )  ;
assign n11341 = state_in[15:8] ;
assign n11342 =  ( n11341 ) == ( bv_8_108_n510 )  ;
assign n11343 = state_in[15:8] ;
assign n11344 =  ( n11343 ) == ( bv_8_107_n370 )  ;
assign n11345 = state_in[15:8] ;
assign n11346 =  ( n11345 ) == ( bv_8_106_n155 )  ;
assign n11347 = state_in[15:8] ;
assign n11348 =  ( n11347 ) == ( bv_8_105_n148 )  ;
assign n11349 = state_in[15:8] ;
assign n11350 =  ( n11349 ) == ( bv_8_104_n520 )  ;
assign n11351 = state_in[15:8] ;
assign n11352 =  ( n11351 ) == ( bv_8_103_n523 )  ;
assign n11353 = state_in[15:8] ;
assign n11354 =  ( n11353 ) == ( bv_8_102_n527 )  ;
assign n11355 = state_in[15:8] ;
assign n11356 =  ( n11355 ) == ( bv_8_101_n49 )  ;
assign n11357 = state_in[15:8] ;
assign n11358 =  ( n11357 ) == ( bv_8_100_n348 )  ;
assign n11359 = state_in[15:8] ;
assign n11360 =  ( n11359 ) == ( bv_8_99_n476 )  ;
assign n11361 = state_in[15:8] ;
assign n11362 =  ( n11361 ) == ( bv_8_98_n536 )  ;
assign n11363 = state_in[15:8] ;
assign n11364 =  ( n11363 ) == ( bv_8_97_n198 )  ;
assign n11365 = state_in[15:8] ;
assign n11366 =  ( n11365 ) == ( bv_8_96_n542 )  ;
assign n11367 = state_in[15:8] ;
assign n11368 =  ( n11367 ) == ( bv_8_95_n545 )  ;
assign n11369 = state_in[15:8] ;
assign n11370 =  ( n11369 ) == ( bv_8_94_n548 )  ;
assign n11371 = state_in[15:8] ;
assign n11372 =  ( n11371 ) == ( bv_8_93_n498 )  ;
assign n11373 = state_in[15:8] ;
assign n11374 =  ( n11373 ) == ( bv_8_92_n234 )  ;
assign n11375 = state_in[15:8] ;
assign n11376 =  ( n11375 ) == ( bv_8_91_n555 )  ;
assign n11377 = state_in[15:8] ;
assign n11378 =  ( n11377 ) == ( bv_8_90_n25 )  ;
assign n11379 = state_in[15:8] ;
assign n11380 =  ( n11379 ) == ( bv_8_89_n61 )  ;
assign n11381 = state_in[15:8] ;
assign n11382 =  ( n11381 ) == ( bv_8_88_n562 )  ;
assign n11383 = state_in[15:8] ;
assign n11384 =  ( n11383 ) == ( bv_8_87_n226 )  ;
assign n11385 = state_in[15:8] ;
assign n11386 =  ( n11385 ) == ( bv_8_86_n567 )  ;
assign n11387 = state_in[15:8] ;
assign n11388 =  ( n11387 ) == ( bv_8_85_n423 )  ;
assign n11389 = state_in[15:8] ;
assign n11390 =  ( n11389 ) == ( bv_8_84_n386 )  ;
assign n11391 = state_in[15:8] ;
assign n11392 =  ( n11391 ) == ( bv_8_83_n575 )  ;
assign n11393 = state_in[15:8] ;
assign n11394 =  ( n11393 ) == ( bv_8_82_n578 )  ;
assign n11395 = state_in[15:8] ;
assign n11396 =  ( n11395 ) == ( bv_8_81_n582 )  ;
assign n11397 = state_in[15:8] ;
assign n11398 =  ( n11397 ) == ( bv_8_80_n73 )  ;
assign n11399 = state_in[15:8] ;
assign n11400 =  ( n11399 ) == ( bv_8_79_n538 )  ;
assign n11401 = state_in[15:8] ;
assign n11402 =  ( n11401 ) == ( bv_8_78_n590 )  ;
assign n11403 = state_in[15:8] ;
assign n11404 =  ( n11403 ) == ( bv_8_77_n593 )  ;
assign n11405 = state_in[15:8] ;
assign n11406 =  ( n11405 ) == ( bv_8_76_n596 )  ;
assign n11407 = state_in[15:8] ;
assign n11408 =  ( n11407 ) == ( bv_8_75_n503 )  ;
assign n11409 = state_in[15:8] ;
assign n11410 =  ( n11409 ) == ( bv_8_74_n237 )  ;
assign n11411 = state_in[15:8] ;
assign n11412 =  ( n11411 ) == ( bv_8_73_n275 )  ;
assign n11413 = state_in[15:8] ;
assign n11414 =  ( n11413 ) == ( bv_8_72_n330 )  ;
assign n11415 = state_in[15:8] ;
assign n11416 =  ( n11415 ) == ( bv_8_71_n252 )  ;
assign n11417 = state_in[15:8] ;
assign n11418 =  ( n11417 ) == ( bv_8_70_n609 )  ;
assign n11419 = state_in[15:8] ;
assign n11420 =  ( n11419 ) == ( bv_8_69_n612 )  ;
assign n11421 = state_in[15:8] ;
assign n11422 =  ( n11421 ) == ( bv_8_68_n390 )  ;
assign n11423 = state_in[15:8] ;
assign n11424 =  ( n11423 ) == ( bv_8_67_n318 )  ;
assign n11425 = state_in[15:8] ;
assign n11426 =  ( n11425 ) == ( bv_8_66_n466 )  ;
assign n11427 = state_in[15:8] ;
assign n11428 =  ( n11427 ) == ( bv_8_65_n623 )  ;
assign n11429 = state_in[15:8] ;
assign n11430 =  ( n11429 ) == ( bv_8_64_n573 )  ;
assign n11431 = state_in[15:8] ;
assign n11432 =  ( n11431 ) == ( bv_8_63_n489 )  ;
assign n11433 = state_in[15:8] ;
assign n11434 =  ( n11433 ) == ( bv_8_62_n205 )  ;
assign n11435 = state_in[15:8] ;
assign n11436 =  ( n11435 ) == ( bv_8_61_n634 )  ;
assign n11437 = state_in[15:8] ;
assign n11438 =  ( n11437 ) == ( bv_8_60_n93 )  ;
assign n11439 = state_in[15:8] ;
assign n11440 =  ( n11439 ) == ( bv_8_59_n382 )  ;
assign n11441 = state_in[15:8] ;
assign n11442 =  ( n11441 ) == ( bv_8_58_n136 )  ;
assign n11443 = state_in[15:8] ;
assign n11444 =  ( n11443 ) == ( bv_8_57_n312 )  ;
assign n11445 = state_in[15:8] ;
assign n11446 =  ( n11445 ) == ( bv_8_56_n230 )  ;
assign n11447 = state_in[15:8] ;
assign n11448 =  ( n11447 ) == ( bv_8_55_n650 )  ;
assign n11449 = state_in[15:8] ;
assign n11450 =  ( n11449 ) == ( bv_8_54_n616 )  ;
assign n11451 = state_in[15:8] ;
assign n11452 =  ( n11451 ) == ( bv_8_53_n436 )  ;
assign n11453 = state_in[15:8] ;
assign n11454 =  ( n11453 ) == ( bv_8_52_n619 )  ;
assign n11455 = state_in[15:8] ;
assign n11456 =  ( n11455 ) == ( bv_8_51_n101 )  ;
assign n11457 = state_in[15:8] ;
assign n11458 =  ( n11457 ) == ( bv_8_50_n408 )  ;
assign n11459 = state_in[15:8] ;
assign n11460 =  ( n11459 ) == ( bv_8_49_n309 )  ;
assign n11461 = state_in[15:8] ;
assign n11462 =  ( n11461 ) == ( bv_8_48_n660 )  ;
assign n11463 = state_in[15:8] ;
assign n11464 =  ( n11463 ) == ( bv_8_47_n652 )  ;
assign n11465 = state_in[15:8] ;
assign n11466 =  ( n11465 ) == ( bv_8_46_n429 )  ;
assign n11467 = state_in[15:8] ;
assign n11468 =  ( n11467 ) == ( bv_8_45_n97 )  ;
assign n11469 = state_in[15:8] ;
assign n11470 =  ( n11469 ) == ( bv_8_44_n5 )  ;
assign n11471 = state_in[15:8] ;
assign n11472 =  ( n11471 ) == ( bv_8_43_n121 )  ;
assign n11473 = state_in[15:8] ;
assign n11474 =  ( n11473 ) == ( bv_8_42_n672 )  ;
assign n11475 = state_in[15:8] ;
assign n11476 =  ( n11475 ) == ( bv_8_41_n29 )  ;
assign n11477 = state_in[15:8] ;
assign n11478 =  ( n11477 ) == ( bv_8_40_n366 )  ;
assign n11479 = state_in[15:8] ;
assign n11480 =  ( n11479 ) == ( bv_8_39_n132 )  ;
assign n11481 = state_in[15:8] ;
assign n11482 =  ( n11481 ) == ( bv_8_38_n444 )  ;
assign n11483 = state_in[15:8] ;
assign n11484 =  ( n11483 ) == ( bv_8_37_n506 )  ;
assign n11485 = state_in[15:8] ;
assign n11486 =  ( n11485 ) == ( bv_8_36_n645 )  ;
assign n11487 = state_in[15:8] ;
assign n11488 =  ( n11487 ) == ( bv_8_35_n696 )  ;
assign n11489 = state_in[15:8] ;
assign n11490 =  ( n11489 ) == ( bv_8_34_n117 )  ;
assign n11491 = state_in[15:8] ;
assign n11492 =  ( n11491 ) == ( bv_8_33_n486 )  ;
assign n11493 = state_in[15:8] ;
assign n11494 =  ( n11493 ) == ( bv_8_32_n463 )  ;
assign n11495 = state_in[15:8] ;
assign n11496 =  ( n11495 ) == ( bv_8_31_n705 )  ;
assign n11497 = state_in[15:8] ;
assign n11498 =  ( n11497 ) == ( bv_8_30_n21 )  ;
assign n11499 = state_in[15:8] ;
assign n11500 =  ( n11499 ) == ( bv_8_29_n625 )  ;
assign n11501 = state_in[15:8] ;
assign n11502 =  ( n11501 ) == ( bv_8_28_n162 )  ;
assign n11503 = state_in[15:8] ;
assign n11504 =  ( n11503 ) == ( bv_8_27_n642 )  ;
assign n11505 = state_in[15:8] ;
assign n11506 =  ( n11505 ) == ( bv_8_26_n53 )  ;
assign n11507 = state_in[15:8] ;
assign n11508 =  ( n11507 ) == ( bv_8_25_n399 )  ;
assign n11509 = state_in[15:8] ;
assign n11510 =  ( n11509 ) == ( bv_8_24_n448 )  ;
assign n11511 = state_in[15:8] ;
assign n11512 =  ( n11511 ) == ( bv_8_23_n144 )  ;
assign n11513 = state_in[15:8] ;
assign n11514 =  ( n11513 ) == ( bv_8_22_n357 )  ;
assign n11515 = state_in[15:8] ;
assign n11516 =  ( n11515 ) == ( bv_8_21_n89 )  ;
assign n11517 = state_in[15:8] ;
assign n11518 =  ( n11517 ) == ( bv_8_20_n341 )  ;
assign n11519 = state_in[15:8] ;
assign n11520 =  ( n11519 ) == ( bv_8_19_n588 )  ;
assign n11521 = state_in[15:8] ;
assign n11522 =  ( n11521 ) == ( bv_8_18_n628 )  ;
assign n11523 = state_in[15:8] ;
assign n11524 =  ( n11523 ) == ( bv_8_17_n525 )  ;
assign n11525 = state_in[15:8] ;
assign n11526 =  ( n11525 ) == ( bv_8_16_n248 )  ;
assign n11527 = state_in[15:8] ;
assign n11528 =  ( n11527 ) == ( bv_8_15_n190 )  ;
assign n11529 = state_in[15:8] ;
assign n11530 =  ( n11529 ) == ( bv_8_14_n648 )  ;
assign n11531 = state_in[15:8] ;
assign n11532 =  ( n11531 ) == ( bv_8_13_n194 )  ;
assign n11533 = state_in[15:8] ;
assign n11534 =  ( n11533 ) == ( bv_8_12_n333 )  ;
assign n11535 = state_in[15:8] ;
assign n11536 =  ( n11535 ) == ( bv_8_11_n379 )  ;
assign n11537 = state_in[15:8] ;
assign n11538 =  ( n11537 ) == ( bv_8_10_n655 )  ;
assign n11539 = state_in[15:8] ;
assign n11540 =  ( n11539 ) == ( bv_8_9_n57 )  ;
assign n11541 = state_in[15:8] ;
assign n11542 =  ( n11541 ) == ( bv_8_8_n669 )  ;
assign n11543 = state_in[15:8] ;
assign n11544 =  ( n11543 ) == ( bv_8_7_n105 )  ;
assign n11545 = state_in[15:8] ;
assign n11546 =  ( n11545 ) == ( bv_8_6_n169 )  ;
assign n11547 = state_in[15:8] ;
assign n11548 =  ( n11547 ) == ( bv_8_5_n492 )  ;
assign n11549 = state_in[15:8] ;
assign n11550 =  ( n11549 ) == ( bv_8_4_n516 )  ;
assign n11551 = state_in[15:8] ;
assign n11552 =  ( n11551 ) == ( bv_8_3_n65 )  ;
assign n11553 = state_in[15:8] ;
assign n11554 =  ( n11553 ) == ( bv_8_2_n751 )  ;
assign n11555 = state_in[15:8] ;
assign n11556 =  ( n11555 ) == ( bv_8_1_n287 )  ;
assign n11557 = state_in[15:8] ;
assign n11558 =  ( n11557 ) == ( bv_8_0_n580 )  ;
assign n11559 =  ( n11558 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n11560 =  ( n11556 ) ? ( bv_8_248_n31 ) : ( n11559 ) ;
assign n11561 =  ( n11554 ) ? ( bv_8_238_n71 ) : ( n11560 ) ;
assign n11562 =  ( n11552 ) ? ( bv_8_246_n39 ) : ( n11561 ) ;
assign n11563 =  ( n11550 ) ? ( bv_8_255_n3 ) : ( n11562 ) ;
assign n11564 =  ( n11548 ) ? ( bv_8_214_n164 ) : ( n11563 ) ;
assign n11565 =  ( n11546 ) ? ( bv_8_222_n134 ) : ( n11564 ) ;
assign n11566 =  ( n11544 ) ? ( bv_8_145_n397 ) : ( n11565 ) ;
assign n11567 =  ( n11542 ) ? ( bv_8_96_n542 ) : ( n11566 ) ;
assign n11568 =  ( n11540 ) ? ( bv_8_2_n751 ) : ( n11567 ) ;
assign n11569 =  ( n11538 ) ? ( bv_8_206_n192 ) : ( n11568 ) ;
assign n11570 =  ( n11536 ) ? ( bv_8_86_n567 ) : ( n11569 ) ;
assign n11571 =  ( n11534 ) ? ( bv_8_231_n99 ) : ( n11570 ) ;
assign n11572 =  ( n11532 ) ? ( bv_8_181_n281 ) : ( n11571 ) ;
assign n11573 =  ( n11530 ) ? ( bv_8_77_n593 ) : ( n11572 ) ;
assign n11574 =  ( n11528 ) ? ( bv_8_236_n79 ) : ( n11573 ) ;
assign n11575 =  ( n11526 ) ? ( bv_8_143_n403 ) : ( n11574 ) ;
assign n11576 =  ( n11524 ) ? ( bv_8_31_n705 ) : ( n11575 ) ;
assign n11577 =  ( n11522 ) ? ( bv_8_137_n421 ) : ( n11576 ) ;
assign n11578 =  ( n11520 ) ? ( bv_8_250_n23 ) : ( n11577 ) ;
assign n11579 =  ( n11518 ) ? ( bv_8_239_n67 ) : ( n11578 ) ;
assign n11580 =  ( n11516 ) ? ( bv_8_178_n292 ) : ( n11579 ) ;
assign n11581 =  ( n11514 ) ? ( bv_8_142_n406 ) : ( n11580 ) ;
assign n11582 =  ( n11512 ) ? ( bv_8_251_n19 ) : ( n11581 ) ;
assign n11583 =  ( n11510 ) ? ( bv_8_65_n623 ) : ( n11582 ) ;
assign n11584 =  ( n11508 ) ? ( bv_8_179_n289 ) : ( n11583 ) ;
assign n11585 =  ( n11506 ) ? ( bv_8_95_n545 ) : ( n11584 ) ;
assign n11586 =  ( n11504 ) ? ( bv_8_69_n612 ) : ( n11585 ) ;
assign n11587 =  ( n11502 ) ? ( bv_8_35_n696 ) : ( n11586 ) ;
assign n11588 =  ( n11500 ) ? ( bv_8_83_n575 ) : ( n11587 ) ;
assign n11589 =  ( n11498 ) ? ( bv_8_228_n111 ) : ( n11588 ) ;
assign n11590 =  ( n11496 ) ? ( bv_8_155_n364 ) : ( n11589 ) ;
assign n11591 =  ( n11494 ) ? ( bv_8_117_n484 ) : ( n11590 ) ;
assign n11592 =  ( n11492 ) ? ( bv_8_225_n123 ) : ( n11591 ) ;
assign n11593 =  ( n11490 ) ? ( bv_8_61_n634 ) : ( n11592 ) ;
assign n11594 =  ( n11488 ) ? ( bv_8_76_n596 ) : ( n11593 ) ;
assign n11595 =  ( n11486 ) ? ( bv_8_108_n510 ) : ( n11594 ) ;
assign n11596 =  ( n11484 ) ? ( bv_8_126_n456 ) : ( n11595 ) ;
assign n11597 =  ( n11482 ) ? ( bv_8_245_n43 ) : ( n11596 ) ;
assign n11598 =  ( n11480 ) ? ( bv_8_131_n440 ) : ( n11597 ) ;
assign n11599 =  ( n11478 ) ? ( bv_8_104_n520 ) : ( n11598 ) ;
assign n11600 =  ( n11476 ) ? ( bv_8_81_n582 ) : ( n11599 ) ;
assign n11601 =  ( n11474 ) ? ( bv_8_209_n182 ) : ( n11600 ) ;
assign n11602 =  ( n11472 ) ? ( bv_8_249_n27 ) : ( n11601 ) ;
assign n11603 =  ( n11470 ) ? ( bv_8_226_n119 ) : ( n11602 ) ;
assign n11604 =  ( n11468 ) ? ( bv_8_171_n314 ) : ( n11603 ) ;
assign n11605 =  ( n11466 ) ? ( bv_8_98_n536 ) : ( n11604 ) ;
assign n11606 =  ( n11464 ) ? ( bv_8_42_n672 ) : ( n11605 ) ;
assign n11607 =  ( n11462 ) ? ( bv_8_8_n669 ) : ( n11606 ) ;
assign n11608 =  ( n11460 ) ? ( bv_8_149_n384 ) : ( n11607 ) ;
assign n11609 =  ( n11458 ) ? ( bv_8_70_n609 ) : ( n11608 ) ;
assign n11610 =  ( n11456 ) ? ( bv_8_157_n359 ) : ( n11609 ) ;
assign n11611 =  ( n11454 ) ? ( bv_8_48_n660 ) : ( n11610 ) ;
assign n11612 =  ( n11452 ) ? ( bv_8_55_n650 ) : ( n11611 ) ;
assign n11613 =  ( n11450 ) ? ( bv_8_10_n655 ) : ( n11612 ) ;
assign n11614 =  ( n11448 ) ? ( bv_8_47_n652 ) : ( n11613 ) ;
assign n11615 =  ( n11446 ) ? ( bv_8_14_n648 ) : ( n11614 ) ;
assign n11616 =  ( n11444 ) ? ( bv_8_36_n645 ) : ( n11615 ) ;
assign n11617 =  ( n11442 ) ? ( bv_8_27_n642 ) : ( n11616 ) ;
assign n11618 =  ( n11440 ) ? ( bv_8_223_n130 ) : ( n11617 ) ;
assign n11619 =  ( n11438 ) ? ( bv_8_205_n196 ) : ( n11618 ) ;
assign n11620 =  ( n11436 ) ? ( bv_8_78_n590 ) : ( n11619 ) ;
assign n11621 =  ( n11434 ) ? ( bv_8_127_n453 ) : ( n11620 ) ;
assign n11622 =  ( n11432 ) ? ( bv_8_234_n87 ) : ( n11621 ) ;
assign n11623 =  ( n11430 ) ? ( bv_8_18_n628 ) : ( n11622 ) ;
assign n11624 =  ( n11428 ) ? ( bv_8_29_n625 ) : ( n11623 ) ;
assign n11625 =  ( n11426 ) ? ( bv_8_88_n562 ) : ( n11624 ) ;
assign n11626 =  ( n11424 ) ? ( bv_8_52_n619 ) : ( n11625 ) ;
assign n11627 =  ( n11422 ) ? ( bv_8_54_n616 ) : ( n11626 ) ;
assign n11628 =  ( n11420 ) ? ( bv_8_220_n142 ) : ( n11627 ) ;
assign n11629 =  ( n11418 ) ? ( bv_8_180_n285 ) : ( n11628 ) ;
assign n11630 =  ( n11416 ) ? ( bv_8_91_n555 ) : ( n11629 ) ;
assign n11631 =  ( n11414 ) ? ( bv_8_164_n335 ) : ( n11630 ) ;
assign n11632 =  ( n11412 ) ? ( bv_8_118_n480 ) : ( n11631 ) ;
assign n11633 =  ( n11410 ) ? ( bv_8_183_n273 ) : ( n11632 ) ;
assign n11634 =  ( n11408 ) ? ( bv_8_125_n459 ) : ( n11633 ) ;
assign n11635 =  ( n11406 ) ? ( bv_8_82_n578 ) : ( n11634 ) ;
assign n11636 =  ( n11404 ) ? ( bv_8_221_n138 ) : ( n11635 ) ;
assign n11637 =  ( n11402 ) ? ( bv_8_94_n548 ) : ( n11636 ) ;
assign n11638 =  ( n11400 ) ? ( bv_8_19_n588 ) : ( n11637 ) ;
assign n11639 =  ( n11398 ) ? ( bv_8_166_n328 ) : ( n11638 ) ;
assign n11640 =  ( n11396 ) ? ( bv_8_185_n266 ) : ( n11639 ) ;
assign n11641 =  ( n11394 ) ? ( bv_8_0_n580 ) : ( n11640 ) ;
assign n11642 =  ( n11392 ) ? ( bv_8_193_n239 ) : ( n11641 ) ;
assign n11643 =  ( n11390 ) ? ( bv_8_64_n573 ) : ( n11642 ) ;
assign n11644 =  ( n11388 ) ? ( bv_8_227_n115 ) : ( n11643 ) ;
assign n11645 =  ( n11386 ) ? ( bv_8_121_n470 ) : ( n11644 ) ;
assign n11646 =  ( n11384 ) ? ( bv_8_182_n277 ) : ( n11645 ) ;
assign n11647 =  ( n11382 ) ? ( bv_8_212_n171 ) : ( n11646 ) ;
assign n11648 =  ( n11380 ) ? ( bv_8_141_n410 ) : ( n11647 ) ;
assign n11649 =  ( n11378 ) ? ( bv_8_103_n523 ) : ( n11648 ) ;
assign n11650 =  ( n11376 ) ? ( bv_8_114_n494 ) : ( n11649 ) ;
assign n11651 =  ( n11374 ) ? ( bv_8_148_n388 ) : ( n11650 ) ;
assign n11652 =  ( n11372 ) ? ( bv_8_152_n374 ) : ( n11651 ) ;
assign n11653 =  ( n11370 ) ? ( bv_8_176_n299 ) : ( n11652 ) ;
assign n11654 =  ( n11368 ) ? ( bv_8_133_n434 ) : ( n11653 ) ;
assign n11655 =  ( n11366 ) ? ( bv_8_187_n260 ) : ( n11654 ) ;
assign n11656 =  ( n11364 ) ? ( bv_8_197_n224 ) : ( n11655 ) ;
assign n11657 =  ( n11362 ) ? ( bv_8_79_n538 ) : ( n11656 ) ;
assign n11658 =  ( n11360 ) ? ( bv_8_237_n75 ) : ( n11657 ) ;
assign n11659 =  ( n11358 ) ? ( bv_8_134_n431 ) : ( n11658 ) ;
assign n11660 =  ( n11356 ) ? ( bv_8_154_n368 ) : ( n11659 ) ;
assign n11661 =  ( n11354 ) ? ( bv_8_102_n527 ) : ( n11660 ) ;
assign n11662 =  ( n11352 ) ? ( bv_8_17_n525 ) : ( n11661 ) ;
assign n11663 =  ( n11350 ) ? ( bv_8_138_n418 ) : ( n11662 ) ;
assign n11664 =  ( n11348 ) ? ( bv_8_233_n91 ) : ( n11663 ) ;
assign n11665 =  ( n11346 ) ? ( bv_8_4_n516 ) : ( n11664 ) ;
assign n11666 =  ( n11344 ) ? ( bv_8_254_n7 ) : ( n11665 ) ;
assign n11667 =  ( n11342 ) ? ( bv_8_160_n350 ) : ( n11666 ) ;
assign n11668 =  ( n11340 ) ? ( bv_8_120_n474 ) : ( n11667 ) ;
assign n11669 =  ( n11338 ) ? ( bv_8_37_n506 ) : ( n11668 ) ;
assign n11670 =  ( n11336 ) ? ( bv_8_75_n503 ) : ( n11669 ) ;
assign n11671 =  ( n11334 ) ? ( bv_8_162_n343 ) : ( n11670 ) ;
assign n11672 =  ( n11332 ) ? ( bv_8_93_n498 ) : ( n11671 ) ;
assign n11673 =  ( n11330 ) ? ( bv_8_128_n450 ) : ( n11672 ) ;
assign n11674 =  ( n11328 ) ? ( bv_8_5_n492 ) : ( n11673 ) ;
assign n11675 =  ( n11326 ) ? ( bv_8_63_n489 ) : ( n11674 ) ;
assign n11676 =  ( n11324 ) ? ( bv_8_33_n486 ) : ( n11675 ) ;
assign n11677 =  ( n11322 ) ? ( bv_8_112_n482 ) : ( n11676 ) ;
assign n11678 =  ( n11320 ) ? ( bv_8_241_n59 ) : ( n11677 ) ;
assign n11679 =  ( n11318 ) ? ( bv_8_99_n476 ) : ( n11678 ) ;
assign n11680 =  ( n11316 ) ? ( bv_8_119_n472 ) : ( n11679 ) ;
assign n11681 =  ( n11314 ) ? ( bv_8_175_n302 ) : ( n11680 ) ;
assign n11682 =  ( n11312 ) ? ( bv_8_66_n466 ) : ( n11681 ) ;
assign n11683 =  ( n11310 ) ? ( bv_8_32_n463 ) : ( n11682 ) ;
assign n11684 =  ( n11308 ) ? ( bv_8_229_n107 ) : ( n11683 ) ;
assign n11685 =  ( n11306 ) ? ( bv_8_253_n11 ) : ( n11684 ) ;
assign n11686 =  ( n11304 ) ? ( bv_8_191_n246 ) : ( n11685 ) ;
assign n11687 =  ( n11302 ) ? ( bv_8_129_n446 ) : ( n11686 ) ;
assign n11688 =  ( n11300 ) ? ( bv_8_24_n448 ) : ( n11687 ) ;
assign n11689 =  ( n11298 ) ? ( bv_8_38_n444 ) : ( n11688 ) ;
assign n11690 =  ( n11296 ) ? ( bv_8_195_n232 ) : ( n11689 ) ;
assign n11691 =  ( n11294 ) ? ( bv_8_190_n250 ) : ( n11690 ) ;
assign n11692 =  ( n11292 ) ? ( bv_8_53_n436 ) : ( n11691 ) ;
assign n11693 =  ( n11290 ) ? ( bv_8_136_n425 ) : ( n11692 ) ;
assign n11694 =  ( n11288 ) ? ( bv_8_46_n429 ) : ( n11693 ) ;
assign n11695 =  ( n11286 ) ? ( bv_8_147_n392 ) : ( n11694 ) ;
assign n11696 =  ( n11284 ) ? ( bv_8_85_n423 ) : ( n11695 ) ;
assign n11697 =  ( n11282 ) ? ( bv_8_252_n15 ) : ( n11696 ) ;
assign n11698 =  ( n11280 ) ? ( bv_8_122_n416 ) : ( n11697 ) ;
assign n11699 =  ( n11278 ) ? ( bv_8_200_n213 ) : ( n11698 ) ;
assign n11700 =  ( n11276 ) ? ( bv_8_186_n263 ) : ( n11699 ) ;
assign n11701 =  ( n11274 ) ? ( bv_8_50_n408 ) : ( n11700 ) ;
assign n11702 =  ( n11272 ) ? ( bv_8_230_n103 ) : ( n11701 ) ;
assign n11703 =  ( n11270 ) ? ( bv_8_192_n242 ) : ( n11702 ) ;
assign n11704 =  ( n11268 ) ? ( bv_8_25_n399 ) : ( n11703 ) ;
assign n11705 =  ( n11266 ) ? ( bv_8_158_n355 ) : ( n11704 ) ;
assign n11706 =  ( n11264 ) ? ( bv_8_163_n339 ) : ( n11705 ) ;
assign n11707 =  ( n11262 ) ? ( bv_8_68_n390 ) : ( n11706 ) ;
assign n11708 =  ( n11260 ) ? ( bv_8_84_n386 ) : ( n11707 ) ;
assign n11709 =  ( n11258 ) ? ( bv_8_59_n382 ) : ( n11708 ) ;
assign n11710 =  ( n11256 ) ? ( bv_8_11_n379 ) : ( n11709 ) ;
assign n11711 =  ( n11254 ) ? ( bv_8_140_n376 ) : ( n11710 ) ;
assign n11712 =  ( n11252 ) ? ( bv_8_199_n216 ) : ( n11711 ) ;
assign n11713 =  ( n11250 ) ? ( bv_8_107_n370 ) : ( n11712 ) ;
assign n11714 =  ( n11248 ) ? ( bv_8_40_n366 ) : ( n11713 ) ;
assign n11715 =  ( n11246 ) ? ( bv_8_167_n325 ) : ( n11714 ) ;
assign n11716 =  ( n11244 ) ? ( bv_8_188_n257 ) : ( n11715 ) ;
assign n11717 =  ( n11242 ) ? ( bv_8_22_n357 ) : ( n11716 ) ;
assign n11718 =  ( n11240 ) ? ( bv_8_173_n307 ) : ( n11717 ) ;
assign n11719 =  ( n11238 ) ? ( bv_8_219_n146 ) : ( n11718 ) ;
assign n11720 =  ( n11236 ) ? ( bv_8_100_n348 ) : ( n11719 ) ;
assign n11721 =  ( n11234 ) ? ( bv_8_116_n345 ) : ( n11720 ) ;
assign n11722 =  ( n11232 ) ? ( bv_8_20_n341 ) : ( n11721 ) ;
assign n11723 =  ( n11230 ) ? ( bv_8_146_n337 ) : ( n11722 ) ;
assign n11724 =  ( n11228 ) ? ( bv_8_12_n333 ) : ( n11723 ) ;
assign n11725 =  ( n11226 ) ? ( bv_8_72_n330 ) : ( n11724 ) ;
assign n11726 =  ( n11224 ) ? ( bv_8_184_n270 ) : ( n11725 ) ;
assign n11727 =  ( n11222 ) ? ( bv_8_159_n323 ) : ( n11726 ) ;
assign n11728 =  ( n11220 ) ? ( bv_8_189_n254 ) : ( n11727 ) ;
assign n11729 =  ( n11218 ) ? ( bv_8_67_n318 ) : ( n11728 ) ;
assign n11730 =  ( n11216 ) ? ( bv_8_196_n228 ) : ( n11729 ) ;
assign n11731 =  ( n11214 ) ? ( bv_8_57_n312 ) : ( n11730 ) ;
assign n11732 =  ( n11212 ) ? ( bv_8_49_n309 ) : ( n11731 ) ;
assign n11733 =  ( n11210 ) ? ( bv_8_211_n175 ) : ( n11732 ) ;
assign n11734 =  ( n11208 ) ? ( bv_8_242_n55 ) : ( n11733 ) ;
assign n11735 =  ( n11206 ) ? ( bv_8_213_n167 ) : ( n11734 ) ;
assign n11736 =  ( n11204 ) ? ( bv_8_139_n297 ) : ( n11735 ) ;
assign n11737 =  ( n11202 ) ? ( bv_8_110_n294 ) : ( n11736 ) ;
assign n11738 =  ( n11200 ) ? ( bv_8_218_n150 ) : ( n11737 ) ;
assign n11739 =  ( n11198 ) ? ( bv_8_1_n287 ) : ( n11738 ) ;
assign n11740 =  ( n11196 ) ? ( bv_8_177_n283 ) : ( n11739 ) ;
assign n11741 =  ( n11194 ) ? ( bv_8_156_n279 ) : ( n11740 ) ;
assign n11742 =  ( n11192 ) ? ( bv_8_73_n275 ) : ( n11741 ) ;
assign n11743 =  ( n11190 ) ? ( bv_8_216_n157 ) : ( n11742 ) ;
assign n11744 =  ( n11188 ) ? ( bv_8_172_n268 ) : ( n11743 ) ;
assign n11745 =  ( n11186 ) ? ( bv_8_243_n51 ) : ( n11744 ) ;
assign n11746 =  ( n11184 ) ? ( bv_8_207_n188 ) : ( n11745 ) ;
assign n11747 =  ( n11182 ) ? ( bv_8_202_n207 ) : ( n11746 ) ;
assign n11748 =  ( n11180 ) ? ( bv_8_244_n47 ) : ( n11747 ) ;
assign n11749 =  ( n11178 ) ? ( bv_8_71_n252 ) : ( n11748 ) ;
assign n11750 =  ( n11176 ) ? ( bv_8_16_n248 ) : ( n11749 ) ;
assign n11751 =  ( n11174 ) ? ( bv_8_111_n244 ) : ( n11750 ) ;
assign n11752 =  ( n11172 ) ? ( bv_8_240_n63 ) : ( n11751 ) ;
assign n11753 =  ( n11170 ) ? ( bv_8_74_n237 ) : ( n11752 ) ;
assign n11754 =  ( n11168 ) ? ( bv_8_92_n234 ) : ( n11753 ) ;
assign n11755 =  ( n11166 ) ? ( bv_8_56_n230 ) : ( n11754 ) ;
assign n11756 =  ( n11164 ) ? ( bv_8_87_n226 ) : ( n11755 ) ;
assign n11757 =  ( n11162 ) ? ( bv_8_115_n222 ) : ( n11756 ) ;
assign n11758 =  ( n11160 ) ? ( bv_8_151_n218 ) : ( n11757 ) ;
assign n11759 =  ( n11158 ) ? ( bv_8_203_n203 ) : ( n11758 ) ;
assign n11760 =  ( n11156 ) ? ( bv_8_161_n211 ) : ( n11759 ) ;
assign n11761 =  ( n11154 ) ? ( bv_8_232_n95 ) : ( n11760 ) ;
assign n11762 =  ( n11152 ) ? ( bv_8_62_n205 ) : ( n11761 ) ;
assign n11763 =  ( n11150 ) ? ( bv_8_150_n201 ) : ( n11762 ) ;
assign n11764 =  ( n11148 ) ? ( bv_8_97_n198 ) : ( n11763 ) ;
assign n11765 =  ( n11146 ) ? ( bv_8_13_n194 ) : ( n11764 ) ;
assign n11766 =  ( n11144 ) ? ( bv_8_15_n190 ) : ( n11765 ) ;
assign n11767 =  ( n11142 ) ? ( bv_8_224_n126 ) : ( n11766 ) ;
assign n11768 =  ( n11140 ) ? ( bv_8_124_n184 ) : ( n11767 ) ;
assign n11769 =  ( n11138 ) ? ( bv_8_113_n180 ) : ( n11768 ) ;
assign n11770 =  ( n11136 ) ? ( bv_8_204_n177 ) : ( n11769 ) ;
assign n11771 =  ( n11134 ) ? ( bv_8_144_n173 ) : ( n11770 ) ;
assign n11772 =  ( n11132 ) ? ( bv_8_6_n169 ) : ( n11771 ) ;
assign n11773 =  ( n11130 ) ? ( bv_8_247_n35 ) : ( n11772 ) ;
assign n11774 =  ( n11128 ) ? ( bv_8_28_n162 ) : ( n11773 ) ;
assign n11775 =  ( n11126 ) ? ( bv_8_194_n159 ) : ( n11774 ) ;
assign n11776 =  ( n11124 ) ? ( bv_8_106_n155 ) : ( n11775 ) ;
assign n11777 =  ( n11122 ) ? ( bv_8_174_n152 ) : ( n11776 ) ;
assign n11778 =  ( n11120 ) ? ( bv_8_105_n148 ) : ( n11777 ) ;
assign n11779 =  ( n11118 ) ? ( bv_8_23_n144 ) : ( n11778 ) ;
assign n11780 =  ( n11116 ) ? ( bv_8_153_n140 ) : ( n11779 ) ;
assign n11781 =  ( n11114 ) ? ( bv_8_58_n136 ) : ( n11780 ) ;
assign n11782 =  ( n11112 ) ? ( bv_8_39_n132 ) : ( n11781 ) ;
assign n11783 =  ( n11110 ) ? ( bv_8_217_n128 ) : ( n11782 ) ;
assign n11784 =  ( n11108 ) ? ( bv_8_235_n83 ) : ( n11783 ) ;
assign n11785 =  ( n11106 ) ? ( bv_8_43_n121 ) : ( n11784 ) ;
assign n11786 =  ( n11104 ) ? ( bv_8_34_n117 ) : ( n11785 ) ;
assign n11787 =  ( n11102 ) ? ( bv_8_210_n113 ) : ( n11786 ) ;
assign n11788 =  ( n11100 ) ? ( bv_8_169_n109 ) : ( n11787 ) ;
assign n11789 =  ( n11098 ) ? ( bv_8_7_n105 ) : ( n11788 ) ;
assign n11790 =  ( n11096 ) ? ( bv_8_51_n101 ) : ( n11789 ) ;
assign n11791 =  ( n11094 ) ? ( bv_8_45_n97 ) : ( n11790 ) ;
assign n11792 =  ( n11092 ) ? ( bv_8_60_n93 ) : ( n11791 ) ;
assign n11793 =  ( n11090 ) ? ( bv_8_21_n89 ) : ( n11792 ) ;
assign n11794 =  ( n11088 ) ? ( bv_8_201_n85 ) : ( n11793 ) ;
assign n11795 =  ( n11086 ) ? ( bv_8_135_n81 ) : ( n11794 ) ;
assign n11796 =  ( n11084 ) ? ( bv_8_170_n77 ) : ( n11795 ) ;
assign n11797 =  ( n11082 ) ? ( bv_8_80_n73 ) : ( n11796 ) ;
assign n11798 =  ( n11080 ) ? ( bv_8_165_n69 ) : ( n11797 ) ;
assign n11799 =  ( n11078 ) ? ( bv_8_3_n65 ) : ( n11798 ) ;
assign n11800 =  ( n11076 ) ? ( bv_8_89_n61 ) : ( n11799 ) ;
assign n11801 =  ( n11074 ) ? ( bv_8_9_n57 ) : ( n11800 ) ;
assign n11802 =  ( n11072 ) ? ( bv_8_26_n53 ) : ( n11801 ) ;
assign n11803 =  ( n11070 ) ? ( bv_8_101_n49 ) : ( n11802 ) ;
assign n11804 =  ( n11068 ) ? ( bv_8_215_n45 ) : ( n11803 ) ;
assign n11805 =  ( n11066 ) ? ( bv_8_132_n41 ) : ( n11804 ) ;
assign n11806 =  ( n11064 ) ? ( bv_8_208_n37 ) : ( n11805 ) ;
assign n11807 =  ( n11062 ) ? ( bv_8_130_n33 ) : ( n11806 ) ;
assign n11808 =  ( n11060 ) ? ( bv_8_41_n29 ) : ( n11807 ) ;
assign n11809 =  ( n11058 ) ? ( bv_8_90_n25 ) : ( n11808 ) ;
assign n11810 =  ( n11056 ) ? ( bv_8_30_n21 ) : ( n11809 ) ;
assign n11811 =  ( n11054 ) ? ( bv_8_123_n17 ) : ( n11810 ) ;
assign n11812 =  ( n11052 ) ? ( bv_8_168_n13 ) : ( n11811 ) ;
assign n11813 =  ( n11050 ) ? ( bv_8_109_n9 ) : ( n11812 ) ;
assign n11814 =  ( n11048 ) ? ( bv_8_44_n5 ) : ( n11813 ) ;
assign n11815 =  ( n11046 ) ^ ( n11814 )  ;
assign n11816 = key[87:80] ;
assign n11817 =  ( n11815 ) ^ ( n11816 )  ;
assign n11818 =  { ( n10275 ) , ( n11817 ) }  ;
assign n11819 = state_in[103:96] ;
assign n11820 =  ( n11819 ) == ( bv_8_255_n3 )  ;
assign n11821 = state_in[103:96] ;
assign n11822 =  ( n11821 ) == ( bv_8_254_n7 )  ;
assign n11823 = state_in[103:96] ;
assign n11824 =  ( n11823 ) == ( bv_8_253_n11 )  ;
assign n11825 = state_in[103:96] ;
assign n11826 =  ( n11825 ) == ( bv_8_252_n15 )  ;
assign n11827 = state_in[103:96] ;
assign n11828 =  ( n11827 ) == ( bv_8_251_n19 )  ;
assign n11829 = state_in[103:96] ;
assign n11830 =  ( n11829 ) == ( bv_8_250_n23 )  ;
assign n11831 = state_in[103:96] ;
assign n11832 =  ( n11831 ) == ( bv_8_249_n27 )  ;
assign n11833 = state_in[103:96] ;
assign n11834 =  ( n11833 ) == ( bv_8_248_n31 )  ;
assign n11835 = state_in[103:96] ;
assign n11836 =  ( n11835 ) == ( bv_8_247_n35 )  ;
assign n11837 = state_in[103:96] ;
assign n11838 =  ( n11837 ) == ( bv_8_246_n39 )  ;
assign n11839 = state_in[103:96] ;
assign n11840 =  ( n11839 ) == ( bv_8_245_n43 )  ;
assign n11841 = state_in[103:96] ;
assign n11842 =  ( n11841 ) == ( bv_8_244_n47 )  ;
assign n11843 = state_in[103:96] ;
assign n11844 =  ( n11843 ) == ( bv_8_243_n51 )  ;
assign n11845 = state_in[103:96] ;
assign n11846 =  ( n11845 ) == ( bv_8_242_n55 )  ;
assign n11847 = state_in[103:96] ;
assign n11848 =  ( n11847 ) == ( bv_8_241_n59 )  ;
assign n11849 = state_in[103:96] ;
assign n11850 =  ( n11849 ) == ( bv_8_240_n63 )  ;
assign n11851 = state_in[103:96] ;
assign n11852 =  ( n11851 ) == ( bv_8_239_n67 )  ;
assign n11853 = state_in[103:96] ;
assign n11854 =  ( n11853 ) == ( bv_8_238_n71 )  ;
assign n11855 = state_in[103:96] ;
assign n11856 =  ( n11855 ) == ( bv_8_237_n75 )  ;
assign n11857 = state_in[103:96] ;
assign n11858 =  ( n11857 ) == ( bv_8_236_n79 )  ;
assign n11859 = state_in[103:96] ;
assign n11860 =  ( n11859 ) == ( bv_8_235_n83 )  ;
assign n11861 = state_in[103:96] ;
assign n11862 =  ( n11861 ) == ( bv_8_234_n87 )  ;
assign n11863 = state_in[103:96] ;
assign n11864 =  ( n11863 ) == ( bv_8_233_n91 )  ;
assign n11865 = state_in[103:96] ;
assign n11866 =  ( n11865 ) == ( bv_8_232_n95 )  ;
assign n11867 = state_in[103:96] ;
assign n11868 =  ( n11867 ) == ( bv_8_231_n99 )  ;
assign n11869 = state_in[103:96] ;
assign n11870 =  ( n11869 ) == ( bv_8_230_n103 )  ;
assign n11871 = state_in[103:96] ;
assign n11872 =  ( n11871 ) == ( bv_8_229_n107 )  ;
assign n11873 = state_in[103:96] ;
assign n11874 =  ( n11873 ) == ( bv_8_228_n111 )  ;
assign n11875 = state_in[103:96] ;
assign n11876 =  ( n11875 ) == ( bv_8_227_n115 )  ;
assign n11877 = state_in[103:96] ;
assign n11878 =  ( n11877 ) == ( bv_8_226_n119 )  ;
assign n11879 = state_in[103:96] ;
assign n11880 =  ( n11879 ) == ( bv_8_225_n123 )  ;
assign n11881 = state_in[103:96] ;
assign n11882 =  ( n11881 ) == ( bv_8_224_n126 )  ;
assign n11883 = state_in[103:96] ;
assign n11884 =  ( n11883 ) == ( bv_8_223_n130 )  ;
assign n11885 = state_in[103:96] ;
assign n11886 =  ( n11885 ) == ( bv_8_222_n134 )  ;
assign n11887 = state_in[103:96] ;
assign n11888 =  ( n11887 ) == ( bv_8_221_n138 )  ;
assign n11889 = state_in[103:96] ;
assign n11890 =  ( n11889 ) == ( bv_8_220_n142 )  ;
assign n11891 = state_in[103:96] ;
assign n11892 =  ( n11891 ) == ( bv_8_219_n146 )  ;
assign n11893 = state_in[103:96] ;
assign n11894 =  ( n11893 ) == ( bv_8_218_n150 )  ;
assign n11895 = state_in[103:96] ;
assign n11896 =  ( n11895 ) == ( bv_8_217_n128 )  ;
assign n11897 = state_in[103:96] ;
assign n11898 =  ( n11897 ) == ( bv_8_216_n157 )  ;
assign n11899 = state_in[103:96] ;
assign n11900 =  ( n11899 ) == ( bv_8_215_n45 )  ;
assign n11901 = state_in[103:96] ;
assign n11902 =  ( n11901 ) == ( bv_8_214_n164 )  ;
assign n11903 = state_in[103:96] ;
assign n11904 =  ( n11903 ) == ( bv_8_213_n167 )  ;
assign n11905 = state_in[103:96] ;
assign n11906 =  ( n11905 ) == ( bv_8_212_n171 )  ;
assign n11907 = state_in[103:96] ;
assign n11908 =  ( n11907 ) == ( bv_8_211_n175 )  ;
assign n11909 = state_in[103:96] ;
assign n11910 =  ( n11909 ) == ( bv_8_210_n113 )  ;
assign n11911 = state_in[103:96] ;
assign n11912 =  ( n11911 ) == ( bv_8_209_n182 )  ;
assign n11913 = state_in[103:96] ;
assign n11914 =  ( n11913 ) == ( bv_8_208_n37 )  ;
assign n11915 = state_in[103:96] ;
assign n11916 =  ( n11915 ) == ( bv_8_207_n188 )  ;
assign n11917 = state_in[103:96] ;
assign n11918 =  ( n11917 ) == ( bv_8_206_n192 )  ;
assign n11919 = state_in[103:96] ;
assign n11920 =  ( n11919 ) == ( bv_8_205_n196 )  ;
assign n11921 = state_in[103:96] ;
assign n11922 =  ( n11921 ) == ( bv_8_204_n177 )  ;
assign n11923 = state_in[103:96] ;
assign n11924 =  ( n11923 ) == ( bv_8_203_n203 )  ;
assign n11925 = state_in[103:96] ;
assign n11926 =  ( n11925 ) == ( bv_8_202_n207 )  ;
assign n11927 = state_in[103:96] ;
assign n11928 =  ( n11927 ) == ( bv_8_201_n85 )  ;
assign n11929 = state_in[103:96] ;
assign n11930 =  ( n11929 ) == ( bv_8_200_n213 )  ;
assign n11931 = state_in[103:96] ;
assign n11932 =  ( n11931 ) == ( bv_8_199_n216 )  ;
assign n11933 = state_in[103:96] ;
assign n11934 =  ( n11933 ) == ( bv_8_198_n220 )  ;
assign n11935 = state_in[103:96] ;
assign n11936 =  ( n11935 ) == ( bv_8_197_n224 )  ;
assign n11937 = state_in[103:96] ;
assign n11938 =  ( n11937 ) == ( bv_8_196_n228 )  ;
assign n11939 = state_in[103:96] ;
assign n11940 =  ( n11939 ) == ( bv_8_195_n232 )  ;
assign n11941 = state_in[103:96] ;
assign n11942 =  ( n11941 ) == ( bv_8_194_n159 )  ;
assign n11943 = state_in[103:96] ;
assign n11944 =  ( n11943 ) == ( bv_8_193_n239 )  ;
assign n11945 = state_in[103:96] ;
assign n11946 =  ( n11945 ) == ( bv_8_192_n242 )  ;
assign n11947 = state_in[103:96] ;
assign n11948 =  ( n11947 ) == ( bv_8_191_n246 )  ;
assign n11949 = state_in[103:96] ;
assign n11950 =  ( n11949 ) == ( bv_8_190_n250 )  ;
assign n11951 = state_in[103:96] ;
assign n11952 =  ( n11951 ) == ( bv_8_189_n254 )  ;
assign n11953 = state_in[103:96] ;
assign n11954 =  ( n11953 ) == ( bv_8_188_n257 )  ;
assign n11955 = state_in[103:96] ;
assign n11956 =  ( n11955 ) == ( bv_8_187_n260 )  ;
assign n11957 = state_in[103:96] ;
assign n11958 =  ( n11957 ) == ( bv_8_186_n263 )  ;
assign n11959 = state_in[103:96] ;
assign n11960 =  ( n11959 ) == ( bv_8_185_n266 )  ;
assign n11961 = state_in[103:96] ;
assign n11962 =  ( n11961 ) == ( bv_8_184_n270 )  ;
assign n11963 = state_in[103:96] ;
assign n11964 =  ( n11963 ) == ( bv_8_183_n273 )  ;
assign n11965 = state_in[103:96] ;
assign n11966 =  ( n11965 ) == ( bv_8_182_n277 )  ;
assign n11967 = state_in[103:96] ;
assign n11968 =  ( n11967 ) == ( bv_8_181_n281 )  ;
assign n11969 = state_in[103:96] ;
assign n11970 =  ( n11969 ) == ( bv_8_180_n285 )  ;
assign n11971 = state_in[103:96] ;
assign n11972 =  ( n11971 ) == ( bv_8_179_n289 )  ;
assign n11973 = state_in[103:96] ;
assign n11974 =  ( n11973 ) == ( bv_8_178_n292 )  ;
assign n11975 = state_in[103:96] ;
assign n11976 =  ( n11975 ) == ( bv_8_177_n283 )  ;
assign n11977 = state_in[103:96] ;
assign n11978 =  ( n11977 ) == ( bv_8_176_n299 )  ;
assign n11979 = state_in[103:96] ;
assign n11980 =  ( n11979 ) == ( bv_8_175_n302 )  ;
assign n11981 = state_in[103:96] ;
assign n11982 =  ( n11981 ) == ( bv_8_174_n152 )  ;
assign n11983 = state_in[103:96] ;
assign n11984 =  ( n11983 ) == ( bv_8_173_n307 )  ;
assign n11985 = state_in[103:96] ;
assign n11986 =  ( n11985 ) == ( bv_8_172_n268 )  ;
assign n11987 = state_in[103:96] ;
assign n11988 =  ( n11987 ) == ( bv_8_171_n314 )  ;
assign n11989 = state_in[103:96] ;
assign n11990 =  ( n11989 ) == ( bv_8_170_n77 )  ;
assign n11991 = state_in[103:96] ;
assign n11992 =  ( n11991 ) == ( bv_8_169_n109 )  ;
assign n11993 = state_in[103:96] ;
assign n11994 =  ( n11993 ) == ( bv_8_168_n13 )  ;
assign n11995 = state_in[103:96] ;
assign n11996 =  ( n11995 ) == ( bv_8_167_n325 )  ;
assign n11997 = state_in[103:96] ;
assign n11998 =  ( n11997 ) == ( bv_8_166_n328 )  ;
assign n11999 = state_in[103:96] ;
assign n12000 =  ( n11999 ) == ( bv_8_165_n69 )  ;
assign n12001 = state_in[103:96] ;
assign n12002 =  ( n12001 ) == ( bv_8_164_n335 )  ;
assign n12003 = state_in[103:96] ;
assign n12004 =  ( n12003 ) == ( bv_8_163_n339 )  ;
assign n12005 = state_in[103:96] ;
assign n12006 =  ( n12005 ) == ( bv_8_162_n343 )  ;
assign n12007 = state_in[103:96] ;
assign n12008 =  ( n12007 ) == ( bv_8_161_n211 )  ;
assign n12009 = state_in[103:96] ;
assign n12010 =  ( n12009 ) == ( bv_8_160_n350 )  ;
assign n12011 = state_in[103:96] ;
assign n12012 =  ( n12011 ) == ( bv_8_159_n323 )  ;
assign n12013 = state_in[103:96] ;
assign n12014 =  ( n12013 ) == ( bv_8_158_n355 )  ;
assign n12015 = state_in[103:96] ;
assign n12016 =  ( n12015 ) == ( bv_8_157_n359 )  ;
assign n12017 = state_in[103:96] ;
assign n12018 =  ( n12017 ) == ( bv_8_156_n279 )  ;
assign n12019 = state_in[103:96] ;
assign n12020 =  ( n12019 ) == ( bv_8_155_n364 )  ;
assign n12021 = state_in[103:96] ;
assign n12022 =  ( n12021 ) == ( bv_8_154_n368 )  ;
assign n12023 = state_in[103:96] ;
assign n12024 =  ( n12023 ) == ( bv_8_153_n140 )  ;
assign n12025 = state_in[103:96] ;
assign n12026 =  ( n12025 ) == ( bv_8_152_n374 )  ;
assign n12027 = state_in[103:96] ;
assign n12028 =  ( n12027 ) == ( bv_8_151_n218 )  ;
assign n12029 = state_in[103:96] ;
assign n12030 =  ( n12029 ) == ( bv_8_150_n201 )  ;
assign n12031 = state_in[103:96] ;
assign n12032 =  ( n12031 ) == ( bv_8_149_n384 )  ;
assign n12033 = state_in[103:96] ;
assign n12034 =  ( n12033 ) == ( bv_8_148_n388 )  ;
assign n12035 = state_in[103:96] ;
assign n12036 =  ( n12035 ) == ( bv_8_147_n392 )  ;
assign n12037 = state_in[103:96] ;
assign n12038 =  ( n12037 ) == ( bv_8_146_n337 )  ;
assign n12039 = state_in[103:96] ;
assign n12040 =  ( n12039 ) == ( bv_8_145_n397 )  ;
assign n12041 = state_in[103:96] ;
assign n12042 =  ( n12041 ) == ( bv_8_144_n173 )  ;
assign n12043 = state_in[103:96] ;
assign n12044 =  ( n12043 ) == ( bv_8_143_n403 )  ;
assign n12045 = state_in[103:96] ;
assign n12046 =  ( n12045 ) == ( bv_8_142_n406 )  ;
assign n12047 = state_in[103:96] ;
assign n12048 =  ( n12047 ) == ( bv_8_141_n410 )  ;
assign n12049 = state_in[103:96] ;
assign n12050 =  ( n12049 ) == ( bv_8_140_n376 )  ;
assign n12051 = state_in[103:96] ;
assign n12052 =  ( n12051 ) == ( bv_8_139_n297 )  ;
assign n12053 = state_in[103:96] ;
assign n12054 =  ( n12053 ) == ( bv_8_138_n418 )  ;
assign n12055 = state_in[103:96] ;
assign n12056 =  ( n12055 ) == ( bv_8_137_n421 )  ;
assign n12057 = state_in[103:96] ;
assign n12058 =  ( n12057 ) == ( bv_8_136_n425 )  ;
assign n12059 = state_in[103:96] ;
assign n12060 =  ( n12059 ) == ( bv_8_135_n81 )  ;
assign n12061 = state_in[103:96] ;
assign n12062 =  ( n12061 ) == ( bv_8_134_n431 )  ;
assign n12063 = state_in[103:96] ;
assign n12064 =  ( n12063 ) == ( bv_8_133_n434 )  ;
assign n12065 = state_in[103:96] ;
assign n12066 =  ( n12065 ) == ( bv_8_132_n41 )  ;
assign n12067 = state_in[103:96] ;
assign n12068 =  ( n12067 ) == ( bv_8_131_n440 )  ;
assign n12069 = state_in[103:96] ;
assign n12070 =  ( n12069 ) == ( bv_8_130_n33 )  ;
assign n12071 = state_in[103:96] ;
assign n12072 =  ( n12071 ) == ( bv_8_129_n446 )  ;
assign n12073 = state_in[103:96] ;
assign n12074 =  ( n12073 ) == ( bv_8_128_n450 )  ;
assign n12075 = state_in[103:96] ;
assign n12076 =  ( n12075 ) == ( bv_8_127_n453 )  ;
assign n12077 = state_in[103:96] ;
assign n12078 =  ( n12077 ) == ( bv_8_126_n456 )  ;
assign n12079 = state_in[103:96] ;
assign n12080 =  ( n12079 ) == ( bv_8_125_n459 )  ;
assign n12081 = state_in[103:96] ;
assign n12082 =  ( n12081 ) == ( bv_8_124_n184 )  ;
assign n12083 = state_in[103:96] ;
assign n12084 =  ( n12083 ) == ( bv_8_123_n17 )  ;
assign n12085 = state_in[103:96] ;
assign n12086 =  ( n12085 ) == ( bv_8_122_n416 )  ;
assign n12087 = state_in[103:96] ;
assign n12088 =  ( n12087 ) == ( bv_8_121_n470 )  ;
assign n12089 = state_in[103:96] ;
assign n12090 =  ( n12089 ) == ( bv_8_120_n474 )  ;
assign n12091 = state_in[103:96] ;
assign n12092 =  ( n12091 ) == ( bv_8_119_n472 )  ;
assign n12093 = state_in[103:96] ;
assign n12094 =  ( n12093 ) == ( bv_8_118_n480 )  ;
assign n12095 = state_in[103:96] ;
assign n12096 =  ( n12095 ) == ( bv_8_117_n484 )  ;
assign n12097 = state_in[103:96] ;
assign n12098 =  ( n12097 ) == ( bv_8_116_n345 )  ;
assign n12099 = state_in[103:96] ;
assign n12100 =  ( n12099 ) == ( bv_8_115_n222 )  ;
assign n12101 = state_in[103:96] ;
assign n12102 =  ( n12101 ) == ( bv_8_114_n494 )  ;
assign n12103 = state_in[103:96] ;
assign n12104 =  ( n12103 ) == ( bv_8_113_n180 )  ;
assign n12105 = state_in[103:96] ;
assign n12106 =  ( n12105 ) == ( bv_8_112_n482 )  ;
assign n12107 = state_in[103:96] ;
assign n12108 =  ( n12107 ) == ( bv_8_111_n244 )  ;
assign n12109 = state_in[103:96] ;
assign n12110 =  ( n12109 ) == ( bv_8_110_n294 )  ;
assign n12111 = state_in[103:96] ;
assign n12112 =  ( n12111 ) == ( bv_8_109_n9 )  ;
assign n12113 = state_in[103:96] ;
assign n12114 =  ( n12113 ) == ( bv_8_108_n510 )  ;
assign n12115 = state_in[103:96] ;
assign n12116 =  ( n12115 ) == ( bv_8_107_n370 )  ;
assign n12117 = state_in[103:96] ;
assign n12118 =  ( n12117 ) == ( bv_8_106_n155 )  ;
assign n12119 = state_in[103:96] ;
assign n12120 =  ( n12119 ) == ( bv_8_105_n148 )  ;
assign n12121 = state_in[103:96] ;
assign n12122 =  ( n12121 ) == ( bv_8_104_n520 )  ;
assign n12123 = state_in[103:96] ;
assign n12124 =  ( n12123 ) == ( bv_8_103_n523 )  ;
assign n12125 = state_in[103:96] ;
assign n12126 =  ( n12125 ) == ( bv_8_102_n527 )  ;
assign n12127 = state_in[103:96] ;
assign n12128 =  ( n12127 ) == ( bv_8_101_n49 )  ;
assign n12129 = state_in[103:96] ;
assign n12130 =  ( n12129 ) == ( bv_8_100_n348 )  ;
assign n12131 = state_in[103:96] ;
assign n12132 =  ( n12131 ) == ( bv_8_99_n476 )  ;
assign n12133 = state_in[103:96] ;
assign n12134 =  ( n12133 ) == ( bv_8_98_n536 )  ;
assign n12135 = state_in[103:96] ;
assign n12136 =  ( n12135 ) == ( bv_8_97_n198 )  ;
assign n12137 = state_in[103:96] ;
assign n12138 =  ( n12137 ) == ( bv_8_96_n542 )  ;
assign n12139 = state_in[103:96] ;
assign n12140 =  ( n12139 ) == ( bv_8_95_n545 )  ;
assign n12141 = state_in[103:96] ;
assign n12142 =  ( n12141 ) == ( bv_8_94_n548 )  ;
assign n12143 = state_in[103:96] ;
assign n12144 =  ( n12143 ) == ( bv_8_93_n498 )  ;
assign n12145 = state_in[103:96] ;
assign n12146 =  ( n12145 ) == ( bv_8_92_n234 )  ;
assign n12147 = state_in[103:96] ;
assign n12148 =  ( n12147 ) == ( bv_8_91_n555 )  ;
assign n12149 = state_in[103:96] ;
assign n12150 =  ( n12149 ) == ( bv_8_90_n25 )  ;
assign n12151 = state_in[103:96] ;
assign n12152 =  ( n12151 ) == ( bv_8_89_n61 )  ;
assign n12153 = state_in[103:96] ;
assign n12154 =  ( n12153 ) == ( bv_8_88_n562 )  ;
assign n12155 = state_in[103:96] ;
assign n12156 =  ( n12155 ) == ( bv_8_87_n226 )  ;
assign n12157 = state_in[103:96] ;
assign n12158 =  ( n12157 ) == ( bv_8_86_n567 )  ;
assign n12159 = state_in[103:96] ;
assign n12160 =  ( n12159 ) == ( bv_8_85_n423 )  ;
assign n12161 = state_in[103:96] ;
assign n12162 =  ( n12161 ) == ( bv_8_84_n386 )  ;
assign n12163 = state_in[103:96] ;
assign n12164 =  ( n12163 ) == ( bv_8_83_n575 )  ;
assign n12165 = state_in[103:96] ;
assign n12166 =  ( n12165 ) == ( bv_8_82_n578 )  ;
assign n12167 = state_in[103:96] ;
assign n12168 =  ( n12167 ) == ( bv_8_81_n582 )  ;
assign n12169 = state_in[103:96] ;
assign n12170 =  ( n12169 ) == ( bv_8_80_n73 )  ;
assign n12171 = state_in[103:96] ;
assign n12172 =  ( n12171 ) == ( bv_8_79_n538 )  ;
assign n12173 = state_in[103:96] ;
assign n12174 =  ( n12173 ) == ( bv_8_78_n590 )  ;
assign n12175 = state_in[103:96] ;
assign n12176 =  ( n12175 ) == ( bv_8_77_n593 )  ;
assign n12177 = state_in[103:96] ;
assign n12178 =  ( n12177 ) == ( bv_8_76_n596 )  ;
assign n12179 = state_in[103:96] ;
assign n12180 =  ( n12179 ) == ( bv_8_75_n503 )  ;
assign n12181 = state_in[103:96] ;
assign n12182 =  ( n12181 ) == ( bv_8_74_n237 )  ;
assign n12183 = state_in[103:96] ;
assign n12184 =  ( n12183 ) == ( bv_8_73_n275 )  ;
assign n12185 = state_in[103:96] ;
assign n12186 =  ( n12185 ) == ( bv_8_72_n330 )  ;
assign n12187 = state_in[103:96] ;
assign n12188 =  ( n12187 ) == ( bv_8_71_n252 )  ;
assign n12189 = state_in[103:96] ;
assign n12190 =  ( n12189 ) == ( bv_8_70_n609 )  ;
assign n12191 = state_in[103:96] ;
assign n12192 =  ( n12191 ) == ( bv_8_69_n612 )  ;
assign n12193 = state_in[103:96] ;
assign n12194 =  ( n12193 ) == ( bv_8_68_n390 )  ;
assign n12195 = state_in[103:96] ;
assign n12196 =  ( n12195 ) == ( bv_8_67_n318 )  ;
assign n12197 = state_in[103:96] ;
assign n12198 =  ( n12197 ) == ( bv_8_66_n466 )  ;
assign n12199 = state_in[103:96] ;
assign n12200 =  ( n12199 ) == ( bv_8_65_n623 )  ;
assign n12201 = state_in[103:96] ;
assign n12202 =  ( n12201 ) == ( bv_8_64_n573 )  ;
assign n12203 = state_in[103:96] ;
assign n12204 =  ( n12203 ) == ( bv_8_63_n489 )  ;
assign n12205 = state_in[103:96] ;
assign n12206 =  ( n12205 ) == ( bv_8_62_n205 )  ;
assign n12207 = state_in[103:96] ;
assign n12208 =  ( n12207 ) == ( bv_8_61_n634 )  ;
assign n12209 = state_in[103:96] ;
assign n12210 =  ( n12209 ) == ( bv_8_60_n93 )  ;
assign n12211 = state_in[103:96] ;
assign n12212 =  ( n12211 ) == ( bv_8_59_n382 )  ;
assign n12213 = state_in[103:96] ;
assign n12214 =  ( n12213 ) == ( bv_8_58_n136 )  ;
assign n12215 = state_in[103:96] ;
assign n12216 =  ( n12215 ) == ( bv_8_57_n312 )  ;
assign n12217 = state_in[103:96] ;
assign n12218 =  ( n12217 ) == ( bv_8_56_n230 )  ;
assign n12219 = state_in[103:96] ;
assign n12220 =  ( n12219 ) == ( bv_8_55_n650 )  ;
assign n12221 = state_in[103:96] ;
assign n12222 =  ( n12221 ) == ( bv_8_54_n616 )  ;
assign n12223 = state_in[103:96] ;
assign n12224 =  ( n12223 ) == ( bv_8_53_n436 )  ;
assign n12225 = state_in[103:96] ;
assign n12226 =  ( n12225 ) == ( bv_8_52_n619 )  ;
assign n12227 = state_in[103:96] ;
assign n12228 =  ( n12227 ) == ( bv_8_51_n101 )  ;
assign n12229 = state_in[103:96] ;
assign n12230 =  ( n12229 ) == ( bv_8_50_n408 )  ;
assign n12231 = state_in[103:96] ;
assign n12232 =  ( n12231 ) == ( bv_8_49_n309 )  ;
assign n12233 = state_in[103:96] ;
assign n12234 =  ( n12233 ) == ( bv_8_48_n660 )  ;
assign n12235 = state_in[103:96] ;
assign n12236 =  ( n12235 ) == ( bv_8_47_n652 )  ;
assign n12237 = state_in[103:96] ;
assign n12238 =  ( n12237 ) == ( bv_8_46_n429 )  ;
assign n12239 = state_in[103:96] ;
assign n12240 =  ( n12239 ) == ( bv_8_45_n97 )  ;
assign n12241 = state_in[103:96] ;
assign n12242 =  ( n12241 ) == ( bv_8_44_n5 )  ;
assign n12243 = state_in[103:96] ;
assign n12244 =  ( n12243 ) == ( bv_8_43_n121 )  ;
assign n12245 = state_in[103:96] ;
assign n12246 =  ( n12245 ) == ( bv_8_42_n672 )  ;
assign n12247 = state_in[103:96] ;
assign n12248 =  ( n12247 ) == ( bv_8_41_n29 )  ;
assign n12249 = state_in[103:96] ;
assign n12250 =  ( n12249 ) == ( bv_8_40_n366 )  ;
assign n12251 = state_in[103:96] ;
assign n12252 =  ( n12251 ) == ( bv_8_39_n132 )  ;
assign n12253 = state_in[103:96] ;
assign n12254 =  ( n12253 ) == ( bv_8_38_n444 )  ;
assign n12255 = state_in[103:96] ;
assign n12256 =  ( n12255 ) == ( bv_8_37_n506 )  ;
assign n12257 = state_in[103:96] ;
assign n12258 =  ( n12257 ) == ( bv_8_36_n645 )  ;
assign n12259 = state_in[103:96] ;
assign n12260 =  ( n12259 ) == ( bv_8_35_n696 )  ;
assign n12261 = state_in[103:96] ;
assign n12262 =  ( n12261 ) == ( bv_8_34_n117 )  ;
assign n12263 = state_in[103:96] ;
assign n12264 =  ( n12263 ) == ( bv_8_33_n486 )  ;
assign n12265 = state_in[103:96] ;
assign n12266 =  ( n12265 ) == ( bv_8_32_n463 )  ;
assign n12267 = state_in[103:96] ;
assign n12268 =  ( n12267 ) == ( bv_8_31_n705 )  ;
assign n12269 = state_in[103:96] ;
assign n12270 =  ( n12269 ) == ( bv_8_30_n21 )  ;
assign n12271 = state_in[103:96] ;
assign n12272 =  ( n12271 ) == ( bv_8_29_n625 )  ;
assign n12273 = state_in[103:96] ;
assign n12274 =  ( n12273 ) == ( bv_8_28_n162 )  ;
assign n12275 = state_in[103:96] ;
assign n12276 =  ( n12275 ) == ( bv_8_27_n642 )  ;
assign n12277 = state_in[103:96] ;
assign n12278 =  ( n12277 ) == ( bv_8_26_n53 )  ;
assign n12279 = state_in[103:96] ;
assign n12280 =  ( n12279 ) == ( bv_8_25_n399 )  ;
assign n12281 = state_in[103:96] ;
assign n12282 =  ( n12281 ) == ( bv_8_24_n448 )  ;
assign n12283 = state_in[103:96] ;
assign n12284 =  ( n12283 ) == ( bv_8_23_n144 )  ;
assign n12285 = state_in[103:96] ;
assign n12286 =  ( n12285 ) == ( bv_8_22_n357 )  ;
assign n12287 = state_in[103:96] ;
assign n12288 =  ( n12287 ) == ( bv_8_21_n89 )  ;
assign n12289 = state_in[103:96] ;
assign n12290 =  ( n12289 ) == ( bv_8_20_n341 )  ;
assign n12291 = state_in[103:96] ;
assign n12292 =  ( n12291 ) == ( bv_8_19_n588 )  ;
assign n12293 = state_in[103:96] ;
assign n12294 =  ( n12293 ) == ( bv_8_18_n628 )  ;
assign n12295 = state_in[103:96] ;
assign n12296 =  ( n12295 ) == ( bv_8_17_n525 )  ;
assign n12297 = state_in[103:96] ;
assign n12298 =  ( n12297 ) == ( bv_8_16_n248 )  ;
assign n12299 = state_in[103:96] ;
assign n12300 =  ( n12299 ) == ( bv_8_15_n190 )  ;
assign n12301 = state_in[103:96] ;
assign n12302 =  ( n12301 ) == ( bv_8_14_n648 )  ;
assign n12303 = state_in[103:96] ;
assign n12304 =  ( n12303 ) == ( bv_8_13_n194 )  ;
assign n12305 = state_in[103:96] ;
assign n12306 =  ( n12305 ) == ( bv_8_12_n333 )  ;
assign n12307 = state_in[103:96] ;
assign n12308 =  ( n12307 ) == ( bv_8_11_n379 )  ;
assign n12309 = state_in[103:96] ;
assign n12310 =  ( n12309 ) == ( bv_8_10_n655 )  ;
assign n12311 = state_in[103:96] ;
assign n12312 =  ( n12311 ) == ( bv_8_9_n57 )  ;
assign n12313 = state_in[103:96] ;
assign n12314 =  ( n12313 ) == ( bv_8_8_n669 )  ;
assign n12315 = state_in[103:96] ;
assign n12316 =  ( n12315 ) == ( bv_8_7_n105 )  ;
assign n12317 = state_in[103:96] ;
assign n12318 =  ( n12317 ) == ( bv_8_6_n169 )  ;
assign n12319 = state_in[103:96] ;
assign n12320 =  ( n12319 ) == ( bv_8_5_n492 )  ;
assign n12321 = state_in[103:96] ;
assign n12322 =  ( n12321 ) == ( bv_8_4_n516 )  ;
assign n12323 = state_in[103:96] ;
assign n12324 =  ( n12323 ) == ( bv_8_3_n65 )  ;
assign n12325 = state_in[103:96] ;
assign n12326 =  ( n12325 ) == ( bv_8_2_n751 )  ;
assign n12327 = state_in[103:96] ;
assign n12328 =  ( n12327 ) == ( bv_8_1_n287 )  ;
assign n12329 = state_in[103:96] ;
assign n12330 =  ( n12329 ) == ( bv_8_0_n580 )  ;
assign n12331 =  ( n12330 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n12332 =  ( n12328 ) ? ( bv_8_248_n31 ) : ( n12331 ) ;
assign n12333 =  ( n12326 ) ? ( bv_8_238_n71 ) : ( n12332 ) ;
assign n12334 =  ( n12324 ) ? ( bv_8_246_n39 ) : ( n12333 ) ;
assign n12335 =  ( n12322 ) ? ( bv_8_255_n3 ) : ( n12334 ) ;
assign n12336 =  ( n12320 ) ? ( bv_8_214_n164 ) : ( n12335 ) ;
assign n12337 =  ( n12318 ) ? ( bv_8_222_n134 ) : ( n12336 ) ;
assign n12338 =  ( n12316 ) ? ( bv_8_145_n397 ) : ( n12337 ) ;
assign n12339 =  ( n12314 ) ? ( bv_8_96_n542 ) : ( n12338 ) ;
assign n12340 =  ( n12312 ) ? ( bv_8_2_n751 ) : ( n12339 ) ;
assign n12341 =  ( n12310 ) ? ( bv_8_206_n192 ) : ( n12340 ) ;
assign n12342 =  ( n12308 ) ? ( bv_8_86_n567 ) : ( n12341 ) ;
assign n12343 =  ( n12306 ) ? ( bv_8_231_n99 ) : ( n12342 ) ;
assign n12344 =  ( n12304 ) ? ( bv_8_181_n281 ) : ( n12343 ) ;
assign n12345 =  ( n12302 ) ? ( bv_8_77_n593 ) : ( n12344 ) ;
assign n12346 =  ( n12300 ) ? ( bv_8_236_n79 ) : ( n12345 ) ;
assign n12347 =  ( n12298 ) ? ( bv_8_143_n403 ) : ( n12346 ) ;
assign n12348 =  ( n12296 ) ? ( bv_8_31_n705 ) : ( n12347 ) ;
assign n12349 =  ( n12294 ) ? ( bv_8_137_n421 ) : ( n12348 ) ;
assign n12350 =  ( n12292 ) ? ( bv_8_250_n23 ) : ( n12349 ) ;
assign n12351 =  ( n12290 ) ? ( bv_8_239_n67 ) : ( n12350 ) ;
assign n12352 =  ( n12288 ) ? ( bv_8_178_n292 ) : ( n12351 ) ;
assign n12353 =  ( n12286 ) ? ( bv_8_142_n406 ) : ( n12352 ) ;
assign n12354 =  ( n12284 ) ? ( bv_8_251_n19 ) : ( n12353 ) ;
assign n12355 =  ( n12282 ) ? ( bv_8_65_n623 ) : ( n12354 ) ;
assign n12356 =  ( n12280 ) ? ( bv_8_179_n289 ) : ( n12355 ) ;
assign n12357 =  ( n12278 ) ? ( bv_8_95_n545 ) : ( n12356 ) ;
assign n12358 =  ( n12276 ) ? ( bv_8_69_n612 ) : ( n12357 ) ;
assign n12359 =  ( n12274 ) ? ( bv_8_35_n696 ) : ( n12358 ) ;
assign n12360 =  ( n12272 ) ? ( bv_8_83_n575 ) : ( n12359 ) ;
assign n12361 =  ( n12270 ) ? ( bv_8_228_n111 ) : ( n12360 ) ;
assign n12362 =  ( n12268 ) ? ( bv_8_155_n364 ) : ( n12361 ) ;
assign n12363 =  ( n12266 ) ? ( bv_8_117_n484 ) : ( n12362 ) ;
assign n12364 =  ( n12264 ) ? ( bv_8_225_n123 ) : ( n12363 ) ;
assign n12365 =  ( n12262 ) ? ( bv_8_61_n634 ) : ( n12364 ) ;
assign n12366 =  ( n12260 ) ? ( bv_8_76_n596 ) : ( n12365 ) ;
assign n12367 =  ( n12258 ) ? ( bv_8_108_n510 ) : ( n12366 ) ;
assign n12368 =  ( n12256 ) ? ( bv_8_126_n456 ) : ( n12367 ) ;
assign n12369 =  ( n12254 ) ? ( bv_8_245_n43 ) : ( n12368 ) ;
assign n12370 =  ( n12252 ) ? ( bv_8_131_n440 ) : ( n12369 ) ;
assign n12371 =  ( n12250 ) ? ( bv_8_104_n520 ) : ( n12370 ) ;
assign n12372 =  ( n12248 ) ? ( bv_8_81_n582 ) : ( n12371 ) ;
assign n12373 =  ( n12246 ) ? ( bv_8_209_n182 ) : ( n12372 ) ;
assign n12374 =  ( n12244 ) ? ( bv_8_249_n27 ) : ( n12373 ) ;
assign n12375 =  ( n12242 ) ? ( bv_8_226_n119 ) : ( n12374 ) ;
assign n12376 =  ( n12240 ) ? ( bv_8_171_n314 ) : ( n12375 ) ;
assign n12377 =  ( n12238 ) ? ( bv_8_98_n536 ) : ( n12376 ) ;
assign n12378 =  ( n12236 ) ? ( bv_8_42_n672 ) : ( n12377 ) ;
assign n12379 =  ( n12234 ) ? ( bv_8_8_n669 ) : ( n12378 ) ;
assign n12380 =  ( n12232 ) ? ( bv_8_149_n384 ) : ( n12379 ) ;
assign n12381 =  ( n12230 ) ? ( bv_8_70_n609 ) : ( n12380 ) ;
assign n12382 =  ( n12228 ) ? ( bv_8_157_n359 ) : ( n12381 ) ;
assign n12383 =  ( n12226 ) ? ( bv_8_48_n660 ) : ( n12382 ) ;
assign n12384 =  ( n12224 ) ? ( bv_8_55_n650 ) : ( n12383 ) ;
assign n12385 =  ( n12222 ) ? ( bv_8_10_n655 ) : ( n12384 ) ;
assign n12386 =  ( n12220 ) ? ( bv_8_47_n652 ) : ( n12385 ) ;
assign n12387 =  ( n12218 ) ? ( bv_8_14_n648 ) : ( n12386 ) ;
assign n12388 =  ( n12216 ) ? ( bv_8_36_n645 ) : ( n12387 ) ;
assign n12389 =  ( n12214 ) ? ( bv_8_27_n642 ) : ( n12388 ) ;
assign n12390 =  ( n12212 ) ? ( bv_8_223_n130 ) : ( n12389 ) ;
assign n12391 =  ( n12210 ) ? ( bv_8_205_n196 ) : ( n12390 ) ;
assign n12392 =  ( n12208 ) ? ( bv_8_78_n590 ) : ( n12391 ) ;
assign n12393 =  ( n12206 ) ? ( bv_8_127_n453 ) : ( n12392 ) ;
assign n12394 =  ( n12204 ) ? ( bv_8_234_n87 ) : ( n12393 ) ;
assign n12395 =  ( n12202 ) ? ( bv_8_18_n628 ) : ( n12394 ) ;
assign n12396 =  ( n12200 ) ? ( bv_8_29_n625 ) : ( n12395 ) ;
assign n12397 =  ( n12198 ) ? ( bv_8_88_n562 ) : ( n12396 ) ;
assign n12398 =  ( n12196 ) ? ( bv_8_52_n619 ) : ( n12397 ) ;
assign n12399 =  ( n12194 ) ? ( bv_8_54_n616 ) : ( n12398 ) ;
assign n12400 =  ( n12192 ) ? ( bv_8_220_n142 ) : ( n12399 ) ;
assign n12401 =  ( n12190 ) ? ( bv_8_180_n285 ) : ( n12400 ) ;
assign n12402 =  ( n12188 ) ? ( bv_8_91_n555 ) : ( n12401 ) ;
assign n12403 =  ( n12186 ) ? ( bv_8_164_n335 ) : ( n12402 ) ;
assign n12404 =  ( n12184 ) ? ( bv_8_118_n480 ) : ( n12403 ) ;
assign n12405 =  ( n12182 ) ? ( bv_8_183_n273 ) : ( n12404 ) ;
assign n12406 =  ( n12180 ) ? ( bv_8_125_n459 ) : ( n12405 ) ;
assign n12407 =  ( n12178 ) ? ( bv_8_82_n578 ) : ( n12406 ) ;
assign n12408 =  ( n12176 ) ? ( bv_8_221_n138 ) : ( n12407 ) ;
assign n12409 =  ( n12174 ) ? ( bv_8_94_n548 ) : ( n12408 ) ;
assign n12410 =  ( n12172 ) ? ( bv_8_19_n588 ) : ( n12409 ) ;
assign n12411 =  ( n12170 ) ? ( bv_8_166_n328 ) : ( n12410 ) ;
assign n12412 =  ( n12168 ) ? ( bv_8_185_n266 ) : ( n12411 ) ;
assign n12413 =  ( n12166 ) ? ( bv_8_0_n580 ) : ( n12412 ) ;
assign n12414 =  ( n12164 ) ? ( bv_8_193_n239 ) : ( n12413 ) ;
assign n12415 =  ( n12162 ) ? ( bv_8_64_n573 ) : ( n12414 ) ;
assign n12416 =  ( n12160 ) ? ( bv_8_227_n115 ) : ( n12415 ) ;
assign n12417 =  ( n12158 ) ? ( bv_8_121_n470 ) : ( n12416 ) ;
assign n12418 =  ( n12156 ) ? ( bv_8_182_n277 ) : ( n12417 ) ;
assign n12419 =  ( n12154 ) ? ( bv_8_212_n171 ) : ( n12418 ) ;
assign n12420 =  ( n12152 ) ? ( bv_8_141_n410 ) : ( n12419 ) ;
assign n12421 =  ( n12150 ) ? ( bv_8_103_n523 ) : ( n12420 ) ;
assign n12422 =  ( n12148 ) ? ( bv_8_114_n494 ) : ( n12421 ) ;
assign n12423 =  ( n12146 ) ? ( bv_8_148_n388 ) : ( n12422 ) ;
assign n12424 =  ( n12144 ) ? ( bv_8_152_n374 ) : ( n12423 ) ;
assign n12425 =  ( n12142 ) ? ( bv_8_176_n299 ) : ( n12424 ) ;
assign n12426 =  ( n12140 ) ? ( bv_8_133_n434 ) : ( n12425 ) ;
assign n12427 =  ( n12138 ) ? ( bv_8_187_n260 ) : ( n12426 ) ;
assign n12428 =  ( n12136 ) ? ( bv_8_197_n224 ) : ( n12427 ) ;
assign n12429 =  ( n12134 ) ? ( bv_8_79_n538 ) : ( n12428 ) ;
assign n12430 =  ( n12132 ) ? ( bv_8_237_n75 ) : ( n12429 ) ;
assign n12431 =  ( n12130 ) ? ( bv_8_134_n431 ) : ( n12430 ) ;
assign n12432 =  ( n12128 ) ? ( bv_8_154_n368 ) : ( n12431 ) ;
assign n12433 =  ( n12126 ) ? ( bv_8_102_n527 ) : ( n12432 ) ;
assign n12434 =  ( n12124 ) ? ( bv_8_17_n525 ) : ( n12433 ) ;
assign n12435 =  ( n12122 ) ? ( bv_8_138_n418 ) : ( n12434 ) ;
assign n12436 =  ( n12120 ) ? ( bv_8_233_n91 ) : ( n12435 ) ;
assign n12437 =  ( n12118 ) ? ( bv_8_4_n516 ) : ( n12436 ) ;
assign n12438 =  ( n12116 ) ? ( bv_8_254_n7 ) : ( n12437 ) ;
assign n12439 =  ( n12114 ) ? ( bv_8_160_n350 ) : ( n12438 ) ;
assign n12440 =  ( n12112 ) ? ( bv_8_120_n474 ) : ( n12439 ) ;
assign n12441 =  ( n12110 ) ? ( bv_8_37_n506 ) : ( n12440 ) ;
assign n12442 =  ( n12108 ) ? ( bv_8_75_n503 ) : ( n12441 ) ;
assign n12443 =  ( n12106 ) ? ( bv_8_162_n343 ) : ( n12442 ) ;
assign n12444 =  ( n12104 ) ? ( bv_8_93_n498 ) : ( n12443 ) ;
assign n12445 =  ( n12102 ) ? ( bv_8_128_n450 ) : ( n12444 ) ;
assign n12446 =  ( n12100 ) ? ( bv_8_5_n492 ) : ( n12445 ) ;
assign n12447 =  ( n12098 ) ? ( bv_8_63_n489 ) : ( n12446 ) ;
assign n12448 =  ( n12096 ) ? ( bv_8_33_n486 ) : ( n12447 ) ;
assign n12449 =  ( n12094 ) ? ( bv_8_112_n482 ) : ( n12448 ) ;
assign n12450 =  ( n12092 ) ? ( bv_8_241_n59 ) : ( n12449 ) ;
assign n12451 =  ( n12090 ) ? ( bv_8_99_n476 ) : ( n12450 ) ;
assign n12452 =  ( n12088 ) ? ( bv_8_119_n472 ) : ( n12451 ) ;
assign n12453 =  ( n12086 ) ? ( bv_8_175_n302 ) : ( n12452 ) ;
assign n12454 =  ( n12084 ) ? ( bv_8_66_n466 ) : ( n12453 ) ;
assign n12455 =  ( n12082 ) ? ( bv_8_32_n463 ) : ( n12454 ) ;
assign n12456 =  ( n12080 ) ? ( bv_8_229_n107 ) : ( n12455 ) ;
assign n12457 =  ( n12078 ) ? ( bv_8_253_n11 ) : ( n12456 ) ;
assign n12458 =  ( n12076 ) ? ( bv_8_191_n246 ) : ( n12457 ) ;
assign n12459 =  ( n12074 ) ? ( bv_8_129_n446 ) : ( n12458 ) ;
assign n12460 =  ( n12072 ) ? ( bv_8_24_n448 ) : ( n12459 ) ;
assign n12461 =  ( n12070 ) ? ( bv_8_38_n444 ) : ( n12460 ) ;
assign n12462 =  ( n12068 ) ? ( bv_8_195_n232 ) : ( n12461 ) ;
assign n12463 =  ( n12066 ) ? ( bv_8_190_n250 ) : ( n12462 ) ;
assign n12464 =  ( n12064 ) ? ( bv_8_53_n436 ) : ( n12463 ) ;
assign n12465 =  ( n12062 ) ? ( bv_8_136_n425 ) : ( n12464 ) ;
assign n12466 =  ( n12060 ) ? ( bv_8_46_n429 ) : ( n12465 ) ;
assign n12467 =  ( n12058 ) ? ( bv_8_147_n392 ) : ( n12466 ) ;
assign n12468 =  ( n12056 ) ? ( bv_8_85_n423 ) : ( n12467 ) ;
assign n12469 =  ( n12054 ) ? ( bv_8_252_n15 ) : ( n12468 ) ;
assign n12470 =  ( n12052 ) ? ( bv_8_122_n416 ) : ( n12469 ) ;
assign n12471 =  ( n12050 ) ? ( bv_8_200_n213 ) : ( n12470 ) ;
assign n12472 =  ( n12048 ) ? ( bv_8_186_n263 ) : ( n12471 ) ;
assign n12473 =  ( n12046 ) ? ( bv_8_50_n408 ) : ( n12472 ) ;
assign n12474 =  ( n12044 ) ? ( bv_8_230_n103 ) : ( n12473 ) ;
assign n12475 =  ( n12042 ) ? ( bv_8_192_n242 ) : ( n12474 ) ;
assign n12476 =  ( n12040 ) ? ( bv_8_25_n399 ) : ( n12475 ) ;
assign n12477 =  ( n12038 ) ? ( bv_8_158_n355 ) : ( n12476 ) ;
assign n12478 =  ( n12036 ) ? ( bv_8_163_n339 ) : ( n12477 ) ;
assign n12479 =  ( n12034 ) ? ( bv_8_68_n390 ) : ( n12478 ) ;
assign n12480 =  ( n12032 ) ? ( bv_8_84_n386 ) : ( n12479 ) ;
assign n12481 =  ( n12030 ) ? ( bv_8_59_n382 ) : ( n12480 ) ;
assign n12482 =  ( n12028 ) ? ( bv_8_11_n379 ) : ( n12481 ) ;
assign n12483 =  ( n12026 ) ? ( bv_8_140_n376 ) : ( n12482 ) ;
assign n12484 =  ( n12024 ) ? ( bv_8_199_n216 ) : ( n12483 ) ;
assign n12485 =  ( n12022 ) ? ( bv_8_107_n370 ) : ( n12484 ) ;
assign n12486 =  ( n12020 ) ? ( bv_8_40_n366 ) : ( n12485 ) ;
assign n12487 =  ( n12018 ) ? ( bv_8_167_n325 ) : ( n12486 ) ;
assign n12488 =  ( n12016 ) ? ( bv_8_188_n257 ) : ( n12487 ) ;
assign n12489 =  ( n12014 ) ? ( bv_8_22_n357 ) : ( n12488 ) ;
assign n12490 =  ( n12012 ) ? ( bv_8_173_n307 ) : ( n12489 ) ;
assign n12491 =  ( n12010 ) ? ( bv_8_219_n146 ) : ( n12490 ) ;
assign n12492 =  ( n12008 ) ? ( bv_8_100_n348 ) : ( n12491 ) ;
assign n12493 =  ( n12006 ) ? ( bv_8_116_n345 ) : ( n12492 ) ;
assign n12494 =  ( n12004 ) ? ( bv_8_20_n341 ) : ( n12493 ) ;
assign n12495 =  ( n12002 ) ? ( bv_8_146_n337 ) : ( n12494 ) ;
assign n12496 =  ( n12000 ) ? ( bv_8_12_n333 ) : ( n12495 ) ;
assign n12497 =  ( n11998 ) ? ( bv_8_72_n330 ) : ( n12496 ) ;
assign n12498 =  ( n11996 ) ? ( bv_8_184_n270 ) : ( n12497 ) ;
assign n12499 =  ( n11994 ) ? ( bv_8_159_n323 ) : ( n12498 ) ;
assign n12500 =  ( n11992 ) ? ( bv_8_189_n254 ) : ( n12499 ) ;
assign n12501 =  ( n11990 ) ? ( bv_8_67_n318 ) : ( n12500 ) ;
assign n12502 =  ( n11988 ) ? ( bv_8_196_n228 ) : ( n12501 ) ;
assign n12503 =  ( n11986 ) ? ( bv_8_57_n312 ) : ( n12502 ) ;
assign n12504 =  ( n11984 ) ? ( bv_8_49_n309 ) : ( n12503 ) ;
assign n12505 =  ( n11982 ) ? ( bv_8_211_n175 ) : ( n12504 ) ;
assign n12506 =  ( n11980 ) ? ( bv_8_242_n55 ) : ( n12505 ) ;
assign n12507 =  ( n11978 ) ? ( bv_8_213_n167 ) : ( n12506 ) ;
assign n12508 =  ( n11976 ) ? ( bv_8_139_n297 ) : ( n12507 ) ;
assign n12509 =  ( n11974 ) ? ( bv_8_110_n294 ) : ( n12508 ) ;
assign n12510 =  ( n11972 ) ? ( bv_8_218_n150 ) : ( n12509 ) ;
assign n12511 =  ( n11970 ) ? ( bv_8_1_n287 ) : ( n12510 ) ;
assign n12512 =  ( n11968 ) ? ( bv_8_177_n283 ) : ( n12511 ) ;
assign n12513 =  ( n11966 ) ? ( bv_8_156_n279 ) : ( n12512 ) ;
assign n12514 =  ( n11964 ) ? ( bv_8_73_n275 ) : ( n12513 ) ;
assign n12515 =  ( n11962 ) ? ( bv_8_216_n157 ) : ( n12514 ) ;
assign n12516 =  ( n11960 ) ? ( bv_8_172_n268 ) : ( n12515 ) ;
assign n12517 =  ( n11958 ) ? ( bv_8_243_n51 ) : ( n12516 ) ;
assign n12518 =  ( n11956 ) ? ( bv_8_207_n188 ) : ( n12517 ) ;
assign n12519 =  ( n11954 ) ? ( bv_8_202_n207 ) : ( n12518 ) ;
assign n12520 =  ( n11952 ) ? ( bv_8_244_n47 ) : ( n12519 ) ;
assign n12521 =  ( n11950 ) ? ( bv_8_71_n252 ) : ( n12520 ) ;
assign n12522 =  ( n11948 ) ? ( bv_8_16_n248 ) : ( n12521 ) ;
assign n12523 =  ( n11946 ) ? ( bv_8_111_n244 ) : ( n12522 ) ;
assign n12524 =  ( n11944 ) ? ( bv_8_240_n63 ) : ( n12523 ) ;
assign n12525 =  ( n11942 ) ? ( bv_8_74_n237 ) : ( n12524 ) ;
assign n12526 =  ( n11940 ) ? ( bv_8_92_n234 ) : ( n12525 ) ;
assign n12527 =  ( n11938 ) ? ( bv_8_56_n230 ) : ( n12526 ) ;
assign n12528 =  ( n11936 ) ? ( bv_8_87_n226 ) : ( n12527 ) ;
assign n12529 =  ( n11934 ) ? ( bv_8_115_n222 ) : ( n12528 ) ;
assign n12530 =  ( n11932 ) ? ( bv_8_151_n218 ) : ( n12529 ) ;
assign n12531 =  ( n11930 ) ? ( bv_8_203_n203 ) : ( n12530 ) ;
assign n12532 =  ( n11928 ) ? ( bv_8_161_n211 ) : ( n12531 ) ;
assign n12533 =  ( n11926 ) ? ( bv_8_232_n95 ) : ( n12532 ) ;
assign n12534 =  ( n11924 ) ? ( bv_8_62_n205 ) : ( n12533 ) ;
assign n12535 =  ( n11922 ) ? ( bv_8_150_n201 ) : ( n12534 ) ;
assign n12536 =  ( n11920 ) ? ( bv_8_97_n198 ) : ( n12535 ) ;
assign n12537 =  ( n11918 ) ? ( bv_8_13_n194 ) : ( n12536 ) ;
assign n12538 =  ( n11916 ) ? ( bv_8_15_n190 ) : ( n12537 ) ;
assign n12539 =  ( n11914 ) ? ( bv_8_224_n126 ) : ( n12538 ) ;
assign n12540 =  ( n11912 ) ? ( bv_8_124_n184 ) : ( n12539 ) ;
assign n12541 =  ( n11910 ) ? ( bv_8_113_n180 ) : ( n12540 ) ;
assign n12542 =  ( n11908 ) ? ( bv_8_204_n177 ) : ( n12541 ) ;
assign n12543 =  ( n11906 ) ? ( bv_8_144_n173 ) : ( n12542 ) ;
assign n12544 =  ( n11904 ) ? ( bv_8_6_n169 ) : ( n12543 ) ;
assign n12545 =  ( n11902 ) ? ( bv_8_247_n35 ) : ( n12544 ) ;
assign n12546 =  ( n11900 ) ? ( bv_8_28_n162 ) : ( n12545 ) ;
assign n12547 =  ( n11898 ) ? ( bv_8_194_n159 ) : ( n12546 ) ;
assign n12548 =  ( n11896 ) ? ( bv_8_106_n155 ) : ( n12547 ) ;
assign n12549 =  ( n11894 ) ? ( bv_8_174_n152 ) : ( n12548 ) ;
assign n12550 =  ( n11892 ) ? ( bv_8_105_n148 ) : ( n12549 ) ;
assign n12551 =  ( n11890 ) ? ( bv_8_23_n144 ) : ( n12550 ) ;
assign n12552 =  ( n11888 ) ? ( bv_8_153_n140 ) : ( n12551 ) ;
assign n12553 =  ( n11886 ) ? ( bv_8_58_n136 ) : ( n12552 ) ;
assign n12554 =  ( n11884 ) ? ( bv_8_39_n132 ) : ( n12553 ) ;
assign n12555 =  ( n11882 ) ? ( bv_8_217_n128 ) : ( n12554 ) ;
assign n12556 =  ( n11880 ) ? ( bv_8_235_n83 ) : ( n12555 ) ;
assign n12557 =  ( n11878 ) ? ( bv_8_43_n121 ) : ( n12556 ) ;
assign n12558 =  ( n11876 ) ? ( bv_8_34_n117 ) : ( n12557 ) ;
assign n12559 =  ( n11874 ) ? ( bv_8_210_n113 ) : ( n12558 ) ;
assign n12560 =  ( n11872 ) ? ( bv_8_169_n109 ) : ( n12559 ) ;
assign n12561 =  ( n11870 ) ? ( bv_8_7_n105 ) : ( n12560 ) ;
assign n12562 =  ( n11868 ) ? ( bv_8_51_n101 ) : ( n12561 ) ;
assign n12563 =  ( n11866 ) ? ( bv_8_45_n97 ) : ( n12562 ) ;
assign n12564 =  ( n11864 ) ? ( bv_8_60_n93 ) : ( n12563 ) ;
assign n12565 =  ( n11862 ) ? ( bv_8_21_n89 ) : ( n12564 ) ;
assign n12566 =  ( n11860 ) ? ( bv_8_201_n85 ) : ( n12565 ) ;
assign n12567 =  ( n11858 ) ? ( bv_8_135_n81 ) : ( n12566 ) ;
assign n12568 =  ( n11856 ) ? ( bv_8_170_n77 ) : ( n12567 ) ;
assign n12569 =  ( n11854 ) ? ( bv_8_80_n73 ) : ( n12568 ) ;
assign n12570 =  ( n11852 ) ? ( bv_8_165_n69 ) : ( n12569 ) ;
assign n12571 =  ( n11850 ) ? ( bv_8_3_n65 ) : ( n12570 ) ;
assign n12572 =  ( n11848 ) ? ( bv_8_89_n61 ) : ( n12571 ) ;
assign n12573 =  ( n11846 ) ? ( bv_8_9_n57 ) : ( n12572 ) ;
assign n12574 =  ( n11844 ) ? ( bv_8_26_n53 ) : ( n12573 ) ;
assign n12575 =  ( n11842 ) ? ( bv_8_101_n49 ) : ( n12574 ) ;
assign n12576 =  ( n11840 ) ? ( bv_8_215_n45 ) : ( n12575 ) ;
assign n12577 =  ( n11838 ) ? ( bv_8_132_n41 ) : ( n12576 ) ;
assign n12578 =  ( n11836 ) ? ( bv_8_208_n37 ) : ( n12577 ) ;
assign n12579 =  ( n11834 ) ? ( bv_8_130_n33 ) : ( n12578 ) ;
assign n12580 =  ( n11832 ) ? ( bv_8_41_n29 ) : ( n12579 ) ;
assign n12581 =  ( n11830 ) ? ( bv_8_90_n25 ) : ( n12580 ) ;
assign n12582 =  ( n11828 ) ? ( bv_8_30_n21 ) : ( n12581 ) ;
assign n12583 =  ( n11826 ) ? ( bv_8_123_n17 ) : ( n12582 ) ;
assign n12584 =  ( n11824 ) ? ( bv_8_168_n13 ) : ( n12583 ) ;
assign n12585 =  ( n11822 ) ? ( bv_8_109_n9 ) : ( n12584 ) ;
assign n12586 =  ( n11820 ) ? ( bv_8_44_n5 ) : ( n12585 ) ;
assign n12587 =  ( n7196 ) ^ ( n12586 )  ;
assign n12588 =  ( n12587 ) ^ ( n11043 )  ;
assign n12589 =  ( n12588 ) ^ ( n8733 )  ;
assign n12590 =  ( n12589 ) ^ ( n11814 )  ;
assign n12591 = key[79:72] ;
assign n12592 =  ( n12590 ) ^ ( n12591 )  ;
assign n12593 =  { ( n11818 ) , ( n12592 ) }  ;
assign n12594 =  ( n12586 ) ^ ( n11043 )  ;
assign n12595 =  ( n12594 ) ^ ( n7964 )  ;
assign n12596 =  ( n12595 ) ^ ( n8733 )  ;
assign n12597 =  ( n12596 ) ^ ( n10271 )  ;
assign n12598 = key[71:64] ;
assign n12599 =  ( n12597 ) ^ ( n12598 )  ;
assign n12600 =  { ( n12593 ) , ( n12599 ) }  ;
assign n12601 = state_in[111:104] ;
assign n12602 =  ( n12601 ) == ( bv_8_255_n3 )  ;
assign n12603 = state_in[111:104] ;
assign n12604 =  ( n12603 ) == ( bv_8_254_n7 )  ;
assign n12605 = state_in[111:104] ;
assign n12606 =  ( n12605 ) == ( bv_8_253_n11 )  ;
assign n12607 = state_in[111:104] ;
assign n12608 =  ( n12607 ) == ( bv_8_252_n15 )  ;
assign n12609 = state_in[111:104] ;
assign n12610 =  ( n12609 ) == ( bv_8_251_n19 )  ;
assign n12611 = state_in[111:104] ;
assign n12612 =  ( n12611 ) == ( bv_8_250_n23 )  ;
assign n12613 = state_in[111:104] ;
assign n12614 =  ( n12613 ) == ( bv_8_249_n27 )  ;
assign n12615 = state_in[111:104] ;
assign n12616 =  ( n12615 ) == ( bv_8_248_n31 )  ;
assign n12617 = state_in[111:104] ;
assign n12618 =  ( n12617 ) == ( bv_8_247_n35 )  ;
assign n12619 = state_in[111:104] ;
assign n12620 =  ( n12619 ) == ( bv_8_246_n39 )  ;
assign n12621 = state_in[111:104] ;
assign n12622 =  ( n12621 ) == ( bv_8_245_n43 )  ;
assign n12623 = state_in[111:104] ;
assign n12624 =  ( n12623 ) == ( bv_8_244_n47 )  ;
assign n12625 = state_in[111:104] ;
assign n12626 =  ( n12625 ) == ( bv_8_243_n51 )  ;
assign n12627 = state_in[111:104] ;
assign n12628 =  ( n12627 ) == ( bv_8_242_n55 )  ;
assign n12629 = state_in[111:104] ;
assign n12630 =  ( n12629 ) == ( bv_8_241_n59 )  ;
assign n12631 = state_in[111:104] ;
assign n12632 =  ( n12631 ) == ( bv_8_240_n63 )  ;
assign n12633 = state_in[111:104] ;
assign n12634 =  ( n12633 ) == ( bv_8_239_n67 )  ;
assign n12635 = state_in[111:104] ;
assign n12636 =  ( n12635 ) == ( bv_8_238_n71 )  ;
assign n12637 = state_in[111:104] ;
assign n12638 =  ( n12637 ) == ( bv_8_237_n75 )  ;
assign n12639 = state_in[111:104] ;
assign n12640 =  ( n12639 ) == ( bv_8_236_n79 )  ;
assign n12641 = state_in[111:104] ;
assign n12642 =  ( n12641 ) == ( bv_8_235_n83 )  ;
assign n12643 = state_in[111:104] ;
assign n12644 =  ( n12643 ) == ( bv_8_234_n87 )  ;
assign n12645 = state_in[111:104] ;
assign n12646 =  ( n12645 ) == ( bv_8_233_n91 )  ;
assign n12647 = state_in[111:104] ;
assign n12648 =  ( n12647 ) == ( bv_8_232_n95 )  ;
assign n12649 = state_in[111:104] ;
assign n12650 =  ( n12649 ) == ( bv_8_231_n99 )  ;
assign n12651 = state_in[111:104] ;
assign n12652 =  ( n12651 ) == ( bv_8_230_n103 )  ;
assign n12653 = state_in[111:104] ;
assign n12654 =  ( n12653 ) == ( bv_8_229_n107 )  ;
assign n12655 = state_in[111:104] ;
assign n12656 =  ( n12655 ) == ( bv_8_228_n111 )  ;
assign n12657 = state_in[111:104] ;
assign n12658 =  ( n12657 ) == ( bv_8_227_n115 )  ;
assign n12659 = state_in[111:104] ;
assign n12660 =  ( n12659 ) == ( bv_8_226_n119 )  ;
assign n12661 = state_in[111:104] ;
assign n12662 =  ( n12661 ) == ( bv_8_225_n123 )  ;
assign n12663 = state_in[111:104] ;
assign n12664 =  ( n12663 ) == ( bv_8_224_n126 )  ;
assign n12665 = state_in[111:104] ;
assign n12666 =  ( n12665 ) == ( bv_8_223_n130 )  ;
assign n12667 = state_in[111:104] ;
assign n12668 =  ( n12667 ) == ( bv_8_222_n134 )  ;
assign n12669 = state_in[111:104] ;
assign n12670 =  ( n12669 ) == ( bv_8_221_n138 )  ;
assign n12671 = state_in[111:104] ;
assign n12672 =  ( n12671 ) == ( bv_8_220_n142 )  ;
assign n12673 = state_in[111:104] ;
assign n12674 =  ( n12673 ) == ( bv_8_219_n146 )  ;
assign n12675 = state_in[111:104] ;
assign n12676 =  ( n12675 ) == ( bv_8_218_n150 )  ;
assign n12677 = state_in[111:104] ;
assign n12678 =  ( n12677 ) == ( bv_8_217_n128 )  ;
assign n12679 = state_in[111:104] ;
assign n12680 =  ( n12679 ) == ( bv_8_216_n157 )  ;
assign n12681 = state_in[111:104] ;
assign n12682 =  ( n12681 ) == ( bv_8_215_n45 )  ;
assign n12683 = state_in[111:104] ;
assign n12684 =  ( n12683 ) == ( bv_8_214_n164 )  ;
assign n12685 = state_in[111:104] ;
assign n12686 =  ( n12685 ) == ( bv_8_213_n167 )  ;
assign n12687 = state_in[111:104] ;
assign n12688 =  ( n12687 ) == ( bv_8_212_n171 )  ;
assign n12689 = state_in[111:104] ;
assign n12690 =  ( n12689 ) == ( bv_8_211_n175 )  ;
assign n12691 = state_in[111:104] ;
assign n12692 =  ( n12691 ) == ( bv_8_210_n113 )  ;
assign n12693 = state_in[111:104] ;
assign n12694 =  ( n12693 ) == ( bv_8_209_n182 )  ;
assign n12695 = state_in[111:104] ;
assign n12696 =  ( n12695 ) == ( bv_8_208_n37 )  ;
assign n12697 = state_in[111:104] ;
assign n12698 =  ( n12697 ) == ( bv_8_207_n188 )  ;
assign n12699 = state_in[111:104] ;
assign n12700 =  ( n12699 ) == ( bv_8_206_n192 )  ;
assign n12701 = state_in[111:104] ;
assign n12702 =  ( n12701 ) == ( bv_8_205_n196 )  ;
assign n12703 = state_in[111:104] ;
assign n12704 =  ( n12703 ) == ( bv_8_204_n177 )  ;
assign n12705 = state_in[111:104] ;
assign n12706 =  ( n12705 ) == ( bv_8_203_n203 )  ;
assign n12707 = state_in[111:104] ;
assign n12708 =  ( n12707 ) == ( bv_8_202_n207 )  ;
assign n12709 = state_in[111:104] ;
assign n12710 =  ( n12709 ) == ( bv_8_201_n85 )  ;
assign n12711 = state_in[111:104] ;
assign n12712 =  ( n12711 ) == ( bv_8_200_n213 )  ;
assign n12713 = state_in[111:104] ;
assign n12714 =  ( n12713 ) == ( bv_8_199_n216 )  ;
assign n12715 = state_in[111:104] ;
assign n12716 =  ( n12715 ) == ( bv_8_198_n220 )  ;
assign n12717 = state_in[111:104] ;
assign n12718 =  ( n12717 ) == ( bv_8_197_n224 )  ;
assign n12719 = state_in[111:104] ;
assign n12720 =  ( n12719 ) == ( bv_8_196_n228 )  ;
assign n12721 = state_in[111:104] ;
assign n12722 =  ( n12721 ) == ( bv_8_195_n232 )  ;
assign n12723 = state_in[111:104] ;
assign n12724 =  ( n12723 ) == ( bv_8_194_n159 )  ;
assign n12725 = state_in[111:104] ;
assign n12726 =  ( n12725 ) == ( bv_8_193_n239 )  ;
assign n12727 = state_in[111:104] ;
assign n12728 =  ( n12727 ) == ( bv_8_192_n242 )  ;
assign n12729 = state_in[111:104] ;
assign n12730 =  ( n12729 ) == ( bv_8_191_n246 )  ;
assign n12731 = state_in[111:104] ;
assign n12732 =  ( n12731 ) == ( bv_8_190_n250 )  ;
assign n12733 = state_in[111:104] ;
assign n12734 =  ( n12733 ) == ( bv_8_189_n254 )  ;
assign n12735 = state_in[111:104] ;
assign n12736 =  ( n12735 ) == ( bv_8_188_n257 )  ;
assign n12737 = state_in[111:104] ;
assign n12738 =  ( n12737 ) == ( bv_8_187_n260 )  ;
assign n12739 = state_in[111:104] ;
assign n12740 =  ( n12739 ) == ( bv_8_186_n263 )  ;
assign n12741 = state_in[111:104] ;
assign n12742 =  ( n12741 ) == ( bv_8_185_n266 )  ;
assign n12743 = state_in[111:104] ;
assign n12744 =  ( n12743 ) == ( bv_8_184_n270 )  ;
assign n12745 = state_in[111:104] ;
assign n12746 =  ( n12745 ) == ( bv_8_183_n273 )  ;
assign n12747 = state_in[111:104] ;
assign n12748 =  ( n12747 ) == ( bv_8_182_n277 )  ;
assign n12749 = state_in[111:104] ;
assign n12750 =  ( n12749 ) == ( bv_8_181_n281 )  ;
assign n12751 = state_in[111:104] ;
assign n12752 =  ( n12751 ) == ( bv_8_180_n285 )  ;
assign n12753 = state_in[111:104] ;
assign n12754 =  ( n12753 ) == ( bv_8_179_n289 )  ;
assign n12755 = state_in[111:104] ;
assign n12756 =  ( n12755 ) == ( bv_8_178_n292 )  ;
assign n12757 = state_in[111:104] ;
assign n12758 =  ( n12757 ) == ( bv_8_177_n283 )  ;
assign n12759 = state_in[111:104] ;
assign n12760 =  ( n12759 ) == ( bv_8_176_n299 )  ;
assign n12761 = state_in[111:104] ;
assign n12762 =  ( n12761 ) == ( bv_8_175_n302 )  ;
assign n12763 = state_in[111:104] ;
assign n12764 =  ( n12763 ) == ( bv_8_174_n152 )  ;
assign n12765 = state_in[111:104] ;
assign n12766 =  ( n12765 ) == ( bv_8_173_n307 )  ;
assign n12767 = state_in[111:104] ;
assign n12768 =  ( n12767 ) == ( bv_8_172_n268 )  ;
assign n12769 = state_in[111:104] ;
assign n12770 =  ( n12769 ) == ( bv_8_171_n314 )  ;
assign n12771 = state_in[111:104] ;
assign n12772 =  ( n12771 ) == ( bv_8_170_n77 )  ;
assign n12773 = state_in[111:104] ;
assign n12774 =  ( n12773 ) == ( bv_8_169_n109 )  ;
assign n12775 = state_in[111:104] ;
assign n12776 =  ( n12775 ) == ( bv_8_168_n13 )  ;
assign n12777 = state_in[111:104] ;
assign n12778 =  ( n12777 ) == ( bv_8_167_n325 )  ;
assign n12779 = state_in[111:104] ;
assign n12780 =  ( n12779 ) == ( bv_8_166_n328 )  ;
assign n12781 = state_in[111:104] ;
assign n12782 =  ( n12781 ) == ( bv_8_165_n69 )  ;
assign n12783 = state_in[111:104] ;
assign n12784 =  ( n12783 ) == ( bv_8_164_n335 )  ;
assign n12785 = state_in[111:104] ;
assign n12786 =  ( n12785 ) == ( bv_8_163_n339 )  ;
assign n12787 = state_in[111:104] ;
assign n12788 =  ( n12787 ) == ( bv_8_162_n343 )  ;
assign n12789 = state_in[111:104] ;
assign n12790 =  ( n12789 ) == ( bv_8_161_n211 )  ;
assign n12791 = state_in[111:104] ;
assign n12792 =  ( n12791 ) == ( bv_8_160_n350 )  ;
assign n12793 = state_in[111:104] ;
assign n12794 =  ( n12793 ) == ( bv_8_159_n323 )  ;
assign n12795 = state_in[111:104] ;
assign n12796 =  ( n12795 ) == ( bv_8_158_n355 )  ;
assign n12797 = state_in[111:104] ;
assign n12798 =  ( n12797 ) == ( bv_8_157_n359 )  ;
assign n12799 = state_in[111:104] ;
assign n12800 =  ( n12799 ) == ( bv_8_156_n279 )  ;
assign n12801 = state_in[111:104] ;
assign n12802 =  ( n12801 ) == ( bv_8_155_n364 )  ;
assign n12803 = state_in[111:104] ;
assign n12804 =  ( n12803 ) == ( bv_8_154_n368 )  ;
assign n12805 = state_in[111:104] ;
assign n12806 =  ( n12805 ) == ( bv_8_153_n140 )  ;
assign n12807 = state_in[111:104] ;
assign n12808 =  ( n12807 ) == ( bv_8_152_n374 )  ;
assign n12809 = state_in[111:104] ;
assign n12810 =  ( n12809 ) == ( bv_8_151_n218 )  ;
assign n12811 = state_in[111:104] ;
assign n12812 =  ( n12811 ) == ( bv_8_150_n201 )  ;
assign n12813 = state_in[111:104] ;
assign n12814 =  ( n12813 ) == ( bv_8_149_n384 )  ;
assign n12815 = state_in[111:104] ;
assign n12816 =  ( n12815 ) == ( bv_8_148_n388 )  ;
assign n12817 = state_in[111:104] ;
assign n12818 =  ( n12817 ) == ( bv_8_147_n392 )  ;
assign n12819 = state_in[111:104] ;
assign n12820 =  ( n12819 ) == ( bv_8_146_n337 )  ;
assign n12821 = state_in[111:104] ;
assign n12822 =  ( n12821 ) == ( bv_8_145_n397 )  ;
assign n12823 = state_in[111:104] ;
assign n12824 =  ( n12823 ) == ( bv_8_144_n173 )  ;
assign n12825 = state_in[111:104] ;
assign n12826 =  ( n12825 ) == ( bv_8_143_n403 )  ;
assign n12827 = state_in[111:104] ;
assign n12828 =  ( n12827 ) == ( bv_8_142_n406 )  ;
assign n12829 = state_in[111:104] ;
assign n12830 =  ( n12829 ) == ( bv_8_141_n410 )  ;
assign n12831 = state_in[111:104] ;
assign n12832 =  ( n12831 ) == ( bv_8_140_n376 )  ;
assign n12833 = state_in[111:104] ;
assign n12834 =  ( n12833 ) == ( bv_8_139_n297 )  ;
assign n12835 = state_in[111:104] ;
assign n12836 =  ( n12835 ) == ( bv_8_138_n418 )  ;
assign n12837 = state_in[111:104] ;
assign n12838 =  ( n12837 ) == ( bv_8_137_n421 )  ;
assign n12839 = state_in[111:104] ;
assign n12840 =  ( n12839 ) == ( bv_8_136_n425 )  ;
assign n12841 = state_in[111:104] ;
assign n12842 =  ( n12841 ) == ( bv_8_135_n81 )  ;
assign n12843 = state_in[111:104] ;
assign n12844 =  ( n12843 ) == ( bv_8_134_n431 )  ;
assign n12845 = state_in[111:104] ;
assign n12846 =  ( n12845 ) == ( bv_8_133_n434 )  ;
assign n12847 = state_in[111:104] ;
assign n12848 =  ( n12847 ) == ( bv_8_132_n41 )  ;
assign n12849 = state_in[111:104] ;
assign n12850 =  ( n12849 ) == ( bv_8_131_n440 )  ;
assign n12851 = state_in[111:104] ;
assign n12852 =  ( n12851 ) == ( bv_8_130_n33 )  ;
assign n12853 = state_in[111:104] ;
assign n12854 =  ( n12853 ) == ( bv_8_129_n446 )  ;
assign n12855 = state_in[111:104] ;
assign n12856 =  ( n12855 ) == ( bv_8_128_n450 )  ;
assign n12857 = state_in[111:104] ;
assign n12858 =  ( n12857 ) == ( bv_8_127_n453 )  ;
assign n12859 = state_in[111:104] ;
assign n12860 =  ( n12859 ) == ( bv_8_126_n456 )  ;
assign n12861 = state_in[111:104] ;
assign n12862 =  ( n12861 ) == ( bv_8_125_n459 )  ;
assign n12863 = state_in[111:104] ;
assign n12864 =  ( n12863 ) == ( bv_8_124_n184 )  ;
assign n12865 = state_in[111:104] ;
assign n12866 =  ( n12865 ) == ( bv_8_123_n17 )  ;
assign n12867 = state_in[111:104] ;
assign n12868 =  ( n12867 ) == ( bv_8_122_n416 )  ;
assign n12869 = state_in[111:104] ;
assign n12870 =  ( n12869 ) == ( bv_8_121_n470 )  ;
assign n12871 = state_in[111:104] ;
assign n12872 =  ( n12871 ) == ( bv_8_120_n474 )  ;
assign n12873 = state_in[111:104] ;
assign n12874 =  ( n12873 ) == ( bv_8_119_n472 )  ;
assign n12875 = state_in[111:104] ;
assign n12876 =  ( n12875 ) == ( bv_8_118_n480 )  ;
assign n12877 = state_in[111:104] ;
assign n12878 =  ( n12877 ) == ( bv_8_117_n484 )  ;
assign n12879 = state_in[111:104] ;
assign n12880 =  ( n12879 ) == ( bv_8_116_n345 )  ;
assign n12881 = state_in[111:104] ;
assign n12882 =  ( n12881 ) == ( bv_8_115_n222 )  ;
assign n12883 = state_in[111:104] ;
assign n12884 =  ( n12883 ) == ( bv_8_114_n494 )  ;
assign n12885 = state_in[111:104] ;
assign n12886 =  ( n12885 ) == ( bv_8_113_n180 )  ;
assign n12887 = state_in[111:104] ;
assign n12888 =  ( n12887 ) == ( bv_8_112_n482 )  ;
assign n12889 = state_in[111:104] ;
assign n12890 =  ( n12889 ) == ( bv_8_111_n244 )  ;
assign n12891 = state_in[111:104] ;
assign n12892 =  ( n12891 ) == ( bv_8_110_n294 )  ;
assign n12893 = state_in[111:104] ;
assign n12894 =  ( n12893 ) == ( bv_8_109_n9 )  ;
assign n12895 = state_in[111:104] ;
assign n12896 =  ( n12895 ) == ( bv_8_108_n510 )  ;
assign n12897 = state_in[111:104] ;
assign n12898 =  ( n12897 ) == ( bv_8_107_n370 )  ;
assign n12899 = state_in[111:104] ;
assign n12900 =  ( n12899 ) == ( bv_8_106_n155 )  ;
assign n12901 = state_in[111:104] ;
assign n12902 =  ( n12901 ) == ( bv_8_105_n148 )  ;
assign n12903 = state_in[111:104] ;
assign n12904 =  ( n12903 ) == ( bv_8_104_n520 )  ;
assign n12905 = state_in[111:104] ;
assign n12906 =  ( n12905 ) == ( bv_8_103_n523 )  ;
assign n12907 = state_in[111:104] ;
assign n12908 =  ( n12907 ) == ( bv_8_102_n527 )  ;
assign n12909 = state_in[111:104] ;
assign n12910 =  ( n12909 ) == ( bv_8_101_n49 )  ;
assign n12911 = state_in[111:104] ;
assign n12912 =  ( n12911 ) == ( bv_8_100_n348 )  ;
assign n12913 = state_in[111:104] ;
assign n12914 =  ( n12913 ) == ( bv_8_99_n476 )  ;
assign n12915 = state_in[111:104] ;
assign n12916 =  ( n12915 ) == ( bv_8_98_n536 )  ;
assign n12917 = state_in[111:104] ;
assign n12918 =  ( n12917 ) == ( bv_8_97_n198 )  ;
assign n12919 = state_in[111:104] ;
assign n12920 =  ( n12919 ) == ( bv_8_96_n542 )  ;
assign n12921 = state_in[111:104] ;
assign n12922 =  ( n12921 ) == ( bv_8_95_n545 )  ;
assign n12923 = state_in[111:104] ;
assign n12924 =  ( n12923 ) == ( bv_8_94_n548 )  ;
assign n12925 = state_in[111:104] ;
assign n12926 =  ( n12925 ) == ( bv_8_93_n498 )  ;
assign n12927 = state_in[111:104] ;
assign n12928 =  ( n12927 ) == ( bv_8_92_n234 )  ;
assign n12929 = state_in[111:104] ;
assign n12930 =  ( n12929 ) == ( bv_8_91_n555 )  ;
assign n12931 = state_in[111:104] ;
assign n12932 =  ( n12931 ) == ( bv_8_90_n25 )  ;
assign n12933 = state_in[111:104] ;
assign n12934 =  ( n12933 ) == ( bv_8_89_n61 )  ;
assign n12935 = state_in[111:104] ;
assign n12936 =  ( n12935 ) == ( bv_8_88_n562 )  ;
assign n12937 = state_in[111:104] ;
assign n12938 =  ( n12937 ) == ( bv_8_87_n226 )  ;
assign n12939 = state_in[111:104] ;
assign n12940 =  ( n12939 ) == ( bv_8_86_n567 )  ;
assign n12941 = state_in[111:104] ;
assign n12942 =  ( n12941 ) == ( bv_8_85_n423 )  ;
assign n12943 = state_in[111:104] ;
assign n12944 =  ( n12943 ) == ( bv_8_84_n386 )  ;
assign n12945 = state_in[111:104] ;
assign n12946 =  ( n12945 ) == ( bv_8_83_n575 )  ;
assign n12947 = state_in[111:104] ;
assign n12948 =  ( n12947 ) == ( bv_8_82_n578 )  ;
assign n12949 = state_in[111:104] ;
assign n12950 =  ( n12949 ) == ( bv_8_81_n582 )  ;
assign n12951 = state_in[111:104] ;
assign n12952 =  ( n12951 ) == ( bv_8_80_n73 )  ;
assign n12953 = state_in[111:104] ;
assign n12954 =  ( n12953 ) == ( bv_8_79_n538 )  ;
assign n12955 = state_in[111:104] ;
assign n12956 =  ( n12955 ) == ( bv_8_78_n590 )  ;
assign n12957 = state_in[111:104] ;
assign n12958 =  ( n12957 ) == ( bv_8_77_n593 )  ;
assign n12959 = state_in[111:104] ;
assign n12960 =  ( n12959 ) == ( bv_8_76_n596 )  ;
assign n12961 = state_in[111:104] ;
assign n12962 =  ( n12961 ) == ( bv_8_75_n503 )  ;
assign n12963 = state_in[111:104] ;
assign n12964 =  ( n12963 ) == ( bv_8_74_n237 )  ;
assign n12965 = state_in[111:104] ;
assign n12966 =  ( n12965 ) == ( bv_8_73_n275 )  ;
assign n12967 = state_in[111:104] ;
assign n12968 =  ( n12967 ) == ( bv_8_72_n330 )  ;
assign n12969 = state_in[111:104] ;
assign n12970 =  ( n12969 ) == ( bv_8_71_n252 )  ;
assign n12971 = state_in[111:104] ;
assign n12972 =  ( n12971 ) == ( bv_8_70_n609 )  ;
assign n12973 = state_in[111:104] ;
assign n12974 =  ( n12973 ) == ( bv_8_69_n612 )  ;
assign n12975 = state_in[111:104] ;
assign n12976 =  ( n12975 ) == ( bv_8_68_n390 )  ;
assign n12977 = state_in[111:104] ;
assign n12978 =  ( n12977 ) == ( bv_8_67_n318 )  ;
assign n12979 = state_in[111:104] ;
assign n12980 =  ( n12979 ) == ( bv_8_66_n466 )  ;
assign n12981 = state_in[111:104] ;
assign n12982 =  ( n12981 ) == ( bv_8_65_n623 )  ;
assign n12983 = state_in[111:104] ;
assign n12984 =  ( n12983 ) == ( bv_8_64_n573 )  ;
assign n12985 = state_in[111:104] ;
assign n12986 =  ( n12985 ) == ( bv_8_63_n489 )  ;
assign n12987 = state_in[111:104] ;
assign n12988 =  ( n12987 ) == ( bv_8_62_n205 )  ;
assign n12989 = state_in[111:104] ;
assign n12990 =  ( n12989 ) == ( bv_8_61_n634 )  ;
assign n12991 = state_in[111:104] ;
assign n12992 =  ( n12991 ) == ( bv_8_60_n93 )  ;
assign n12993 = state_in[111:104] ;
assign n12994 =  ( n12993 ) == ( bv_8_59_n382 )  ;
assign n12995 = state_in[111:104] ;
assign n12996 =  ( n12995 ) == ( bv_8_58_n136 )  ;
assign n12997 = state_in[111:104] ;
assign n12998 =  ( n12997 ) == ( bv_8_57_n312 )  ;
assign n12999 = state_in[111:104] ;
assign n13000 =  ( n12999 ) == ( bv_8_56_n230 )  ;
assign n13001 = state_in[111:104] ;
assign n13002 =  ( n13001 ) == ( bv_8_55_n650 )  ;
assign n13003 = state_in[111:104] ;
assign n13004 =  ( n13003 ) == ( bv_8_54_n616 )  ;
assign n13005 = state_in[111:104] ;
assign n13006 =  ( n13005 ) == ( bv_8_53_n436 )  ;
assign n13007 = state_in[111:104] ;
assign n13008 =  ( n13007 ) == ( bv_8_52_n619 )  ;
assign n13009 = state_in[111:104] ;
assign n13010 =  ( n13009 ) == ( bv_8_51_n101 )  ;
assign n13011 = state_in[111:104] ;
assign n13012 =  ( n13011 ) == ( bv_8_50_n408 )  ;
assign n13013 = state_in[111:104] ;
assign n13014 =  ( n13013 ) == ( bv_8_49_n309 )  ;
assign n13015 = state_in[111:104] ;
assign n13016 =  ( n13015 ) == ( bv_8_48_n660 )  ;
assign n13017 = state_in[111:104] ;
assign n13018 =  ( n13017 ) == ( bv_8_47_n652 )  ;
assign n13019 = state_in[111:104] ;
assign n13020 =  ( n13019 ) == ( bv_8_46_n429 )  ;
assign n13021 = state_in[111:104] ;
assign n13022 =  ( n13021 ) == ( bv_8_45_n97 )  ;
assign n13023 = state_in[111:104] ;
assign n13024 =  ( n13023 ) == ( bv_8_44_n5 )  ;
assign n13025 = state_in[111:104] ;
assign n13026 =  ( n13025 ) == ( bv_8_43_n121 )  ;
assign n13027 = state_in[111:104] ;
assign n13028 =  ( n13027 ) == ( bv_8_42_n672 )  ;
assign n13029 = state_in[111:104] ;
assign n13030 =  ( n13029 ) == ( bv_8_41_n29 )  ;
assign n13031 = state_in[111:104] ;
assign n13032 =  ( n13031 ) == ( bv_8_40_n366 )  ;
assign n13033 = state_in[111:104] ;
assign n13034 =  ( n13033 ) == ( bv_8_39_n132 )  ;
assign n13035 = state_in[111:104] ;
assign n13036 =  ( n13035 ) == ( bv_8_38_n444 )  ;
assign n13037 = state_in[111:104] ;
assign n13038 =  ( n13037 ) == ( bv_8_37_n506 )  ;
assign n13039 = state_in[111:104] ;
assign n13040 =  ( n13039 ) == ( bv_8_36_n645 )  ;
assign n13041 = state_in[111:104] ;
assign n13042 =  ( n13041 ) == ( bv_8_35_n696 )  ;
assign n13043 = state_in[111:104] ;
assign n13044 =  ( n13043 ) == ( bv_8_34_n117 )  ;
assign n13045 = state_in[111:104] ;
assign n13046 =  ( n13045 ) == ( bv_8_33_n486 )  ;
assign n13047 = state_in[111:104] ;
assign n13048 =  ( n13047 ) == ( bv_8_32_n463 )  ;
assign n13049 = state_in[111:104] ;
assign n13050 =  ( n13049 ) == ( bv_8_31_n705 )  ;
assign n13051 = state_in[111:104] ;
assign n13052 =  ( n13051 ) == ( bv_8_30_n21 )  ;
assign n13053 = state_in[111:104] ;
assign n13054 =  ( n13053 ) == ( bv_8_29_n625 )  ;
assign n13055 = state_in[111:104] ;
assign n13056 =  ( n13055 ) == ( bv_8_28_n162 )  ;
assign n13057 = state_in[111:104] ;
assign n13058 =  ( n13057 ) == ( bv_8_27_n642 )  ;
assign n13059 = state_in[111:104] ;
assign n13060 =  ( n13059 ) == ( bv_8_26_n53 )  ;
assign n13061 = state_in[111:104] ;
assign n13062 =  ( n13061 ) == ( bv_8_25_n399 )  ;
assign n13063 = state_in[111:104] ;
assign n13064 =  ( n13063 ) == ( bv_8_24_n448 )  ;
assign n13065 = state_in[111:104] ;
assign n13066 =  ( n13065 ) == ( bv_8_23_n144 )  ;
assign n13067 = state_in[111:104] ;
assign n13068 =  ( n13067 ) == ( bv_8_22_n357 )  ;
assign n13069 = state_in[111:104] ;
assign n13070 =  ( n13069 ) == ( bv_8_21_n89 )  ;
assign n13071 = state_in[111:104] ;
assign n13072 =  ( n13071 ) == ( bv_8_20_n341 )  ;
assign n13073 = state_in[111:104] ;
assign n13074 =  ( n13073 ) == ( bv_8_19_n588 )  ;
assign n13075 = state_in[111:104] ;
assign n13076 =  ( n13075 ) == ( bv_8_18_n628 )  ;
assign n13077 = state_in[111:104] ;
assign n13078 =  ( n13077 ) == ( bv_8_17_n525 )  ;
assign n13079 = state_in[111:104] ;
assign n13080 =  ( n13079 ) == ( bv_8_16_n248 )  ;
assign n13081 = state_in[111:104] ;
assign n13082 =  ( n13081 ) == ( bv_8_15_n190 )  ;
assign n13083 = state_in[111:104] ;
assign n13084 =  ( n13083 ) == ( bv_8_14_n648 )  ;
assign n13085 = state_in[111:104] ;
assign n13086 =  ( n13085 ) == ( bv_8_13_n194 )  ;
assign n13087 = state_in[111:104] ;
assign n13088 =  ( n13087 ) == ( bv_8_12_n333 )  ;
assign n13089 = state_in[111:104] ;
assign n13090 =  ( n13089 ) == ( bv_8_11_n379 )  ;
assign n13091 = state_in[111:104] ;
assign n13092 =  ( n13091 ) == ( bv_8_10_n655 )  ;
assign n13093 = state_in[111:104] ;
assign n13094 =  ( n13093 ) == ( bv_8_9_n57 )  ;
assign n13095 = state_in[111:104] ;
assign n13096 =  ( n13095 ) == ( bv_8_8_n669 )  ;
assign n13097 = state_in[111:104] ;
assign n13098 =  ( n13097 ) == ( bv_8_7_n105 )  ;
assign n13099 = state_in[111:104] ;
assign n13100 =  ( n13099 ) == ( bv_8_6_n169 )  ;
assign n13101 = state_in[111:104] ;
assign n13102 =  ( n13101 ) == ( bv_8_5_n492 )  ;
assign n13103 = state_in[111:104] ;
assign n13104 =  ( n13103 ) == ( bv_8_4_n516 )  ;
assign n13105 = state_in[111:104] ;
assign n13106 =  ( n13105 ) == ( bv_8_3_n65 )  ;
assign n13107 = state_in[111:104] ;
assign n13108 =  ( n13107 ) == ( bv_8_2_n751 )  ;
assign n13109 = state_in[111:104] ;
assign n13110 =  ( n13109 ) == ( bv_8_1_n287 )  ;
assign n13111 = state_in[111:104] ;
assign n13112 =  ( n13111 ) == ( bv_8_0_n580 )  ;
assign n13113 =  ( n13112 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n13114 =  ( n13110 ) ? ( bv_8_124_n184 ) : ( n13113 ) ;
assign n13115 =  ( n13108 ) ? ( bv_8_119_n472 ) : ( n13114 ) ;
assign n13116 =  ( n13106 ) ? ( bv_8_123_n17 ) : ( n13115 ) ;
assign n13117 =  ( n13104 ) ? ( bv_8_242_n55 ) : ( n13116 ) ;
assign n13118 =  ( n13102 ) ? ( bv_8_107_n370 ) : ( n13117 ) ;
assign n13119 =  ( n13100 ) ? ( bv_8_111_n244 ) : ( n13118 ) ;
assign n13120 =  ( n13098 ) ? ( bv_8_197_n224 ) : ( n13119 ) ;
assign n13121 =  ( n13096 ) ? ( bv_8_48_n660 ) : ( n13120 ) ;
assign n13122 =  ( n13094 ) ? ( bv_8_1_n287 ) : ( n13121 ) ;
assign n13123 =  ( n13092 ) ? ( bv_8_103_n523 ) : ( n13122 ) ;
assign n13124 =  ( n13090 ) ? ( bv_8_43_n121 ) : ( n13123 ) ;
assign n13125 =  ( n13088 ) ? ( bv_8_254_n7 ) : ( n13124 ) ;
assign n13126 =  ( n13086 ) ? ( bv_8_215_n45 ) : ( n13125 ) ;
assign n13127 =  ( n13084 ) ? ( bv_8_171_n314 ) : ( n13126 ) ;
assign n13128 =  ( n13082 ) ? ( bv_8_118_n480 ) : ( n13127 ) ;
assign n13129 =  ( n13080 ) ? ( bv_8_202_n207 ) : ( n13128 ) ;
assign n13130 =  ( n13078 ) ? ( bv_8_130_n33 ) : ( n13129 ) ;
assign n13131 =  ( n13076 ) ? ( bv_8_201_n85 ) : ( n13130 ) ;
assign n13132 =  ( n13074 ) ? ( bv_8_125_n459 ) : ( n13131 ) ;
assign n13133 =  ( n13072 ) ? ( bv_8_250_n23 ) : ( n13132 ) ;
assign n13134 =  ( n13070 ) ? ( bv_8_89_n61 ) : ( n13133 ) ;
assign n13135 =  ( n13068 ) ? ( bv_8_71_n252 ) : ( n13134 ) ;
assign n13136 =  ( n13066 ) ? ( bv_8_240_n63 ) : ( n13135 ) ;
assign n13137 =  ( n13064 ) ? ( bv_8_173_n307 ) : ( n13136 ) ;
assign n13138 =  ( n13062 ) ? ( bv_8_212_n171 ) : ( n13137 ) ;
assign n13139 =  ( n13060 ) ? ( bv_8_162_n343 ) : ( n13138 ) ;
assign n13140 =  ( n13058 ) ? ( bv_8_175_n302 ) : ( n13139 ) ;
assign n13141 =  ( n13056 ) ? ( bv_8_156_n279 ) : ( n13140 ) ;
assign n13142 =  ( n13054 ) ? ( bv_8_164_n335 ) : ( n13141 ) ;
assign n13143 =  ( n13052 ) ? ( bv_8_114_n494 ) : ( n13142 ) ;
assign n13144 =  ( n13050 ) ? ( bv_8_192_n242 ) : ( n13143 ) ;
assign n13145 =  ( n13048 ) ? ( bv_8_183_n273 ) : ( n13144 ) ;
assign n13146 =  ( n13046 ) ? ( bv_8_253_n11 ) : ( n13145 ) ;
assign n13147 =  ( n13044 ) ? ( bv_8_147_n392 ) : ( n13146 ) ;
assign n13148 =  ( n13042 ) ? ( bv_8_38_n444 ) : ( n13147 ) ;
assign n13149 =  ( n13040 ) ? ( bv_8_54_n616 ) : ( n13148 ) ;
assign n13150 =  ( n13038 ) ? ( bv_8_63_n489 ) : ( n13149 ) ;
assign n13151 =  ( n13036 ) ? ( bv_8_247_n35 ) : ( n13150 ) ;
assign n13152 =  ( n13034 ) ? ( bv_8_204_n177 ) : ( n13151 ) ;
assign n13153 =  ( n13032 ) ? ( bv_8_52_n619 ) : ( n13152 ) ;
assign n13154 =  ( n13030 ) ? ( bv_8_165_n69 ) : ( n13153 ) ;
assign n13155 =  ( n13028 ) ? ( bv_8_229_n107 ) : ( n13154 ) ;
assign n13156 =  ( n13026 ) ? ( bv_8_241_n59 ) : ( n13155 ) ;
assign n13157 =  ( n13024 ) ? ( bv_8_113_n180 ) : ( n13156 ) ;
assign n13158 =  ( n13022 ) ? ( bv_8_216_n157 ) : ( n13157 ) ;
assign n13159 =  ( n13020 ) ? ( bv_8_49_n309 ) : ( n13158 ) ;
assign n13160 =  ( n13018 ) ? ( bv_8_21_n89 ) : ( n13159 ) ;
assign n13161 =  ( n13016 ) ? ( bv_8_4_n516 ) : ( n13160 ) ;
assign n13162 =  ( n13014 ) ? ( bv_8_199_n216 ) : ( n13161 ) ;
assign n13163 =  ( n13012 ) ? ( bv_8_35_n696 ) : ( n13162 ) ;
assign n13164 =  ( n13010 ) ? ( bv_8_195_n232 ) : ( n13163 ) ;
assign n13165 =  ( n13008 ) ? ( bv_8_24_n448 ) : ( n13164 ) ;
assign n13166 =  ( n13006 ) ? ( bv_8_150_n201 ) : ( n13165 ) ;
assign n13167 =  ( n13004 ) ? ( bv_8_5_n492 ) : ( n13166 ) ;
assign n13168 =  ( n13002 ) ? ( bv_8_154_n368 ) : ( n13167 ) ;
assign n13169 =  ( n13000 ) ? ( bv_8_7_n105 ) : ( n13168 ) ;
assign n13170 =  ( n12998 ) ? ( bv_8_18_n628 ) : ( n13169 ) ;
assign n13171 =  ( n12996 ) ? ( bv_8_128_n450 ) : ( n13170 ) ;
assign n13172 =  ( n12994 ) ? ( bv_8_226_n119 ) : ( n13171 ) ;
assign n13173 =  ( n12992 ) ? ( bv_8_235_n83 ) : ( n13172 ) ;
assign n13174 =  ( n12990 ) ? ( bv_8_39_n132 ) : ( n13173 ) ;
assign n13175 =  ( n12988 ) ? ( bv_8_178_n292 ) : ( n13174 ) ;
assign n13176 =  ( n12986 ) ? ( bv_8_117_n484 ) : ( n13175 ) ;
assign n13177 =  ( n12984 ) ? ( bv_8_9_n57 ) : ( n13176 ) ;
assign n13178 =  ( n12982 ) ? ( bv_8_131_n440 ) : ( n13177 ) ;
assign n13179 =  ( n12980 ) ? ( bv_8_44_n5 ) : ( n13178 ) ;
assign n13180 =  ( n12978 ) ? ( bv_8_26_n53 ) : ( n13179 ) ;
assign n13181 =  ( n12976 ) ? ( bv_8_27_n642 ) : ( n13180 ) ;
assign n13182 =  ( n12974 ) ? ( bv_8_110_n294 ) : ( n13181 ) ;
assign n13183 =  ( n12972 ) ? ( bv_8_90_n25 ) : ( n13182 ) ;
assign n13184 =  ( n12970 ) ? ( bv_8_160_n350 ) : ( n13183 ) ;
assign n13185 =  ( n12968 ) ? ( bv_8_82_n578 ) : ( n13184 ) ;
assign n13186 =  ( n12966 ) ? ( bv_8_59_n382 ) : ( n13185 ) ;
assign n13187 =  ( n12964 ) ? ( bv_8_214_n164 ) : ( n13186 ) ;
assign n13188 =  ( n12962 ) ? ( bv_8_179_n289 ) : ( n13187 ) ;
assign n13189 =  ( n12960 ) ? ( bv_8_41_n29 ) : ( n13188 ) ;
assign n13190 =  ( n12958 ) ? ( bv_8_227_n115 ) : ( n13189 ) ;
assign n13191 =  ( n12956 ) ? ( bv_8_47_n652 ) : ( n13190 ) ;
assign n13192 =  ( n12954 ) ? ( bv_8_132_n41 ) : ( n13191 ) ;
assign n13193 =  ( n12952 ) ? ( bv_8_83_n575 ) : ( n13192 ) ;
assign n13194 =  ( n12950 ) ? ( bv_8_209_n182 ) : ( n13193 ) ;
assign n13195 =  ( n12948 ) ? ( bv_8_0_n580 ) : ( n13194 ) ;
assign n13196 =  ( n12946 ) ? ( bv_8_237_n75 ) : ( n13195 ) ;
assign n13197 =  ( n12944 ) ? ( bv_8_32_n463 ) : ( n13196 ) ;
assign n13198 =  ( n12942 ) ? ( bv_8_252_n15 ) : ( n13197 ) ;
assign n13199 =  ( n12940 ) ? ( bv_8_177_n283 ) : ( n13198 ) ;
assign n13200 =  ( n12938 ) ? ( bv_8_91_n555 ) : ( n13199 ) ;
assign n13201 =  ( n12936 ) ? ( bv_8_106_n155 ) : ( n13200 ) ;
assign n13202 =  ( n12934 ) ? ( bv_8_203_n203 ) : ( n13201 ) ;
assign n13203 =  ( n12932 ) ? ( bv_8_190_n250 ) : ( n13202 ) ;
assign n13204 =  ( n12930 ) ? ( bv_8_57_n312 ) : ( n13203 ) ;
assign n13205 =  ( n12928 ) ? ( bv_8_74_n237 ) : ( n13204 ) ;
assign n13206 =  ( n12926 ) ? ( bv_8_76_n596 ) : ( n13205 ) ;
assign n13207 =  ( n12924 ) ? ( bv_8_88_n562 ) : ( n13206 ) ;
assign n13208 =  ( n12922 ) ? ( bv_8_207_n188 ) : ( n13207 ) ;
assign n13209 =  ( n12920 ) ? ( bv_8_208_n37 ) : ( n13208 ) ;
assign n13210 =  ( n12918 ) ? ( bv_8_239_n67 ) : ( n13209 ) ;
assign n13211 =  ( n12916 ) ? ( bv_8_170_n77 ) : ( n13210 ) ;
assign n13212 =  ( n12914 ) ? ( bv_8_251_n19 ) : ( n13211 ) ;
assign n13213 =  ( n12912 ) ? ( bv_8_67_n318 ) : ( n13212 ) ;
assign n13214 =  ( n12910 ) ? ( bv_8_77_n593 ) : ( n13213 ) ;
assign n13215 =  ( n12908 ) ? ( bv_8_51_n101 ) : ( n13214 ) ;
assign n13216 =  ( n12906 ) ? ( bv_8_133_n434 ) : ( n13215 ) ;
assign n13217 =  ( n12904 ) ? ( bv_8_69_n612 ) : ( n13216 ) ;
assign n13218 =  ( n12902 ) ? ( bv_8_249_n27 ) : ( n13217 ) ;
assign n13219 =  ( n12900 ) ? ( bv_8_2_n751 ) : ( n13218 ) ;
assign n13220 =  ( n12898 ) ? ( bv_8_127_n453 ) : ( n13219 ) ;
assign n13221 =  ( n12896 ) ? ( bv_8_80_n73 ) : ( n13220 ) ;
assign n13222 =  ( n12894 ) ? ( bv_8_60_n93 ) : ( n13221 ) ;
assign n13223 =  ( n12892 ) ? ( bv_8_159_n323 ) : ( n13222 ) ;
assign n13224 =  ( n12890 ) ? ( bv_8_168_n13 ) : ( n13223 ) ;
assign n13225 =  ( n12888 ) ? ( bv_8_81_n582 ) : ( n13224 ) ;
assign n13226 =  ( n12886 ) ? ( bv_8_163_n339 ) : ( n13225 ) ;
assign n13227 =  ( n12884 ) ? ( bv_8_64_n573 ) : ( n13226 ) ;
assign n13228 =  ( n12882 ) ? ( bv_8_143_n403 ) : ( n13227 ) ;
assign n13229 =  ( n12880 ) ? ( bv_8_146_n337 ) : ( n13228 ) ;
assign n13230 =  ( n12878 ) ? ( bv_8_157_n359 ) : ( n13229 ) ;
assign n13231 =  ( n12876 ) ? ( bv_8_56_n230 ) : ( n13230 ) ;
assign n13232 =  ( n12874 ) ? ( bv_8_245_n43 ) : ( n13231 ) ;
assign n13233 =  ( n12872 ) ? ( bv_8_188_n257 ) : ( n13232 ) ;
assign n13234 =  ( n12870 ) ? ( bv_8_182_n277 ) : ( n13233 ) ;
assign n13235 =  ( n12868 ) ? ( bv_8_218_n150 ) : ( n13234 ) ;
assign n13236 =  ( n12866 ) ? ( bv_8_33_n486 ) : ( n13235 ) ;
assign n13237 =  ( n12864 ) ? ( bv_8_16_n248 ) : ( n13236 ) ;
assign n13238 =  ( n12862 ) ? ( bv_8_255_n3 ) : ( n13237 ) ;
assign n13239 =  ( n12860 ) ? ( bv_8_243_n51 ) : ( n13238 ) ;
assign n13240 =  ( n12858 ) ? ( bv_8_210_n113 ) : ( n13239 ) ;
assign n13241 =  ( n12856 ) ? ( bv_8_205_n196 ) : ( n13240 ) ;
assign n13242 =  ( n12854 ) ? ( bv_8_12_n333 ) : ( n13241 ) ;
assign n13243 =  ( n12852 ) ? ( bv_8_19_n588 ) : ( n13242 ) ;
assign n13244 =  ( n12850 ) ? ( bv_8_236_n79 ) : ( n13243 ) ;
assign n13245 =  ( n12848 ) ? ( bv_8_95_n545 ) : ( n13244 ) ;
assign n13246 =  ( n12846 ) ? ( bv_8_151_n218 ) : ( n13245 ) ;
assign n13247 =  ( n12844 ) ? ( bv_8_68_n390 ) : ( n13246 ) ;
assign n13248 =  ( n12842 ) ? ( bv_8_23_n144 ) : ( n13247 ) ;
assign n13249 =  ( n12840 ) ? ( bv_8_196_n228 ) : ( n13248 ) ;
assign n13250 =  ( n12838 ) ? ( bv_8_167_n325 ) : ( n13249 ) ;
assign n13251 =  ( n12836 ) ? ( bv_8_126_n456 ) : ( n13250 ) ;
assign n13252 =  ( n12834 ) ? ( bv_8_61_n634 ) : ( n13251 ) ;
assign n13253 =  ( n12832 ) ? ( bv_8_100_n348 ) : ( n13252 ) ;
assign n13254 =  ( n12830 ) ? ( bv_8_93_n498 ) : ( n13253 ) ;
assign n13255 =  ( n12828 ) ? ( bv_8_25_n399 ) : ( n13254 ) ;
assign n13256 =  ( n12826 ) ? ( bv_8_115_n222 ) : ( n13255 ) ;
assign n13257 =  ( n12824 ) ? ( bv_8_96_n542 ) : ( n13256 ) ;
assign n13258 =  ( n12822 ) ? ( bv_8_129_n446 ) : ( n13257 ) ;
assign n13259 =  ( n12820 ) ? ( bv_8_79_n538 ) : ( n13258 ) ;
assign n13260 =  ( n12818 ) ? ( bv_8_220_n142 ) : ( n13259 ) ;
assign n13261 =  ( n12816 ) ? ( bv_8_34_n117 ) : ( n13260 ) ;
assign n13262 =  ( n12814 ) ? ( bv_8_42_n672 ) : ( n13261 ) ;
assign n13263 =  ( n12812 ) ? ( bv_8_144_n173 ) : ( n13262 ) ;
assign n13264 =  ( n12810 ) ? ( bv_8_136_n425 ) : ( n13263 ) ;
assign n13265 =  ( n12808 ) ? ( bv_8_70_n609 ) : ( n13264 ) ;
assign n13266 =  ( n12806 ) ? ( bv_8_238_n71 ) : ( n13265 ) ;
assign n13267 =  ( n12804 ) ? ( bv_8_184_n270 ) : ( n13266 ) ;
assign n13268 =  ( n12802 ) ? ( bv_8_20_n341 ) : ( n13267 ) ;
assign n13269 =  ( n12800 ) ? ( bv_8_222_n134 ) : ( n13268 ) ;
assign n13270 =  ( n12798 ) ? ( bv_8_94_n548 ) : ( n13269 ) ;
assign n13271 =  ( n12796 ) ? ( bv_8_11_n379 ) : ( n13270 ) ;
assign n13272 =  ( n12794 ) ? ( bv_8_219_n146 ) : ( n13271 ) ;
assign n13273 =  ( n12792 ) ? ( bv_8_224_n126 ) : ( n13272 ) ;
assign n13274 =  ( n12790 ) ? ( bv_8_50_n408 ) : ( n13273 ) ;
assign n13275 =  ( n12788 ) ? ( bv_8_58_n136 ) : ( n13274 ) ;
assign n13276 =  ( n12786 ) ? ( bv_8_10_n655 ) : ( n13275 ) ;
assign n13277 =  ( n12784 ) ? ( bv_8_73_n275 ) : ( n13276 ) ;
assign n13278 =  ( n12782 ) ? ( bv_8_6_n169 ) : ( n13277 ) ;
assign n13279 =  ( n12780 ) ? ( bv_8_36_n645 ) : ( n13278 ) ;
assign n13280 =  ( n12778 ) ? ( bv_8_92_n234 ) : ( n13279 ) ;
assign n13281 =  ( n12776 ) ? ( bv_8_194_n159 ) : ( n13280 ) ;
assign n13282 =  ( n12774 ) ? ( bv_8_211_n175 ) : ( n13281 ) ;
assign n13283 =  ( n12772 ) ? ( bv_8_172_n268 ) : ( n13282 ) ;
assign n13284 =  ( n12770 ) ? ( bv_8_98_n536 ) : ( n13283 ) ;
assign n13285 =  ( n12768 ) ? ( bv_8_145_n397 ) : ( n13284 ) ;
assign n13286 =  ( n12766 ) ? ( bv_8_149_n384 ) : ( n13285 ) ;
assign n13287 =  ( n12764 ) ? ( bv_8_228_n111 ) : ( n13286 ) ;
assign n13288 =  ( n12762 ) ? ( bv_8_121_n470 ) : ( n13287 ) ;
assign n13289 =  ( n12760 ) ? ( bv_8_231_n99 ) : ( n13288 ) ;
assign n13290 =  ( n12758 ) ? ( bv_8_200_n213 ) : ( n13289 ) ;
assign n13291 =  ( n12756 ) ? ( bv_8_55_n650 ) : ( n13290 ) ;
assign n13292 =  ( n12754 ) ? ( bv_8_109_n9 ) : ( n13291 ) ;
assign n13293 =  ( n12752 ) ? ( bv_8_141_n410 ) : ( n13292 ) ;
assign n13294 =  ( n12750 ) ? ( bv_8_213_n167 ) : ( n13293 ) ;
assign n13295 =  ( n12748 ) ? ( bv_8_78_n590 ) : ( n13294 ) ;
assign n13296 =  ( n12746 ) ? ( bv_8_169_n109 ) : ( n13295 ) ;
assign n13297 =  ( n12744 ) ? ( bv_8_108_n510 ) : ( n13296 ) ;
assign n13298 =  ( n12742 ) ? ( bv_8_86_n567 ) : ( n13297 ) ;
assign n13299 =  ( n12740 ) ? ( bv_8_244_n47 ) : ( n13298 ) ;
assign n13300 =  ( n12738 ) ? ( bv_8_234_n87 ) : ( n13299 ) ;
assign n13301 =  ( n12736 ) ? ( bv_8_101_n49 ) : ( n13300 ) ;
assign n13302 =  ( n12734 ) ? ( bv_8_122_n416 ) : ( n13301 ) ;
assign n13303 =  ( n12732 ) ? ( bv_8_174_n152 ) : ( n13302 ) ;
assign n13304 =  ( n12730 ) ? ( bv_8_8_n669 ) : ( n13303 ) ;
assign n13305 =  ( n12728 ) ? ( bv_8_186_n263 ) : ( n13304 ) ;
assign n13306 =  ( n12726 ) ? ( bv_8_120_n474 ) : ( n13305 ) ;
assign n13307 =  ( n12724 ) ? ( bv_8_37_n506 ) : ( n13306 ) ;
assign n13308 =  ( n12722 ) ? ( bv_8_46_n429 ) : ( n13307 ) ;
assign n13309 =  ( n12720 ) ? ( bv_8_28_n162 ) : ( n13308 ) ;
assign n13310 =  ( n12718 ) ? ( bv_8_166_n328 ) : ( n13309 ) ;
assign n13311 =  ( n12716 ) ? ( bv_8_180_n285 ) : ( n13310 ) ;
assign n13312 =  ( n12714 ) ? ( bv_8_198_n220 ) : ( n13311 ) ;
assign n13313 =  ( n12712 ) ? ( bv_8_232_n95 ) : ( n13312 ) ;
assign n13314 =  ( n12710 ) ? ( bv_8_221_n138 ) : ( n13313 ) ;
assign n13315 =  ( n12708 ) ? ( bv_8_116_n345 ) : ( n13314 ) ;
assign n13316 =  ( n12706 ) ? ( bv_8_31_n705 ) : ( n13315 ) ;
assign n13317 =  ( n12704 ) ? ( bv_8_75_n503 ) : ( n13316 ) ;
assign n13318 =  ( n12702 ) ? ( bv_8_189_n254 ) : ( n13317 ) ;
assign n13319 =  ( n12700 ) ? ( bv_8_139_n297 ) : ( n13318 ) ;
assign n13320 =  ( n12698 ) ? ( bv_8_138_n418 ) : ( n13319 ) ;
assign n13321 =  ( n12696 ) ? ( bv_8_112_n482 ) : ( n13320 ) ;
assign n13322 =  ( n12694 ) ? ( bv_8_62_n205 ) : ( n13321 ) ;
assign n13323 =  ( n12692 ) ? ( bv_8_181_n281 ) : ( n13322 ) ;
assign n13324 =  ( n12690 ) ? ( bv_8_102_n527 ) : ( n13323 ) ;
assign n13325 =  ( n12688 ) ? ( bv_8_72_n330 ) : ( n13324 ) ;
assign n13326 =  ( n12686 ) ? ( bv_8_3_n65 ) : ( n13325 ) ;
assign n13327 =  ( n12684 ) ? ( bv_8_246_n39 ) : ( n13326 ) ;
assign n13328 =  ( n12682 ) ? ( bv_8_14_n648 ) : ( n13327 ) ;
assign n13329 =  ( n12680 ) ? ( bv_8_97_n198 ) : ( n13328 ) ;
assign n13330 =  ( n12678 ) ? ( bv_8_53_n436 ) : ( n13329 ) ;
assign n13331 =  ( n12676 ) ? ( bv_8_87_n226 ) : ( n13330 ) ;
assign n13332 =  ( n12674 ) ? ( bv_8_185_n266 ) : ( n13331 ) ;
assign n13333 =  ( n12672 ) ? ( bv_8_134_n431 ) : ( n13332 ) ;
assign n13334 =  ( n12670 ) ? ( bv_8_193_n239 ) : ( n13333 ) ;
assign n13335 =  ( n12668 ) ? ( bv_8_29_n625 ) : ( n13334 ) ;
assign n13336 =  ( n12666 ) ? ( bv_8_158_n355 ) : ( n13335 ) ;
assign n13337 =  ( n12664 ) ? ( bv_8_225_n123 ) : ( n13336 ) ;
assign n13338 =  ( n12662 ) ? ( bv_8_248_n31 ) : ( n13337 ) ;
assign n13339 =  ( n12660 ) ? ( bv_8_152_n374 ) : ( n13338 ) ;
assign n13340 =  ( n12658 ) ? ( bv_8_17_n525 ) : ( n13339 ) ;
assign n13341 =  ( n12656 ) ? ( bv_8_105_n148 ) : ( n13340 ) ;
assign n13342 =  ( n12654 ) ? ( bv_8_217_n128 ) : ( n13341 ) ;
assign n13343 =  ( n12652 ) ? ( bv_8_142_n406 ) : ( n13342 ) ;
assign n13344 =  ( n12650 ) ? ( bv_8_148_n388 ) : ( n13343 ) ;
assign n13345 =  ( n12648 ) ? ( bv_8_155_n364 ) : ( n13344 ) ;
assign n13346 =  ( n12646 ) ? ( bv_8_30_n21 ) : ( n13345 ) ;
assign n13347 =  ( n12644 ) ? ( bv_8_135_n81 ) : ( n13346 ) ;
assign n13348 =  ( n12642 ) ? ( bv_8_233_n91 ) : ( n13347 ) ;
assign n13349 =  ( n12640 ) ? ( bv_8_206_n192 ) : ( n13348 ) ;
assign n13350 =  ( n12638 ) ? ( bv_8_85_n423 ) : ( n13349 ) ;
assign n13351 =  ( n12636 ) ? ( bv_8_40_n366 ) : ( n13350 ) ;
assign n13352 =  ( n12634 ) ? ( bv_8_223_n130 ) : ( n13351 ) ;
assign n13353 =  ( n12632 ) ? ( bv_8_140_n376 ) : ( n13352 ) ;
assign n13354 =  ( n12630 ) ? ( bv_8_161_n211 ) : ( n13353 ) ;
assign n13355 =  ( n12628 ) ? ( bv_8_137_n421 ) : ( n13354 ) ;
assign n13356 =  ( n12626 ) ? ( bv_8_13_n194 ) : ( n13355 ) ;
assign n13357 =  ( n12624 ) ? ( bv_8_191_n246 ) : ( n13356 ) ;
assign n13358 =  ( n12622 ) ? ( bv_8_230_n103 ) : ( n13357 ) ;
assign n13359 =  ( n12620 ) ? ( bv_8_66_n466 ) : ( n13358 ) ;
assign n13360 =  ( n12618 ) ? ( bv_8_104_n520 ) : ( n13359 ) ;
assign n13361 =  ( n12616 ) ? ( bv_8_65_n623 ) : ( n13360 ) ;
assign n13362 =  ( n12614 ) ? ( bv_8_153_n140 ) : ( n13361 ) ;
assign n13363 =  ( n12612 ) ? ( bv_8_45_n97 ) : ( n13362 ) ;
assign n13364 =  ( n12610 ) ? ( bv_8_15_n190 ) : ( n13363 ) ;
assign n13365 =  ( n12608 ) ? ( bv_8_176_n299 ) : ( n13364 ) ;
assign n13366 =  ( n12606 ) ? ( bv_8_84_n386 ) : ( n13365 ) ;
assign n13367 =  ( n12604 ) ? ( bv_8_187_n260 ) : ( n13366 ) ;
assign n13368 =  ( n12602 ) ? ( bv_8_22_n357 ) : ( n13367 ) ;
assign n13369 = state_in[71:64] ;
assign n13370 =  ( n13369 ) == ( bv_8_255_n3 )  ;
assign n13371 = state_in[71:64] ;
assign n13372 =  ( n13371 ) == ( bv_8_254_n7 )  ;
assign n13373 = state_in[71:64] ;
assign n13374 =  ( n13373 ) == ( bv_8_253_n11 )  ;
assign n13375 = state_in[71:64] ;
assign n13376 =  ( n13375 ) == ( bv_8_252_n15 )  ;
assign n13377 = state_in[71:64] ;
assign n13378 =  ( n13377 ) == ( bv_8_251_n19 )  ;
assign n13379 = state_in[71:64] ;
assign n13380 =  ( n13379 ) == ( bv_8_250_n23 )  ;
assign n13381 = state_in[71:64] ;
assign n13382 =  ( n13381 ) == ( bv_8_249_n27 )  ;
assign n13383 = state_in[71:64] ;
assign n13384 =  ( n13383 ) == ( bv_8_248_n31 )  ;
assign n13385 = state_in[71:64] ;
assign n13386 =  ( n13385 ) == ( bv_8_247_n35 )  ;
assign n13387 = state_in[71:64] ;
assign n13388 =  ( n13387 ) == ( bv_8_246_n39 )  ;
assign n13389 = state_in[71:64] ;
assign n13390 =  ( n13389 ) == ( bv_8_245_n43 )  ;
assign n13391 = state_in[71:64] ;
assign n13392 =  ( n13391 ) == ( bv_8_244_n47 )  ;
assign n13393 = state_in[71:64] ;
assign n13394 =  ( n13393 ) == ( bv_8_243_n51 )  ;
assign n13395 = state_in[71:64] ;
assign n13396 =  ( n13395 ) == ( bv_8_242_n55 )  ;
assign n13397 = state_in[71:64] ;
assign n13398 =  ( n13397 ) == ( bv_8_241_n59 )  ;
assign n13399 = state_in[71:64] ;
assign n13400 =  ( n13399 ) == ( bv_8_240_n63 )  ;
assign n13401 = state_in[71:64] ;
assign n13402 =  ( n13401 ) == ( bv_8_239_n67 )  ;
assign n13403 = state_in[71:64] ;
assign n13404 =  ( n13403 ) == ( bv_8_238_n71 )  ;
assign n13405 = state_in[71:64] ;
assign n13406 =  ( n13405 ) == ( bv_8_237_n75 )  ;
assign n13407 = state_in[71:64] ;
assign n13408 =  ( n13407 ) == ( bv_8_236_n79 )  ;
assign n13409 = state_in[71:64] ;
assign n13410 =  ( n13409 ) == ( bv_8_235_n83 )  ;
assign n13411 = state_in[71:64] ;
assign n13412 =  ( n13411 ) == ( bv_8_234_n87 )  ;
assign n13413 = state_in[71:64] ;
assign n13414 =  ( n13413 ) == ( bv_8_233_n91 )  ;
assign n13415 = state_in[71:64] ;
assign n13416 =  ( n13415 ) == ( bv_8_232_n95 )  ;
assign n13417 = state_in[71:64] ;
assign n13418 =  ( n13417 ) == ( bv_8_231_n99 )  ;
assign n13419 = state_in[71:64] ;
assign n13420 =  ( n13419 ) == ( bv_8_230_n103 )  ;
assign n13421 = state_in[71:64] ;
assign n13422 =  ( n13421 ) == ( bv_8_229_n107 )  ;
assign n13423 = state_in[71:64] ;
assign n13424 =  ( n13423 ) == ( bv_8_228_n111 )  ;
assign n13425 = state_in[71:64] ;
assign n13426 =  ( n13425 ) == ( bv_8_227_n115 )  ;
assign n13427 = state_in[71:64] ;
assign n13428 =  ( n13427 ) == ( bv_8_226_n119 )  ;
assign n13429 = state_in[71:64] ;
assign n13430 =  ( n13429 ) == ( bv_8_225_n123 )  ;
assign n13431 = state_in[71:64] ;
assign n13432 =  ( n13431 ) == ( bv_8_224_n126 )  ;
assign n13433 = state_in[71:64] ;
assign n13434 =  ( n13433 ) == ( bv_8_223_n130 )  ;
assign n13435 = state_in[71:64] ;
assign n13436 =  ( n13435 ) == ( bv_8_222_n134 )  ;
assign n13437 = state_in[71:64] ;
assign n13438 =  ( n13437 ) == ( bv_8_221_n138 )  ;
assign n13439 = state_in[71:64] ;
assign n13440 =  ( n13439 ) == ( bv_8_220_n142 )  ;
assign n13441 = state_in[71:64] ;
assign n13442 =  ( n13441 ) == ( bv_8_219_n146 )  ;
assign n13443 = state_in[71:64] ;
assign n13444 =  ( n13443 ) == ( bv_8_218_n150 )  ;
assign n13445 = state_in[71:64] ;
assign n13446 =  ( n13445 ) == ( bv_8_217_n128 )  ;
assign n13447 = state_in[71:64] ;
assign n13448 =  ( n13447 ) == ( bv_8_216_n157 )  ;
assign n13449 = state_in[71:64] ;
assign n13450 =  ( n13449 ) == ( bv_8_215_n45 )  ;
assign n13451 = state_in[71:64] ;
assign n13452 =  ( n13451 ) == ( bv_8_214_n164 )  ;
assign n13453 = state_in[71:64] ;
assign n13454 =  ( n13453 ) == ( bv_8_213_n167 )  ;
assign n13455 = state_in[71:64] ;
assign n13456 =  ( n13455 ) == ( bv_8_212_n171 )  ;
assign n13457 = state_in[71:64] ;
assign n13458 =  ( n13457 ) == ( bv_8_211_n175 )  ;
assign n13459 = state_in[71:64] ;
assign n13460 =  ( n13459 ) == ( bv_8_210_n113 )  ;
assign n13461 = state_in[71:64] ;
assign n13462 =  ( n13461 ) == ( bv_8_209_n182 )  ;
assign n13463 = state_in[71:64] ;
assign n13464 =  ( n13463 ) == ( bv_8_208_n37 )  ;
assign n13465 = state_in[71:64] ;
assign n13466 =  ( n13465 ) == ( bv_8_207_n188 )  ;
assign n13467 = state_in[71:64] ;
assign n13468 =  ( n13467 ) == ( bv_8_206_n192 )  ;
assign n13469 = state_in[71:64] ;
assign n13470 =  ( n13469 ) == ( bv_8_205_n196 )  ;
assign n13471 = state_in[71:64] ;
assign n13472 =  ( n13471 ) == ( bv_8_204_n177 )  ;
assign n13473 = state_in[71:64] ;
assign n13474 =  ( n13473 ) == ( bv_8_203_n203 )  ;
assign n13475 = state_in[71:64] ;
assign n13476 =  ( n13475 ) == ( bv_8_202_n207 )  ;
assign n13477 = state_in[71:64] ;
assign n13478 =  ( n13477 ) == ( bv_8_201_n85 )  ;
assign n13479 = state_in[71:64] ;
assign n13480 =  ( n13479 ) == ( bv_8_200_n213 )  ;
assign n13481 = state_in[71:64] ;
assign n13482 =  ( n13481 ) == ( bv_8_199_n216 )  ;
assign n13483 = state_in[71:64] ;
assign n13484 =  ( n13483 ) == ( bv_8_198_n220 )  ;
assign n13485 = state_in[71:64] ;
assign n13486 =  ( n13485 ) == ( bv_8_197_n224 )  ;
assign n13487 = state_in[71:64] ;
assign n13488 =  ( n13487 ) == ( bv_8_196_n228 )  ;
assign n13489 = state_in[71:64] ;
assign n13490 =  ( n13489 ) == ( bv_8_195_n232 )  ;
assign n13491 = state_in[71:64] ;
assign n13492 =  ( n13491 ) == ( bv_8_194_n159 )  ;
assign n13493 = state_in[71:64] ;
assign n13494 =  ( n13493 ) == ( bv_8_193_n239 )  ;
assign n13495 = state_in[71:64] ;
assign n13496 =  ( n13495 ) == ( bv_8_192_n242 )  ;
assign n13497 = state_in[71:64] ;
assign n13498 =  ( n13497 ) == ( bv_8_191_n246 )  ;
assign n13499 = state_in[71:64] ;
assign n13500 =  ( n13499 ) == ( bv_8_190_n250 )  ;
assign n13501 = state_in[71:64] ;
assign n13502 =  ( n13501 ) == ( bv_8_189_n254 )  ;
assign n13503 = state_in[71:64] ;
assign n13504 =  ( n13503 ) == ( bv_8_188_n257 )  ;
assign n13505 = state_in[71:64] ;
assign n13506 =  ( n13505 ) == ( bv_8_187_n260 )  ;
assign n13507 = state_in[71:64] ;
assign n13508 =  ( n13507 ) == ( bv_8_186_n263 )  ;
assign n13509 = state_in[71:64] ;
assign n13510 =  ( n13509 ) == ( bv_8_185_n266 )  ;
assign n13511 = state_in[71:64] ;
assign n13512 =  ( n13511 ) == ( bv_8_184_n270 )  ;
assign n13513 = state_in[71:64] ;
assign n13514 =  ( n13513 ) == ( bv_8_183_n273 )  ;
assign n13515 = state_in[71:64] ;
assign n13516 =  ( n13515 ) == ( bv_8_182_n277 )  ;
assign n13517 = state_in[71:64] ;
assign n13518 =  ( n13517 ) == ( bv_8_181_n281 )  ;
assign n13519 = state_in[71:64] ;
assign n13520 =  ( n13519 ) == ( bv_8_180_n285 )  ;
assign n13521 = state_in[71:64] ;
assign n13522 =  ( n13521 ) == ( bv_8_179_n289 )  ;
assign n13523 = state_in[71:64] ;
assign n13524 =  ( n13523 ) == ( bv_8_178_n292 )  ;
assign n13525 = state_in[71:64] ;
assign n13526 =  ( n13525 ) == ( bv_8_177_n283 )  ;
assign n13527 = state_in[71:64] ;
assign n13528 =  ( n13527 ) == ( bv_8_176_n299 )  ;
assign n13529 = state_in[71:64] ;
assign n13530 =  ( n13529 ) == ( bv_8_175_n302 )  ;
assign n13531 = state_in[71:64] ;
assign n13532 =  ( n13531 ) == ( bv_8_174_n152 )  ;
assign n13533 = state_in[71:64] ;
assign n13534 =  ( n13533 ) == ( bv_8_173_n307 )  ;
assign n13535 = state_in[71:64] ;
assign n13536 =  ( n13535 ) == ( bv_8_172_n268 )  ;
assign n13537 = state_in[71:64] ;
assign n13538 =  ( n13537 ) == ( bv_8_171_n314 )  ;
assign n13539 = state_in[71:64] ;
assign n13540 =  ( n13539 ) == ( bv_8_170_n77 )  ;
assign n13541 = state_in[71:64] ;
assign n13542 =  ( n13541 ) == ( bv_8_169_n109 )  ;
assign n13543 = state_in[71:64] ;
assign n13544 =  ( n13543 ) == ( bv_8_168_n13 )  ;
assign n13545 = state_in[71:64] ;
assign n13546 =  ( n13545 ) == ( bv_8_167_n325 )  ;
assign n13547 = state_in[71:64] ;
assign n13548 =  ( n13547 ) == ( bv_8_166_n328 )  ;
assign n13549 = state_in[71:64] ;
assign n13550 =  ( n13549 ) == ( bv_8_165_n69 )  ;
assign n13551 = state_in[71:64] ;
assign n13552 =  ( n13551 ) == ( bv_8_164_n335 )  ;
assign n13553 = state_in[71:64] ;
assign n13554 =  ( n13553 ) == ( bv_8_163_n339 )  ;
assign n13555 = state_in[71:64] ;
assign n13556 =  ( n13555 ) == ( bv_8_162_n343 )  ;
assign n13557 = state_in[71:64] ;
assign n13558 =  ( n13557 ) == ( bv_8_161_n211 )  ;
assign n13559 = state_in[71:64] ;
assign n13560 =  ( n13559 ) == ( bv_8_160_n350 )  ;
assign n13561 = state_in[71:64] ;
assign n13562 =  ( n13561 ) == ( bv_8_159_n323 )  ;
assign n13563 = state_in[71:64] ;
assign n13564 =  ( n13563 ) == ( bv_8_158_n355 )  ;
assign n13565 = state_in[71:64] ;
assign n13566 =  ( n13565 ) == ( bv_8_157_n359 )  ;
assign n13567 = state_in[71:64] ;
assign n13568 =  ( n13567 ) == ( bv_8_156_n279 )  ;
assign n13569 = state_in[71:64] ;
assign n13570 =  ( n13569 ) == ( bv_8_155_n364 )  ;
assign n13571 = state_in[71:64] ;
assign n13572 =  ( n13571 ) == ( bv_8_154_n368 )  ;
assign n13573 = state_in[71:64] ;
assign n13574 =  ( n13573 ) == ( bv_8_153_n140 )  ;
assign n13575 = state_in[71:64] ;
assign n13576 =  ( n13575 ) == ( bv_8_152_n374 )  ;
assign n13577 = state_in[71:64] ;
assign n13578 =  ( n13577 ) == ( bv_8_151_n218 )  ;
assign n13579 = state_in[71:64] ;
assign n13580 =  ( n13579 ) == ( bv_8_150_n201 )  ;
assign n13581 = state_in[71:64] ;
assign n13582 =  ( n13581 ) == ( bv_8_149_n384 )  ;
assign n13583 = state_in[71:64] ;
assign n13584 =  ( n13583 ) == ( bv_8_148_n388 )  ;
assign n13585 = state_in[71:64] ;
assign n13586 =  ( n13585 ) == ( bv_8_147_n392 )  ;
assign n13587 = state_in[71:64] ;
assign n13588 =  ( n13587 ) == ( bv_8_146_n337 )  ;
assign n13589 = state_in[71:64] ;
assign n13590 =  ( n13589 ) == ( bv_8_145_n397 )  ;
assign n13591 = state_in[71:64] ;
assign n13592 =  ( n13591 ) == ( bv_8_144_n173 )  ;
assign n13593 = state_in[71:64] ;
assign n13594 =  ( n13593 ) == ( bv_8_143_n403 )  ;
assign n13595 = state_in[71:64] ;
assign n13596 =  ( n13595 ) == ( bv_8_142_n406 )  ;
assign n13597 = state_in[71:64] ;
assign n13598 =  ( n13597 ) == ( bv_8_141_n410 )  ;
assign n13599 = state_in[71:64] ;
assign n13600 =  ( n13599 ) == ( bv_8_140_n376 )  ;
assign n13601 = state_in[71:64] ;
assign n13602 =  ( n13601 ) == ( bv_8_139_n297 )  ;
assign n13603 = state_in[71:64] ;
assign n13604 =  ( n13603 ) == ( bv_8_138_n418 )  ;
assign n13605 = state_in[71:64] ;
assign n13606 =  ( n13605 ) == ( bv_8_137_n421 )  ;
assign n13607 = state_in[71:64] ;
assign n13608 =  ( n13607 ) == ( bv_8_136_n425 )  ;
assign n13609 = state_in[71:64] ;
assign n13610 =  ( n13609 ) == ( bv_8_135_n81 )  ;
assign n13611 = state_in[71:64] ;
assign n13612 =  ( n13611 ) == ( bv_8_134_n431 )  ;
assign n13613 = state_in[71:64] ;
assign n13614 =  ( n13613 ) == ( bv_8_133_n434 )  ;
assign n13615 = state_in[71:64] ;
assign n13616 =  ( n13615 ) == ( bv_8_132_n41 )  ;
assign n13617 = state_in[71:64] ;
assign n13618 =  ( n13617 ) == ( bv_8_131_n440 )  ;
assign n13619 = state_in[71:64] ;
assign n13620 =  ( n13619 ) == ( bv_8_130_n33 )  ;
assign n13621 = state_in[71:64] ;
assign n13622 =  ( n13621 ) == ( bv_8_129_n446 )  ;
assign n13623 = state_in[71:64] ;
assign n13624 =  ( n13623 ) == ( bv_8_128_n450 )  ;
assign n13625 = state_in[71:64] ;
assign n13626 =  ( n13625 ) == ( bv_8_127_n453 )  ;
assign n13627 = state_in[71:64] ;
assign n13628 =  ( n13627 ) == ( bv_8_126_n456 )  ;
assign n13629 = state_in[71:64] ;
assign n13630 =  ( n13629 ) == ( bv_8_125_n459 )  ;
assign n13631 = state_in[71:64] ;
assign n13632 =  ( n13631 ) == ( bv_8_124_n184 )  ;
assign n13633 = state_in[71:64] ;
assign n13634 =  ( n13633 ) == ( bv_8_123_n17 )  ;
assign n13635 = state_in[71:64] ;
assign n13636 =  ( n13635 ) == ( bv_8_122_n416 )  ;
assign n13637 = state_in[71:64] ;
assign n13638 =  ( n13637 ) == ( bv_8_121_n470 )  ;
assign n13639 = state_in[71:64] ;
assign n13640 =  ( n13639 ) == ( bv_8_120_n474 )  ;
assign n13641 = state_in[71:64] ;
assign n13642 =  ( n13641 ) == ( bv_8_119_n472 )  ;
assign n13643 = state_in[71:64] ;
assign n13644 =  ( n13643 ) == ( bv_8_118_n480 )  ;
assign n13645 = state_in[71:64] ;
assign n13646 =  ( n13645 ) == ( bv_8_117_n484 )  ;
assign n13647 = state_in[71:64] ;
assign n13648 =  ( n13647 ) == ( bv_8_116_n345 )  ;
assign n13649 = state_in[71:64] ;
assign n13650 =  ( n13649 ) == ( bv_8_115_n222 )  ;
assign n13651 = state_in[71:64] ;
assign n13652 =  ( n13651 ) == ( bv_8_114_n494 )  ;
assign n13653 = state_in[71:64] ;
assign n13654 =  ( n13653 ) == ( bv_8_113_n180 )  ;
assign n13655 = state_in[71:64] ;
assign n13656 =  ( n13655 ) == ( bv_8_112_n482 )  ;
assign n13657 = state_in[71:64] ;
assign n13658 =  ( n13657 ) == ( bv_8_111_n244 )  ;
assign n13659 = state_in[71:64] ;
assign n13660 =  ( n13659 ) == ( bv_8_110_n294 )  ;
assign n13661 = state_in[71:64] ;
assign n13662 =  ( n13661 ) == ( bv_8_109_n9 )  ;
assign n13663 = state_in[71:64] ;
assign n13664 =  ( n13663 ) == ( bv_8_108_n510 )  ;
assign n13665 = state_in[71:64] ;
assign n13666 =  ( n13665 ) == ( bv_8_107_n370 )  ;
assign n13667 = state_in[71:64] ;
assign n13668 =  ( n13667 ) == ( bv_8_106_n155 )  ;
assign n13669 = state_in[71:64] ;
assign n13670 =  ( n13669 ) == ( bv_8_105_n148 )  ;
assign n13671 = state_in[71:64] ;
assign n13672 =  ( n13671 ) == ( bv_8_104_n520 )  ;
assign n13673 = state_in[71:64] ;
assign n13674 =  ( n13673 ) == ( bv_8_103_n523 )  ;
assign n13675 = state_in[71:64] ;
assign n13676 =  ( n13675 ) == ( bv_8_102_n527 )  ;
assign n13677 = state_in[71:64] ;
assign n13678 =  ( n13677 ) == ( bv_8_101_n49 )  ;
assign n13679 = state_in[71:64] ;
assign n13680 =  ( n13679 ) == ( bv_8_100_n348 )  ;
assign n13681 = state_in[71:64] ;
assign n13682 =  ( n13681 ) == ( bv_8_99_n476 )  ;
assign n13683 = state_in[71:64] ;
assign n13684 =  ( n13683 ) == ( bv_8_98_n536 )  ;
assign n13685 = state_in[71:64] ;
assign n13686 =  ( n13685 ) == ( bv_8_97_n198 )  ;
assign n13687 = state_in[71:64] ;
assign n13688 =  ( n13687 ) == ( bv_8_96_n542 )  ;
assign n13689 = state_in[71:64] ;
assign n13690 =  ( n13689 ) == ( bv_8_95_n545 )  ;
assign n13691 = state_in[71:64] ;
assign n13692 =  ( n13691 ) == ( bv_8_94_n548 )  ;
assign n13693 = state_in[71:64] ;
assign n13694 =  ( n13693 ) == ( bv_8_93_n498 )  ;
assign n13695 = state_in[71:64] ;
assign n13696 =  ( n13695 ) == ( bv_8_92_n234 )  ;
assign n13697 = state_in[71:64] ;
assign n13698 =  ( n13697 ) == ( bv_8_91_n555 )  ;
assign n13699 = state_in[71:64] ;
assign n13700 =  ( n13699 ) == ( bv_8_90_n25 )  ;
assign n13701 = state_in[71:64] ;
assign n13702 =  ( n13701 ) == ( bv_8_89_n61 )  ;
assign n13703 = state_in[71:64] ;
assign n13704 =  ( n13703 ) == ( bv_8_88_n562 )  ;
assign n13705 = state_in[71:64] ;
assign n13706 =  ( n13705 ) == ( bv_8_87_n226 )  ;
assign n13707 = state_in[71:64] ;
assign n13708 =  ( n13707 ) == ( bv_8_86_n567 )  ;
assign n13709 = state_in[71:64] ;
assign n13710 =  ( n13709 ) == ( bv_8_85_n423 )  ;
assign n13711 = state_in[71:64] ;
assign n13712 =  ( n13711 ) == ( bv_8_84_n386 )  ;
assign n13713 = state_in[71:64] ;
assign n13714 =  ( n13713 ) == ( bv_8_83_n575 )  ;
assign n13715 = state_in[71:64] ;
assign n13716 =  ( n13715 ) == ( bv_8_82_n578 )  ;
assign n13717 = state_in[71:64] ;
assign n13718 =  ( n13717 ) == ( bv_8_81_n582 )  ;
assign n13719 = state_in[71:64] ;
assign n13720 =  ( n13719 ) == ( bv_8_80_n73 )  ;
assign n13721 = state_in[71:64] ;
assign n13722 =  ( n13721 ) == ( bv_8_79_n538 )  ;
assign n13723 = state_in[71:64] ;
assign n13724 =  ( n13723 ) == ( bv_8_78_n590 )  ;
assign n13725 = state_in[71:64] ;
assign n13726 =  ( n13725 ) == ( bv_8_77_n593 )  ;
assign n13727 = state_in[71:64] ;
assign n13728 =  ( n13727 ) == ( bv_8_76_n596 )  ;
assign n13729 = state_in[71:64] ;
assign n13730 =  ( n13729 ) == ( bv_8_75_n503 )  ;
assign n13731 = state_in[71:64] ;
assign n13732 =  ( n13731 ) == ( bv_8_74_n237 )  ;
assign n13733 = state_in[71:64] ;
assign n13734 =  ( n13733 ) == ( bv_8_73_n275 )  ;
assign n13735 = state_in[71:64] ;
assign n13736 =  ( n13735 ) == ( bv_8_72_n330 )  ;
assign n13737 = state_in[71:64] ;
assign n13738 =  ( n13737 ) == ( bv_8_71_n252 )  ;
assign n13739 = state_in[71:64] ;
assign n13740 =  ( n13739 ) == ( bv_8_70_n609 )  ;
assign n13741 = state_in[71:64] ;
assign n13742 =  ( n13741 ) == ( bv_8_69_n612 )  ;
assign n13743 = state_in[71:64] ;
assign n13744 =  ( n13743 ) == ( bv_8_68_n390 )  ;
assign n13745 = state_in[71:64] ;
assign n13746 =  ( n13745 ) == ( bv_8_67_n318 )  ;
assign n13747 = state_in[71:64] ;
assign n13748 =  ( n13747 ) == ( bv_8_66_n466 )  ;
assign n13749 = state_in[71:64] ;
assign n13750 =  ( n13749 ) == ( bv_8_65_n623 )  ;
assign n13751 = state_in[71:64] ;
assign n13752 =  ( n13751 ) == ( bv_8_64_n573 )  ;
assign n13753 = state_in[71:64] ;
assign n13754 =  ( n13753 ) == ( bv_8_63_n489 )  ;
assign n13755 = state_in[71:64] ;
assign n13756 =  ( n13755 ) == ( bv_8_62_n205 )  ;
assign n13757 = state_in[71:64] ;
assign n13758 =  ( n13757 ) == ( bv_8_61_n634 )  ;
assign n13759 = state_in[71:64] ;
assign n13760 =  ( n13759 ) == ( bv_8_60_n93 )  ;
assign n13761 = state_in[71:64] ;
assign n13762 =  ( n13761 ) == ( bv_8_59_n382 )  ;
assign n13763 = state_in[71:64] ;
assign n13764 =  ( n13763 ) == ( bv_8_58_n136 )  ;
assign n13765 = state_in[71:64] ;
assign n13766 =  ( n13765 ) == ( bv_8_57_n312 )  ;
assign n13767 = state_in[71:64] ;
assign n13768 =  ( n13767 ) == ( bv_8_56_n230 )  ;
assign n13769 = state_in[71:64] ;
assign n13770 =  ( n13769 ) == ( bv_8_55_n650 )  ;
assign n13771 = state_in[71:64] ;
assign n13772 =  ( n13771 ) == ( bv_8_54_n616 )  ;
assign n13773 = state_in[71:64] ;
assign n13774 =  ( n13773 ) == ( bv_8_53_n436 )  ;
assign n13775 = state_in[71:64] ;
assign n13776 =  ( n13775 ) == ( bv_8_52_n619 )  ;
assign n13777 = state_in[71:64] ;
assign n13778 =  ( n13777 ) == ( bv_8_51_n101 )  ;
assign n13779 = state_in[71:64] ;
assign n13780 =  ( n13779 ) == ( bv_8_50_n408 )  ;
assign n13781 = state_in[71:64] ;
assign n13782 =  ( n13781 ) == ( bv_8_49_n309 )  ;
assign n13783 = state_in[71:64] ;
assign n13784 =  ( n13783 ) == ( bv_8_48_n660 )  ;
assign n13785 = state_in[71:64] ;
assign n13786 =  ( n13785 ) == ( bv_8_47_n652 )  ;
assign n13787 = state_in[71:64] ;
assign n13788 =  ( n13787 ) == ( bv_8_46_n429 )  ;
assign n13789 = state_in[71:64] ;
assign n13790 =  ( n13789 ) == ( bv_8_45_n97 )  ;
assign n13791 = state_in[71:64] ;
assign n13792 =  ( n13791 ) == ( bv_8_44_n5 )  ;
assign n13793 = state_in[71:64] ;
assign n13794 =  ( n13793 ) == ( bv_8_43_n121 )  ;
assign n13795 = state_in[71:64] ;
assign n13796 =  ( n13795 ) == ( bv_8_42_n672 )  ;
assign n13797 = state_in[71:64] ;
assign n13798 =  ( n13797 ) == ( bv_8_41_n29 )  ;
assign n13799 = state_in[71:64] ;
assign n13800 =  ( n13799 ) == ( bv_8_40_n366 )  ;
assign n13801 = state_in[71:64] ;
assign n13802 =  ( n13801 ) == ( bv_8_39_n132 )  ;
assign n13803 = state_in[71:64] ;
assign n13804 =  ( n13803 ) == ( bv_8_38_n444 )  ;
assign n13805 = state_in[71:64] ;
assign n13806 =  ( n13805 ) == ( bv_8_37_n506 )  ;
assign n13807 = state_in[71:64] ;
assign n13808 =  ( n13807 ) == ( bv_8_36_n645 )  ;
assign n13809 = state_in[71:64] ;
assign n13810 =  ( n13809 ) == ( bv_8_35_n696 )  ;
assign n13811 = state_in[71:64] ;
assign n13812 =  ( n13811 ) == ( bv_8_34_n117 )  ;
assign n13813 = state_in[71:64] ;
assign n13814 =  ( n13813 ) == ( bv_8_33_n486 )  ;
assign n13815 = state_in[71:64] ;
assign n13816 =  ( n13815 ) == ( bv_8_32_n463 )  ;
assign n13817 = state_in[71:64] ;
assign n13818 =  ( n13817 ) == ( bv_8_31_n705 )  ;
assign n13819 = state_in[71:64] ;
assign n13820 =  ( n13819 ) == ( bv_8_30_n21 )  ;
assign n13821 = state_in[71:64] ;
assign n13822 =  ( n13821 ) == ( bv_8_29_n625 )  ;
assign n13823 = state_in[71:64] ;
assign n13824 =  ( n13823 ) == ( bv_8_28_n162 )  ;
assign n13825 = state_in[71:64] ;
assign n13826 =  ( n13825 ) == ( bv_8_27_n642 )  ;
assign n13827 = state_in[71:64] ;
assign n13828 =  ( n13827 ) == ( bv_8_26_n53 )  ;
assign n13829 = state_in[71:64] ;
assign n13830 =  ( n13829 ) == ( bv_8_25_n399 )  ;
assign n13831 = state_in[71:64] ;
assign n13832 =  ( n13831 ) == ( bv_8_24_n448 )  ;
assign n13833 = state_in[71:64] ;
assign n13834 =  ( n13833 ) == ( bv_8_23_n144 )  ;
assign n13835 = state_in[71:64] ;
assign n13836 =  ( n13835 ) == ( bv_8_22_n357 )  ;
assign n13837 = state_in[71:64] ;
assign n13838 =  ( n13837 ) == ( bv_8_21_n89 )  ;
assign n13839 = state_in[71:64] ;
assign n13840 =  ( n13839 ) == ( bv_8_20_n341 )  ;
assign n13841 = state_in[71:64] ;
assign n13842 =  ( n13841 ) == ( bv_8_19_n588 )  ;
assign n13843 = state_in[71:64] ;
assign n13844 =  ( n13843 ) == ( bv_8_18_n628 )  ;
assign n13845 = state_in[71:64] ;
assign n13846 =  ( n13845 ) == ( bv_8_17_n525 )  ;
assign n13847 = state_in[71:64] ;
assign n13848 =  ( n13847 ) == ( bv_8_16_n248 )  ;
assign n13849 = state_in[71:64] ;
assign n13850 =  ( n13849 ) == ( bv_8_15_n190 )  ;
assign n13851 = state_in[71:64] ;
assign n13852 =  ( n13851 ) == ( bv_8_14_n648 )  ;
assign n13853 = state_in[71:64] ;
assign n13854 =  ( n13853 ) == ( bv_8_13_n194 )  ;
assign n13855 = state_in[71:64] ;
assign n13856 =  ( n13855 ) == ( bv_8_12_n333 )  ;
assign n13857 = state_in[71:64] ;
assign n13858 =  ( n13857 ) == ( bv_8_11_n379 )  ;
assign n13859 = state_in[71:64] ;
assign n13860 =  ( n13859 ) == ( bv_8_10_n655 )  ;
assign n13861 = state_in[71:64] ;
assign n13862 =  ( n13861 ) == ( bv_8_9_n57 )  ;
assign n13863 = state_in[71:64] ;
assign n13864 =  ( n13863 ) == ( bv_8_8_n669 )  ;
assign n13865 = state_in[71:64] ;
assign n13866 =  ( n13865 ) == ( bv_8_7_n105 )  ;
assign n13867 = state_in[71:64] ;
assign n13868 =  ( n13867 ) == ( bv_8_6_n169 )  ;
assign n13869 = state_in[71:64] ;
assign n13870 =  ( n13869 ) == ( bv_8_5_n492 )  ;
assign n13871 = state_in[71:64] ;
assign n13872 =  ( n13871 ) == ( bv_8_4_n516 )  ;
assign n13873 = state_in[71:64] ;
assign n13874 =  ( n13873 ) == ( bv_8_3_n65 )  ;
assign n13875 = state_in[71:64] ;
assign n13876 =  ( n13875 ) == ( bv_8_2_n751 )  ;
assign n13877 = state_in[71:64] ;
assign n13878 =  ( n13877 ) == ( bv_8_1_n287 )  ;
assign n13879 = state_in[71:64] ;
assign n13880 =  ( n13879 ) == ( bv_8_0_n580 )  ;
assign n13881 =  ( n13880 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n13882 =  ( n13878 ) ? ( bv_8_124_n184 ) : ( n13881 ) ;
assign n13883 =  ( n13876 ) ? ( bv_8_119_n472 ) : ( n13882 ) ;
assign n13884 =  ( n13874 ) ? ( bv_8_123_n17 ) : ( n13883 ) ;
assign n13885 =  ( n13872 ) ? ( bv_8_242_n55 ) : ( n13884 ) ;
assign n13886 =  ( n13870 ) ? ( bv_8_107_n370 ) : ( n13885 ) ;
assign n13887 =  ( n13868 ) ? ( bv_8_111_n244 ) : ( n13886 ) ;
assign n13888 =  ( n13866 ) ? ( bv_8_197_n224 ) : ( n13887 ) ;
assign n13889 =  ( n13864 ) ? ( bv_8_48_n660 ) : ( n13888 ) ;
assign n13890 =  ( n13862 ) ? ( bv_8_1_n287 ) : ( n13889 ) ;
assign n13891 =  ( n13860 ) ? ( bv_8_103_n523 ) : ( n13890 ) ;
assign n13892 =  ( n13858 ) ? ( bv_8_43_n121 ) : ( n13891 ) ;
assign n13893 =  ( n13856 ) ? ( bv_8_254_n7 ) : ( n13892 ) ;
assign n13894 =  ( n13854 ) ? ( bv_8_215_n45 ) : ( n13893 ) ;
assign n13895 =  ( n13852 ) ? ( bv_8_171_n314 ) : ( n13894 ) ;
assign n13896 =  ( n13850 ) ? ( bv_8_118_n480 ) : ( n13895 ) ;
assign n13897 =  ( n13848 ) ? ( bv_8_202_n207 ) : ( n13896 ) ;
assign n13898 =  ( n13846 ) ? ( bv_8_130_n33 ) : ( n13897 ) ;
assign n13899 =  ( n13844 ) ? ( bv_8_201_n85 ) : ( n13898 ) ;
assign n13900 =  ( n13842 ) ? ( bv_8_125_n459 ) : ( n13899 ) ;
assign n13901 =  ( n13840 ) ? ( bv_8_250_n23 ) : ( n13900 ) ;
assign n13902 =  ( n13838 ) ? ( bv_8_89_n61 ) : ( n13901 ) ;
assign n13903 =  ( n13836 ) ? ( bv_8_71_n252 ) : ( n13902 ) ;
assign n13904 =  ( n13834 ) ? ( bv_8_240_n63 ) : ( n13903 ) ;
assign n13905 =  ( n13832 ) ? ( bv_8_173_n307 ) : ( n13904 ) ;
assign n13906 =  ( n13830 ) ? ( bv_8_212_n171 ) : ( n13905 ) ;
assign n13907 =  ( n13828 ) ? ( bv_8_162_n343 ) : ( n13906 ) ;
assign n13908 =  ( n13826 ) ? ( bv_8_175_n302 ) : ( n13907 ) ;
assign n13909 =  ( n13824 ) ? ( bv_8_156_n279 ) : ( n13908 ) ;
assign n13910 =  ( n13822 ) ? ( bv_8_164_n335 ) : ( n13909 ) ;
assign n13911 =  ( n13820 ) ? ( bv_8_114_n494 ) : ( n13910 ) ;
assign n13912 =  ( n13818 ) ? ( bv_8_192_n242 ) : ( n13911 ) ;
assign n13913 =  ( n13816 ) ? ( bv_8_183_n273 ) : ( n13912 ) ;
assign n13914 =  ( n13814 ) ? ( bv_8_253_n11 ) : ( n13913 ) ;
assign n13915 =  ( n13812 ) ? ( bv_8_147_n392 ) : ( n13914 ) ;
assign n13916 =  ( n13810 ) ? ( bv_8_38_n444 ) : ( n13915 ) ;
assign n13917 =  ( n13808 ) ? ( bv_8_54_n616 ) : ( n13916 ) ;
assign n13918 =  ( n13806 ) ? ( bv_8_63_n489 ) : ( n13917 ) ;
assign n13919 =  ( n13804 ) ? ( bv_8_247_n35 ) : ( n13918 ) ;
assign n13920 =  ( n13802 ) ? ( bv_8_204_n177 ) : ( n13919 ) ;
assign n13921 =  ( n13800 ) ? ( bv_8_52_n619 ) : ( n13920 ) ;
assign n13922 =  ( n13798 ) ? ( bv_8_165_n69 ) : ( n13921 ) ;
assign n13923 =  ( n13796 ) ? ( bv_8_229_n107 ) : ( n13922 ) ;
assign n13924 =  ( n13794 ) ? ( bv_8_241_n59 ) : ( n13923 ) ;
assign n13925 =  ( n13792 ) ? ( bv_8_113_n180 ) : ( n13924 ) ;
assign n13926 =  ( n13790 ) ? ( bv_8_216_n157 ) : ( n13925 ) ;
assign n13927 =  ( n13788 ) ? ( bv_8_49_n309 ) : ( n13926 ) ;
assign n13928 =  ( n13786 ) ? ( bv_8_21_n89 ) : ( n13927 ) ;
assign n13929 =  ( n13784 ) ? ( bv_8_4_n516 ) : ( n13928 ) ;
assign n13930 =  ( n13782 ) ? ( bv_8_199_n216 ) : ( n13929 ) ;
assign n13931 =  ( n13780 ) ? ( bv_8_35_n696 ) : ( n13930 ) ;
assign n13932 =  ( n13778 ) ? ( bv_8_195_n232 ) : ( n13931 ) ;
assign n13933 =  ( n13776 ) ? ( bv_8_24_n448 ) : ( n13932 ) ;
assign n13934 =  ( n13774 ) ? ( bv_8_150_n201 ) : ( n13933 ) ;
assign n13935 =  ( n13772 ) ? ( bv_8_5_n492 ) : ( n13934 ) ;
assign n13936 =  ( n13770 ) ? ( bv_8_154_n368 ) : ( n13935 ) ;
assign n13937 =  ( n13768 ) ? ( bv_8_7_n105 ) : ( n13936 ) ;
assign n13938 =  ( n13766 ) ? ( bv_8_18_n628 ) : ( n13937 ) ;
assign n13939 =  ( n13764 ) ? ( bv_8_128_n450 ) : ( n13938 ) ;
assign n13940 =  ( n13762 ) ? ( bv_8_226_n119 ) : ( n13939 ) ;
assign n13941 =  ( n13760 ) ? ( bv_8_235_n83 ) : ( n13940 ) ;
assign n13942 =  ( n13758 ) ? ( bv_8_39_n132 ) : ( n13941 ) ;
assign n13943 =  ( n13756 ) ? ( bv_8_178_n292 ) : ( n13942 ) ;
assign n13944 =  ( n13754 ) ? ( bv_8_117_n484 ) : ( n13943 ) ;
assign n13945 =  ( n13752 ) ? ( bv_8_9_n57 ) : ( n13944 ) ;
assign n13946 =  ( n13750 ) ? ( bv_8_131_n440 ) : ( n13945 ) ;
assign n13947 =  ( n13748 ) ? ( bv_8_44_n5 ) : ( n13946 ) ;
assign n13948 =  ( n13746 ) ? ( bv_8_26_n53 ) : ( n13947 ) ;
assign n13949 =  ( n13744 ) ? ( bv_8_27_n642 ) : ( n13948 ) ;
assign n13950 =  ( n13742 ) ? ( bv_8_110_n294 ) : ( n13949 ) ;
assign n13951 =  ( n13740 ) ? ( bv_8_90_n25 ) : ( n13950 ) ;
assign n13952 =  ( n13738 ) ? ( bv_8_160_n350 ) : ( n13951 ) ;
assign n13953 =  ( n13736 ) ? ( bv_8_82_n578 ) : ( n13952 ) ;
assign n13954 =  ( n13734 ) ? ( bv_8_59_n382 ) : ( n13953 ) ;
assign n13955 =  ( n13732 ) ? ( bv_8_214_n164 ) : ( n13954 ) ;
assign n13956 =  ( n13730 ) ? ( bv_8_179_n289 ) : ( n13955 ) ;
assign n13957 =  ( n13728 ) ? ( bv_8_41_n29 ) : ( n13956 ) ;
assign n13958 =  ( n13726 ) ? ( bv_8_227_n115 ) : ( n13957 ) ;
assign n13959 =  ( n13724 ) ? ( bv_8_47_n652 ) : ( n13958 ) ;
assign n13960 =  ( n13722 ) ? ( bv_8_132_n41 ) : ( n13959 ) ;
assign n13961 =  ( n13720 ) ? ( bv_8_83_n575 ) : ( n13960 ) ;
assign n13962 =  ( n13718 ) ? ( bv_8_209_n182 ) : ( n13961 ) ;
assign n13963 =  ( n13716 ) ? ( bv_8_0_n580 ) : ( n13962 ) ;
assign n13964 =  ( n13714 ) ? ( bv_8_237_n75 ) : ( n13963 ) ;
assign n13965 =  ( n13712 ) ? ( bv_8_32_n463 ) : ( n13964 ) ;
assign n13966 =  ( n13710 ) ? ( bv_8_252_n15 ) : ( n13965 ) ;
assign n13967 =  ( n13708 ) ? ( bv_8_177_n283 ) : ( n13966 ) ;
assign n13968 =  ( n13706 ) ? ( bv_8_91_n555 ) : ( n13967 ) ;
assign n13969 =  ( n13704 ) ? ( bv_8_106_n155 ) : ( n13968 ) ;
assign n13970 =  ( n13702 ) ? ( bv_8_203_n203 ) : ( n13969 ) ;
assign n13971 =  ( n13700 ) ? ( bv_8_190_n250 ) : ( n13970 ) ;
assign n13972 =  ( n13698 ) ? ( bv_8_57_n312 ) : ( n13971 ) ;
assign n13973 =  ( n13696 ) ? ( bv_8_74_n237 ) : ( n13972 ) ;
assign n13974 =  ( n13694 ) ? ( bv_8_76_n596 ) : ( n13973 ) ;
assign n13975 =  ( n13692 ) ? ( bv_8_88_n562 ) : ( n13974 ) ;
assign n13976 =  ( n13690 ) ? ( bv_8_207_n188 ) : ( n13975 ) ;
assign n13977 =  ( n13688 ) ? ( bv_8_208_n37 ) : ( n13976 ) ;
assign n13978 =  ( n13686 ) ? ( bv_8_239_n67 ) : ( n13977 ) ;
assign n13979 =  ( n13684 ) ? ( bv_8_170_n77 ) : ( n13978 ) ;
assign n13980 =  ( n13682 ) ? ( bv_8_251_n19 ) : ( n13979 ) ;
assign n13981 =  ( n13680 ) ? ( bv_8_67_n318 ) : ( n13980 ) ;
assign n13982 =  ( n13678 ) ? ( bv_8_77_n593 ) : ( n13981 ) ;
assign n13983 =  ( n13676 ) ? ( bv_8_51_n101 ) : ( n13982 ) ;
assign n13984 =  ( n13674 ) ? ( bv_8_133_n434 ) : ( n13983 ) ;
assign n13985 =  ( n13672 ) ? ( bv_8_69_n612 ) : ( n13984 ) ;
assign n13986 =  ( n13670 ) ? ( bv_8_249_n27 ) : ( n13985 ) ;
assign n13987 =  ( n13668 ) ? ( bv_8_2_n751 ) : ( n13986 ) ;
assign n13988 =  ( n13666 ) ? ( bv_8_127_n453 ) : ( n13987 ) ;
assign n13989 =  ( n13664 ) ? ( bv_8_80_n73 ) : ( n13988 ) ;
assign n13990 =  ( n13662 ) ? ( bv_8_60_n93 ) : ( n13989 ) ;
assign n13991 =  ( n13660 ) ? ( bv_8_159_n323 ) : ( n13990 ) ;
assign n13992 =  ( n13658 ) ? ( bv_8_168_n13 ) : ( n13991 ) ;
assign n13993 =  ( n13656 ) ? ( bv_8_81_n582 ) : ( n13992 ) ;
assign n13994 =  ( n13654 ) ? ( bv_8_163_n339 ) : ( n13993 ) ;
assign n13995 =  ( n13652 ) ? ( bv_8_64_n573 ) : ( n13994 ) ;
assign n13996 =  ( n13650 ) ? ( bv_8_143_n403 ) : ( n13995 ) ;
assign n13997 =  ( n13648 ) ? ( bv_8_146_n337 ) : ( n13996 ) ;
assign n13998 =  ( n13646 ) ? ( bv_8_157_n359 ) : ( n13997 ) ;
assign n13999 =  ( n13644 ) ? ( bv_8_56_n230 ) : ( n13998 ) ;
assign n14000 =  ( n13642 ) ? ( bv_8_245_n43 ) : ( n13999 ) ;
assign n14001 =  ( n13640 ) ? ( bv_8_188_n257 ) : ( n14000 ) ;
assign n14002 =  ( n13638 ) ? ( bv_8_182_n277 ) : ( n14001 ) ;
assign n14003 =  ( n13636 ) ? ( bv_8_218_n150 ) : ( n14002 ) ;
assign n14004 =  ( n13634 ) ? ( bv_8_33_n486 ) : ( n14003 ) ;
assign n14005 =  ( n13632 ) ? ( bv_8_16_n248 ) : ( n14004 ) ;
assign n14006 =  ( n13630 ) ? ( bv_8_255_n3 ) : ( n14005 ) ;
assign n14007 =  ( n13628 ) ? ( bv_8_243_n51 ) : ( n14006 ) ;
assign n14008 =  ( n13626 ) ? ( bv_8_210_n113 ) : ( n14007 ) ;
assign n14009 =  ( n13624 ) ? ( bv_8_205_n196 ) : ( n14008 ) ;
assign n14010 =  ( n13622 ) ? ( bv_8_12_n333 ) : ( n14009 ) ;
assign n14011 =  ( n13620 ) ? ( bv_8_19_n588 ) : ( n14010 ) ;
assign n14012 =  ( n13618 ) ? ( bv_8_236_n79 ) : ( n14011 ) ;
assign n14013 =  ( n13616 ) ? ( bv_8_95_n545 ) : ( n14012 ) ;
assign n14014 =  ( n13614 ) ? ( bv_8_151_n218 ) : ( n14013 ) ;
assign n14015 =  ( n13612 ) ? ( bv_8_68_n390 ) : ( n14014 ) ;
assign n14016 =  ( n13610 ) ? ( bv_8_23_n144 ) : ( n14015 ) ;
assign n14017 =  ( n13608 ) ? ( bv_8_196_n228 ) : ( n14016 ) ;
assign n14018 =  ( n13606 ) ? ( bv_8_167_n325 ) : ( n14017 ) ;
assign n14019 =  ( n13604 ) ? ( bv_8_126_n456 ) : ( n14018 ) ;
assign n14020 =  ( n13602 ) ? ( bv_8_61_n634 ) : ( n14019 ) ;
assign n14021 =  ( n13600 ) ? ( bv_8_100_n348 ) : ( n14020 ) ;
assign n14022 =  ( n13598 ) ? ( bv_8_93_n498 ) : ( n14021 ) ;
assign n14023 =  ( n13596 ) ? ( bv_8_25_n399 ) : ( n14022 ) ;
assign n14024 =  ( n13594 ) ? ( bv_8_115_n222 ) : ( n14023 ) ;
assign n14025 =  ( n13592 ) ? ( bv_8_96_n542 ) : ( n14024 ) ;
assign n14026 =  ( n13590 ) ? ( bv_8_129_n446 ) : ( n14025 ) ;
assign n14027 =  ( n13588 ) ? ( bv_8_79_n538 ) : ( n14026 ) ;
assign n14028 =  ( n13586 ) ? ( bv_8_220_n142 ) : ( n14027 ) ;
assign n14029 =  ( n13584 ) ? ( bv_8_34_n117 ) : ( n14028 ) ;
assign n14030 =  ( n13582 ) ? ( bv_8_42_n672 ) : ( n14029 ) ;
assign n14031 =  ( n13580 ) ? ( bv_8_144_n173 ) : ( n14030 ) ;
assign n14032 =  ( n13578 ) ? ( bv_8_136_n425 ) : ( n14031 ) ;
assign n14033 =  ( n13576 ) ? ( bv_8_70_n609 ) : ( n14032 ) ;
assign n14034 =  ( n13574 ) ? ( bv_8_238_n71 ) : ( n14033 ) ;
assign n14035 =  ( n13572 ) ? ( bv_8_184_n270 ) : ( n14034 ) ;
assign n14036 =  ( n13570 ) ? ( bv_8_20_n341 ) : ( n14035 ) ;
assign n14037 =  ( n13568 ) ? ( bv_8_222_n134 ) : ( n14036 ) ;
assign n14038 =  ( n13566 ) ? ( bv_8_94_n548 ) : ( n14037 ) ;
assign n14039 =  ( n13564 ) ? ( bv_8_11_n379 ) : ( n14038 ) ;
assign n14040 =  ( n13562 ) ? ( bv_8_219_n146 ) : ( n14039 ) ;
assign n14041 =  ( n13560 ) ? ( bv_8_224_n126 ) : ( n14040 ) ;
assign n14042 =  ( n13558 ) ? ( bv_8_50_n408 ) : ( n14041 ) ;
assign n14043 =  ( n13556 ) ? ( bv_8_58_n136 ) : ( n14042 ) ;
assign n14044 =  ( n13554 ) ? ( bv_8_10_n655 ) : ( n14043 ) ;
assign n14045 =  ( n13552 ) ? ( bv_8_73_n275 ) : ( n14044 ) ;
assign n14046 =  ( n13550 ) ? ( bv_8_6_n169 ) : ( n14045 ) ;
assign n14047 =  ( n13548 ) ? ( bv_8_36_n645 ) : ( n14046 ) ;
assign n14048 =  ( n13546 ) ? ( bv_8_92_n234 ) : ( n14047 ) ;
assign n14049 =  ( n13544 ) ? ( bv_8_194_n159 ) : ( n14048 ) ;
assign n14050 =  ( n13542 ) ? ( bv_8_211_n175 ) : ( n14049 ) ;
assign n14051 =  ( n13540 ) ? ( bv_8_172_n268 ) : ( n14050 ) ;
assign n14052 =  ( n13538 ) ? ( bv_8_98_n536 ) : ( n14051 ) ;
assign n14053 =  ( n13536 ) ? ( bv_8_145_n397 ) : ( n14052 ) ;
assign n14054 =  ( n13534 ) ? ( bv_8_149_n384 ) : ( n14053 ) ;
assign n14055 =  ( n13532 ) ? ( bv_8_228_n111 ) : ( n14054 ) ;
assign n14056 =  ( n13530 ) ? ( bv_8_121_n470 ) : ( n14055 ) ;
assign n14057 =  ( n13528 ) ? ( bv_8_231_n99 ) : ( n14056 ) ;
assign n14058 =  ( n13526 ) ? ( bv_8_200_n213 ) : ( n14057 ) ;
assign n14059 =  ( n13524 ) ? ( bv_8_55_n650 ) : ( n14058 ) ;
assign n14060 =  ( n13522 ) ? ( bv_8_109_n9 ) : ( n14059 ) ;
assign n14061 =  ( n13520 ) ? ( bv_8_141_n410 ) : ( n14060 ) ;
assign n14062 =  ( n13518 ) ? ( bv_8_213_n167 ) : ( n14061 ) ;
assign n14063 =  ( n13516 ) ? ( bv_8_78_n590 ) : ( n14062 ) ;
assign n14064 =  ( n13514 ) ? ( bv_8_169_n109 ) : ( n14063 ) ;
assign n14065 =  ( n13512 ) ? ( bv_8_108_n510 ) : ( n14064 ) ;
assign n14066 =  ( n13510 ) ? ( bv_8_86_n567 ) : ( n14065 ) ;
assign n14067 =  ( n13508 ) ? ( bv_8_244_n47 ) : ( n14066 ) ;
assign n14068 =  ( n13506 ) ? ( bv_8_234_n87 ) : ( n14067 ) ;
assign n14069 =  ( n13504 ) ? ( bv_8_101_n49 ) : ( n14068 ) ;
assign n14070 =  ( n13502 ) ? ( bv_8_122_n416 ) : ( n14069 ) ;
assign n14071 =  ( n13500 ) ? ( bv_8_174_n152 ) : ( n14070 ) ;
assign n14072 =  ( n13498 ) ? ( bv_8_8_n669 ) : ( n14071 ) ;
assign n14073 =  ( n13496 ) ? ( bv_8_186_n263 ) : ( n14072 ) ;
assign n14074 =  ( n13494 ) ? ( bv_8_120_n474 ) : ( n14073 ) ;
assign n14075 =  ( n13492 ) ? ( bv_8_37_n506 ) : ( n14074 ) ;
assign n14076 =  ( n13490 ) ? ( bv_8_46_n429 ) : ( n14075 ) ;
assign n14077 =  ( n13488 ) ? ( bv_8_28_n162 ) : ( n14076 ) ;
assign n14078 =  ( n13486 ) ? ( bv_8_166_n328 ) : ( n14077 ) ;
assign n14079 =  ( n13484 ) ? ( bv_8_180_n285 ) : ( n14078 ) ;
assign n14080 =  ( n13482 ) ? ( bv_8_198_n220 ) : ( n14079 ) ;
assign n14081 =  ( n13480 ) ? ( bv_8_232_n95 ) : ( n14080 ) ;
assign n14082 =  ( n13478 ) ? ( bv_8_221_n138 ) : ( n14081 ) ;
assign n14083 =  ( n13476 ) ? ( bv_8_116_n345 ) : ( n14082 ) ;
assign n14084 =  ( n13474 ) ? ( bv_8_31_n705 ) : ( n14083 ) ;
assign n14085 =  ( n13472 ) ? ( bv_8_75_n503 ) : ( n14084 ) ;
assign n14086 =  ( n13470 ) ? ( bv_8_189_n254 ) : ( n14085 ) ;
assign n14087 =  ( n13468 ) ? ( bv_8_139_n297 ) : ( n14086 ) ;
assign n14088 =  ( n13466 ) ? ( bv_8_138_n418 ) : ( n14087 ) ;
assign n14089 =  ( n13464 ) ? ( bv_8_112_n482 ) : ( n14088 ) ;
assign n14090 =  ( n13462 ) ? ( bv_8_62_n205 ) : ( n14089 ) ;
assign n14091 =  ( n13460 ) ? ( bv_8_181_n281 ) : ( n14090 ) ;
assign n14092 =  ( n13458 ) ? ( bv_8_102_n527 ) : ( n14091 ) ;
assign n14093 =  ( n13456 ) ? ( bv_8_72_n330 ) : ( n14092 ) ;
assign n14094 =  ( n13454 ) ? ( bv_8_3_n65 ) : ( n14093 ) ;
assign n14095 =  ( n13452 ) ? ( bv_8_246_n39 ) : ( n14094 ) ;
assign n14096 =  ( n13450 ) ? ( bv_8_14_n648 ) : ( n14095 ) ;
assign n14097 =  ( n13448 ) ? ( bv_8_97_n198 ) : ( n14096 ) ;
assign n14098 =  ( n13446 ) ? ( bv_8_53_n436 ) : ( n14097 ) ;
assign n14099 =  ( n13444 ) ? ( bv_8_87_n226 ) : ( n14098 ) ;
assign n14100 =  ( n13442 ) ? ( bv_8_185_n266 ) : ( n14099 ) ;
assign n14101 =  ( n13440 ) ? ( bv_8_134_n431 ) : ( n14100 ) ;
assign n14102 =  ( n13438 ) ? ( bv_8_193_n239 ) : ( n14101 ) ;
assign n14103 =  ( n13436 ) ? ( bv_8_29_n625 ) : ( n14102 ) ;
assign n14104 =  ( n13434 ) ? ( bv_8_158_n355 ) : ( n14103 ) ;
assign n14105 =  ( n13432 ) ? ( bv_8_225_n123 ) : ( n14104 ) ;
assign n14106 =  ( n13430 ) ? ( bv_8_248_n31 ) : ( n14105 ) ;
assign n14107 =  ( n13428 ) ? ( bv_8_152_n374 ) : ( n14106 ) ;
assign n14108 =  ( n13426 ) ? ( bv_8_17_n525 ) : ( n14107 ) ;
assign n14109 =  ( n13424 ) ? ( bv_8_105_n148 ) : ( n14108 ) ;
assign n14110 =  ( n13422 ) ? ( bv_8_217_n128 ) : ( n14109 ) ;
assign n14111 =  ( n13420 ) ? ( bv_8_142_n406 ) : ( n14110 ) ;
assign n14112 =  ( n13418 ) ? ( bv_8_148_n388 ) : ( n14111 ) ;
assign n14113 =  ( n13416 ) ? ( bv_8_155_n364 ) : ( n14112 ) ;
assign n14114 =  ( n13414 ) ? ( bv_8_30_n21 ) : ( n14113 ) ;
assign n14115 =  ( n13412 ) ? ( bv_8_135_n81 ) : ( n14114 ) ;
assign n14116 =  ( n13410 ) ? ( bv_8_233_n91 ) : ( n14115 ) ;
assign n14117 =  ( n13408 ) ? ( bv_8_206_n192 ) : ( n14116 ) ;
assign n14118 =  ( n13406 ) ? ( bv_8_85_n423 ) : ( n14117 ) ;
assign n14119 =  ( n13404 ) ? ( bv_8_40_n366 ) : ( n14118 ) ;
assign n14120 =  ( n13402 ) ? ( bv_8_223_n130 ) : ( n14119 ) ;
assign n14121 =  ( n13400 ) ? ( bv_8_140_n376 ) : ( n14120 ) ;
assign n14122 =  ( n13398 ) ? ( bv_8_161_n211 ) : ( n14121 ) ;
assign n14123 =  ( n13396 ) ? ( bv_8_137_n421 ) : ( n14122 ) ;
assign n14124 =  ( n13394 ) ? ( bv_8_13_n194 ) : ( n14123 ) ;
assign n14125 =  ( n13392 ) ? ( bv_8_191_n246 ) : ( n14124 ) ;
assign n14126 =  ( n13390 ) ? ( bv_8_230_n103 ) : ( n14125 ) ;
assign n14127 =  ( n13388 ) ? ( bv_8_66_n466 ) : ( n14126 ) ;
assign n14128 =  ( n13386 ) ? ( bv_8_104_n520 ) : ( n14127 ) ;
assign n14129 =  ( n13384 ) ? ( bv_8_65_n623 ) : ( n14128 ) ;
assign n14130 =  ( n13382 ) ? ( bv_8_153_n140 ) : ( n14129 ) ;
assign n14131 =  ( n13380 ) ? ( bv_8_45_n97 ) : ( n14130 ) ;
assign n14132 =  ( n13378 ) ? ( bv_8_15_n190 ) : ( n14131 ) ;
assign n14133 =  ( n13376 ) ? ( bv_8_176_n299 ) : ( n14132 ) ;
assign n14134 =  ( n13374 ) ? ( bv_8_84_n386 ) : ( n14133 ) ;
assign n14135 =  ( n13372 ) ? ( bv_8_187_n260 ) : ( n14134 ) ;
assign n14136 =  ( n13370 ) ? ( bv_8_22_n357 ) : ( n14135 ) ;
assign n14137 =  ( n13368 ) ^ ( n14136 )  ;
assign n14138 = state_in[63:56] ;
assign n14139 =  ( n14138 ) == ( bv_8_255_n3 )  ;
assign n14140 = state_in[63:56] ;
assign n14141 =  ( n14140 ) == ( bv_8_254_n7 )  ;
assign n14142 = state_in[63:56] ;
assign n14143 =  ( n14142 ) == ( bv_8_253_n11 )  ;
assign n14144 = state_in[63:56] ;
assign n14145 =  ( n14144 ) == ( bv_8_252_n15 )  ;
assign n14146 = state_in[63:56] ;
assign n14147 =  ( n14146 ) == ( bv_8_251_n19 )  ;
assign n14148 = state_in[63:56] ;
assign n14149 =  ( n14148 ) == ( bv_8_250_n23 )  ;
assign n14150 = state_in[63:56] ;
assign n14151 =  ( n14150 ) == ( bv_8_249_n27 )  ;
assign n14152 = state_in[63:56] ;
assign n14153 =  ( n14152 ) == ( bv_8_248_n31 )  ;
assign n14154 = state_in[63:56] ;
assign n14155 =  ( n14154 ) == ( bv_8_247_n35 )  ;
assign n14156 = state_in[63:56] ;
assign n14157 =  ( n14156 ) == ( bv_8_246_n39 )  ;
assign n14158 = state_in[63:56] ;
assign n14159 =  ( n14158 ) == ( bv_8_245_n43 )  ;
assign n14160 = state_in[63:56] ;
assign n14161 =  ( n14160 ) == ( bv_8_244_n47 )  ;
assign n14162 = state_in[63:56] ;
assign n14163 =  ( n14162 ) == ( bv_8_243_n51 )  ;
assign n14164 = state_in[63:56] ;
assign n14165 =  ( n14164 ) == ( bv_8_242_n55 )  ;
assign n14166 = state_in[63:56] ;
assign n14167 =  ( n14166 ) == ( bv_8_241_n59 )  ;
assign n14168 = state_in[63:56] ;
assign n14169 =  ( n14168 ) == ( bv_8_240_n63 )  ;
assign n14170 = state_in[63:56] ;
assign n14171 =  ( n14170 ) == ( bv_8_239_n67 )  ;
assign n14172 = state_in[63:56] ;
assign n14173 =  ( n14172 ) == ( bv_8_238_n71 )  ;
assign n14174 = state_in[63:56] ;
assign n14175 =  ( n14174 ) == ( bv_8_237_n75 )  ;
assign n14176 = state_in[63:56] ;
assign n14177 =  ( n14176 ) == ( bv_8_236_n79 )  ;
assign n14178 = state_in[63:56] ;
assign n14179 =  ( n14178 ) == ( bv_8_235_n83 )  ;
assign n14180 = state_in[63:56] ;
assign n14181 =  ( n14180 ) == ( bv_8_234_n87 )  ;
assign n14182 = state_in[63:56] ;
assign n14183 =  ( n14182 ) == ( bv_8_233_n91 )  ;
assign n14184 = state_in[63:56] ;
assign n14185 =  ( n14184 ) == ( bv_8_232_n95 )  ;
assign n14186 = state_in[63:56] ;
assign n14187 =  ( n14186 ) == ( bv_8_231_n99 )  ;
assign n14188 = state_in[63:56] ;
assign n14189 =  ( n14188 ) == ( bv_8_230_n103 )  ;
assign n14190 = state_in[63:56] ;
assign n14191 =  ( n14190 ) == ( bv_8_229_n107 )  ;
assign n14192 = state_in[63:56] ;
assign n14193 =  ( n14192 ) == ( bv_8_228_n111 )  ;
assign n14194 = state_in[63:56] ;
assign n14195 =  ( n14194 ) == ( bv_8_227_n115 )  ;
assign n14196 = state_in[63:56] ;
assign n14197 =  ( n14196 ) == ( bv_8_226_n119 )  ;
assign n14198 = state_in[63:56] ;
assign n14199 =  ( n14198 ) == ( bv_8_225_n123 )  ;
assign n14200 = state_in[63:56] ;
assign n14201 =  ( n14200 ) == ( bv_8_224_n126 )  ;
assign n14202 = state_in[63:56] ;
assign n14203 =  ( n14202 ) == ( bv_8_223_n130 )  ;
assign n14204 = state_in[63:56] ;
assign n14205 =  ( n14204 ) == ( bv_8_222_n134 )  ;
assign n14206 = state_in[63:56] ;
assign n14207 =  ( n14206 ) == ( bv_8_221_n138 )  ;
assign n14208 = state_in[63:56] ;
assign n14209 =  ( n14208 ) == ( bv_8_220_n142 )  ;
assign n14210 = state_in[63:56] ;
assign n14211 =  ( n14210 ) == ( bv_8_219_n146 )  ;
assign n14212 = state_in[63:56] ;
assign n14213 =  ( n14212 ) == ( bv_8_218_n150 )  ;
assign n14214 = state_in[63:56] ;
assign n14215 =  ( n14214 ) == ( bv_8_217_n128 )  ;
assign n14216 = state_in[63:56] ;
assign n14217 =  ( n14216 ) == ( bv_8_216_n157 )  ;
assign n14218 = state_in[63:56] ;
assign n14219 =  ( n14218 ) == ( bv_8_215_n45 )  ;
assign n14220 = state_in[63:56] ;
assign n14221 =  ( n14220 ) == ( bv_8_214_n164 )  ;
assign n14222 = state_in[63:56] ;
assign n14223 =  ( n14222 ) == ( bv_8_213_n167 )  ;
assign n14224 = state_in[63:56] ;
assign n14225 =  ( n14224 ) == ( bv_8_212_n171 )  ;
assign n14226 = state_in[63:56] ;
assign n14227 =  ( n14226 ) == ( bv_8_211_n175 )  ;
assign n14228 = state_in[63:56] ;
assign n14229 =  ( n14228 ) == ( bv_8_210_n113 )  ;
assign n14230 = state_in[63:56] ;
assign n14231 =  ( n14230 ) == ( bv_8_209_n182 )  ;
assign n14232 = state_in[63:56] ;
assign n14233 =  ( n14232 ) == ( bv_8_208_n37 )  ;
assign n14234 = state_in[63:56] ;
assign n14235 =  ( n14234 ) == ( bv_8_207_n188 )  ;
assign n14236 = state_in[63:56] ;
assign n14237 =  ( n14236 ) == ( bv_8_206_n192 )  ;
assign n14238 = state_in[63:56] ;
assign n14239 =  ( n14238 ) == ( bv_8_205_n196 )  ;
assign n14240 = state_in[63:56] ;
assign n14241 =  ( n14240 ) == ( bv_8_204_n177 )  ;
assign n14242 = state_in[63:56] ;
assign n14243 =  ( n14242 ) == ( bv_8_203_n203 )  ;
assign n14244 = state_in[63:56] ;
assign n14245 =  ( n14244 ) == ( bv_8_202_n207 )  ;
assign n14246 = state_in[63:56] ;
assign n14247 =  ( n14246 ) == ( bv_8_201_n85 )  ;
assign n14248 = state_in[63:56] ;
assign n14249 =  ( n14248 ) == ( bv_8_200_n213 )  ;
assign n14250 = state_in[63:56] ;
assign n14251 =  ( n14250 ) == ( bv_8_199_n216 )  ;
assign n14252 = state_in[63:56] ;
assign n14253 =  ( n14252 ) == ( bv_8_198_n220 )  ;
assign n14254 = state_in[63:56] ;
assign n14255 =  ( n14254 ) == ( bv_8_197_n224 )  ;
assign n14256 = state_in[63:56] ;
assign n14257 =  ( n14256 ) == ( bv_8_196_n228 )  ;
assign n14258 = state_in[63:56] ;
assign n14259 =  ( n14258 ) == ( bv_8_195_n232 )  ;
assign n14260 = state_in[63:56] ;
assign n14261 =  ( n14260 ) == ( bv_8_194_n159 )  ;
assign n14262 = state_in[63:56] ;
assign n14263 =  ( n14262 ) == ( bv_8_193_n239 )  ;
assign n14264 = state_in[63:56] ;
assign n14265 =  ( n14264 ) == ( bv_8_192_n242 )  ;
assign n14266 = state_in[63:56] ;
assign n14267 =  ( n14266 ) == ( bv_8_191_n246 )  ;
assign n14268 = state_in[63:56] ;
assign n14269 =  ( n14268 ) == ( bv_8_190_n250 )  ;
assign n14270 = state_in[63:56] ;
assign n14271 =  ( n14270 ) == ( bv_8_189_n254 )  ;
assign n14272 = state_in[63:56] ;
assign n14273 =  ( n14272 ) == ( bv_8_188_n257 )  ;
assign n14274 = state_in[63:56] ;
assign n14275 =  ( n14274 ) == ( bv_8_187_n260 )  ;
assign n14276 = state_in[63:56] ;
assign n14277 =  ( n14276 ) == ( bv_8_186_n263 )  ;
assign n14278 = state_in[63:56] ;
assign n14279 =  ( n14278 ) == ( bv_8_185_n266 )  ;
assign n14280 = state_in[63:56] ;
assign n14281 =  ( n14280 ) == ( bv_8_184_n270 )  ;
assign n14282 = state_in[63:56] ;
assign n14283 =  ( n14282 ) == ( bv_8_183_n273 )  ;
assign n14284 = state_in[63:56] ;
assign n14285 =  ( n14284 ) == ( bv_8_182_n277 )  ;
assign n14286 = state_in[63:56] ;
assign n14287 =  ( n14286 ) == ( bv_8_181_n281 )  ;
assign n14288 = state_in[63:56] ;
assign n14289 =  ( n14288 ) == ( bv_8_180_n285 )  ;
assign n14290 = state_in[63:56] ;
assign n14291 =  ( n14290 ) == ( bv_8_179_n289 )  ;
assign n14292 = state_in[63:56] ;
assign n14293 =  ( n14292 ) == ( bv_8_178_n292 )  ;
assign n14294 = state_in[63:56] ;
assign n14295 =  ( n14294 ) == ( bv_8_177_n283 )  ;
assign n14296 = state_in[63:56] ;
assign n14297 =  ( n14296 ) == ( bv_8_176_n299 )  ;
assign n14298 = state_in[63:56] ;
assign n14299 =  ( n14298 ) == ( bv_8_175_n302 )  ;
assign n14300 = state_in[63:56] ;
assign n14301 =  ( n14300 ) == ( bv_8_174_n152 )  ;
assign n14302 = state_in[63:56] ;
assign n14303 =  ( n14302 ) == ( bv_8_173_n307 )  ;
assign n14304 = state_in[63:56] ;
assign n14305 =  ( n14304 ) == ( bv_8_172_n268 )  ;
assign n14306 = state_in[63:56] ;
assign n14307 =  ( n14306 ) == ( bv_8_171_n314 )  ;
assign n14308 = state_in[63:56] ;
assign n14309 =  ( n14308 ) == ( bv_8_170_n77 )  ;
assign n14310 = state_in[63:56] ;
assign n14311 =  ( n14310 ) == ( bv_8_169_n109 )  ;
assign n14312 = state_in[63:56] ;
assign n14313 =  ( n14312 ) == ( bv_8_168_n13 )  ;
assign n14314 = state_in[63:56] ;
assign n14315 =  ( n14314 ) == ( bv_8_167_n325 )  ;
assign n14316 = state_in[63:56] ;
assign n14317 =  ( n14316 ) == ( bv_8_166_n328 )  ;
assign n14318 = state_in[63:56] ;
assign n14319 =  ( n14318 ) == ( bv_8_165_n69 )  ;
assign n14320 = state_in[63:56] ;
assign n14321 =  ( n14320 ) == ( bv_8_164_n335 )  ;
assign n14322 = state_in[63:56] ;
assign n14323 =  ( n14322 ) == ( bv_8_163_n339 )  ;
assign n14324 = state_in[63:56] ;
assign n14325 =  ( n14324 ) == ( bv_8_162_n343 )  ;
assign n14326 = state_in[63:56] ;
assign n14327 =  ( n14326 ) == ( bv_8_161_n211 )  ;
assign n14328 = state_in[63:56] ;
assign n14329 =  ( n14328 ) == ( bv_8_160_n350 )  ;
assign n14330 = state_in[63:56] ;
assign n14331 =  ( n14330 ) == ( bv_8_159_n323 )  ;
assign n14332 = state_in[63:56] ;
assign n14333 =  ( n14332 ) == ( bv_8_158_n355 )  ;
assign n14334 = state_in[63:56] ;
assign n14335 =  ( n14334 ) == ( bv_8_157_n359 )  ;
assign n14336 = state_in[63:56] ;
assign n14337 =  ( n14336 ) == ( bv_8_156_n279 )  ;
assign n14338 = state_in[63:56] ;
assign n14339 =  ( n14338 ) == ( bv_8_155_n364 )  ;
assign n14340 = state_in[63:56] ;
assign n14341 =  ( n14340 ) == ( bv_8_154_n368 )  ;
assign n14342 = state_in[63:56] ;
assign n14343 =  ( n14342 ) == ( bv_8_153_n140 )  ;
assign n14344 = state_in[63:56] ;
assign n14345 =  ( n14344 ) == ( bv_8_152_n374 )  ;
assign n14346 = state_in[63:56] ;
assign n14347 =  ( n14346 ) == ( bv_8_151_n218 )  ;
assign n14348 = state_in[63:56] ;
assign n14349 =  ( n14348 ) == ( bv_8_150_n201 )  ;
assign n14350 = state_in[63:56] ;
assign n14351 =  ( n14350 ) == ( bv_8_149_n384 )  ;
assign n14352 = state_in[63:56] ;
assign n14353 =  ( n14352 ) == ( bv_8_148_n388 )  ;
assign n14354 = state_in[63:56] ;
assign n14355 =  ( n14354 ) == ( bv_8_147_n392 )  ;
assign n14356 = state_in[63:56] ;
assign n14357 =  ( n14356 ) == ( bv_8_146_n337 )  ;
assign n14358 = state_in[63:56] ;
assign n14359 =  ( n14358 ) == ( bv_8_145_n397 )  ;
assign n14360 = state_in[63:56] ;
assign n14361 =  ( n14360 ) == ( bv_8_144_n173 )  ;
assign n14362 = state_in[63:56] ;
assign n14363 =  ( n14362 ) == ( bv_8_143_n403 )  ;
assign n14364 = state_in[63:56] ;
assign n14365 =  ( n14364 ) == ( bv_8_142_n406 )  ;
assign n14366 = state_in[63:56] ;
assign n14367 =  ( n14366 ) == ( bv_8_141_n410 )  ;
assign n14368 = state_in[63:56] ;
assign n14369 =  ( n14368 ) == ( bv_8_140_n376 )  ;
assign n14370 = state_in[63:56] ;
assign n14371 =  ( n14370 ) == ( bv_8_139_n297 )  ;
assign n14372 = state_in[63:56] ;
assign n14373 =  ( n14372 ) == ( bv_8_138_n418 )  ;
assign n14374 = state_in[63:56] ;
assign n14375 =  ( n14374 ) == ( bv_8_137_n421 )  ;
assign n14376 = state_in[63:56] ;
assign n14377 =  ( n14376 ) == ( bv_8_136_n425 )  ;
assign n14378 = state_in[63:56] ;
assign n14379 =  ( n14378 ) == ( bv_8_135_n81 )  ;
assign n14380 = state_in[63:56] ;
assign n14381 =  ( n14380 ) == ( bv_8_134_n431 )  ;
assign n14382 = state_in[63:56] ;
assign n14383 =  ( n14382 ) == ( bv_8_133_n434 )  ;
assign n14384 = state_in[63:56] ;
assign n14385 =  ( n14384 ) == ( bv_8_132_n41 )  ;
assign n14386 = state_in[63:56] ;
assign n14387 =  ( n14386 ) == ( bv_8_131_n440 )  ;
assign n14388 = state_in[63:56] ;
assign n14389 =  ( n14388 ) == ( bv_8_130_n33 )  ;
assign n14390 = state_in[63:56] ;
assign n14391 =  ( n14390 ) == ( bv_8_129_n446 )  ;
assign n14392 = state_in[63:56] ;
assign n14393 =  ( n14392 ) == ( bv_8_128_n450 )  ;
assign n14394 = state_in[63:56] ;
assign n14395 =  ( n14394 ) == ( bv_8_127_n453 )  ;
assign n14396 = state_in[63:56] ;
assign n14397 =  ( n14396 ) == ( bv_8_126_n456 )  ;
assign n14398 = state_in[63:56] ;
assign n14399 =  ( n14398 ) == ( bv_8_125_n459 )  ;
assign n14400 = state_in[63:56] ;
assign n14401 =  ( n14400 ) == ( bv_8_124_n184 )  ;
assign n14402 = state_in[63:56] ;
assign n14403 =  ( n14402 ) == ( bv_8_123_n17 )  ;
assign n14404 = state_in[63:56] ;
assign n14405 =  ( n14404 ) == ( bv_8_122_n416 )  ;
assign n14406 = state_in[63:56] ;
assign n14407 =  ( n14406 ) == ( bv_8_121_n470 )  ;
assign n14408 = state_in[63:56] ;
assign n14409 =  ( n14408 ) == ( bv_8_120_n474 )  ;
assign n14410 = state_in[63:56] ;
assign n14411 =  ( n14410 ) == ( bv_8_119_n472 )  ;
assign n14412 = state_in[63:56] ;
assign n14413 =  ( n14412 ) == ( bv_8_118_n480 )  ;
assign n14414 = state_in[63:56] ;
assign n14415 =  ( n14414 ) == ( bv_8_117_n484 )  ;
assign n14416 = state_in[63:56] ;
assign n14417 =  ( n14416 ) == ( bv_8_116_n345 )  ;
assign n14418 = state_in[63:56] ;
assign n14419 =  ( n14418 ) == ( bv_8_115_n222 )  ;
assign n14420 = state_in[63:56] ;
assign n14421 =  ( n14420 ) == ( bv_8_114_n494 )  ;
assign n14422 = state_in[63:56] ;
assign n14423 =  ( n14422 ) == ( bv_8_113_n180 )  ;
assign n14424 = state_in[63:56] ;
assign n14425 =  ( n14424 ) == ( bv_8_112_n482 )  ;
assign n14426 = state_in[63:56] ;
assign n14427 =  ( n14426 ) == ( bv_8_111_n244 )  ;
assign n14428 = state_in[63:56] ;
assign n14429 =  ( n14428 ) == ( bv_8_110_n294 )  ;
assign n14430 = state_in[63:56] ;
assign n14431 =  ( n14430 ) == ( bv_8_109_n9 )  ;
assign n14432 = state_in[63:56] ;
assign n14433 =  ( n14432 ) == ( bv_8_108_n510 )  ;
assign n14434 = state_in[63:56] ;
assign n14435 =  ( n14434 ) == ( bv_8_107_n370 )  ;
assign n14436 = state_in[63:56] ;
assign n14437 =  ( n14436 ) == ( bv_8_106_n155 )  ;
assign n14438 = state_in[63:56] ;
assign n14439 =  ( n14438 ) == ( bv_8_105_n148 )  ;
assign n14440 = state_in[63:56] ;
assign n14441 =  ( n14440 ) == ( bv_8_104_n520 )  ;
assign n14442 = state_in[63:56] ;
assign n14443 =  ( n14442 ) == ( bv_8_103_n523 )  ;
assign n14444 = state_in[63:56] ;
assign n14445 =  ( n14444 ) == ( bv_8_102_n527 )  ;
assign n14446 = state_in[63:56] ;
assign n14447 =  ( n14446 ) == ( bv_8_101_n49 )  ;
assign n14448 = state_in[63:56] ;
assign n14449 =  ( n14448 ) == ( bv_8_100_n348 )  ;
assign n14450 = state_in[63:56] ;
assign n14451 =  ( n14450 ) == ( bv_8_99_n476 )  ;
assign n14452 = state_in[63:56] ;
assign n14453 =  ( n14452 ) == ( bv_8_98_n536 )  ;
assign n14454 = state_in[63:56] ;
assign n14455 =  ( n14454 ) == ( bv_8_97_n198 )  ;
assign n14456 = state_in[63:56] ;
assign n14457 =  ( n14456 ) == ( bv_8_96_n542 )  ;
assign n14458 = state_in[63:56] ;
assign n14459 =  ( n14458 ) == ( bv_8_95_n545 )  ;
assign n14460 = state_in[63:56] ;
assign n14461 =  ( n14460 ) == ( bv_8_94_n548 )  ;
assign n14462 = state_in[63:56] ;
assign n14463 =  ( n14462 ) == ( bv_8_93_n498 )  ;
assign n14464 = state_in[63:56] ;
assign n14465 =  ( n14464 ) == ( bv_8_92_n234 )  ;
assign n14466 = state_in[63:56] ;
assign n14467 =  ( n14466 ) == ( bv_8_91_n555 )  ;
assign n14468 = state_in[63:56] ;
assign n14469 =  ( n14468 ) == ( bv_8_90_n25 )  ;
assign n14470 = state_in[63:56] ;
assign n14471 =  ( n14470 ) == ( bv_8_89_n61 )  ;
assign n14472 = state_in[63:56] ;
assign n14473 =  ( n14472 ) == ( bv_8_88_n562 )  ;
assign n14474 = state_in[63:56] ;
assign n14475 =  ( n14474 ) == ( bv_8_87_n226 )  ;
assign n14476 = state_in[63:56] ;
assign n14477 =  ( n14476 ) == ( bv_8_86_n567 )  ;
assign n14478 = state_in[63:56] ;
assign n14479 =  ( n14478 ) == ( bv_8_85_n423 )  ;
assign n14480 = state_in[63:56] ;
assign n14481 =  ( n14480 ) == ( bv_8_84_n386 )  ;
assign n14482 = state_in[63:56] ;
assign n14483 =  ( n14482 ) == ( bv_8_83_n575 )  ;
assign n14484 = state_in[63:56] ;
assign n14485 =  ( n14484 ) == ( bv_8_82_n578 )  ;
assign n14486 = state_in[63:56] ;
assign n14487 =  ( n14486 ) == ( bv_8_81_n582 )  ;
assign n14488 = state_in[63:56] ;
assign n14489 =  ( n14488 ) == ( bv_8_80_n73 )  ;
assign n14490 = state_in[63:56] ;
assign n14491 =  ( n14490 ) == ( bv_8_79_n538 )  ;
assign n14492 = state_in[63:56] ;
assign n14493 =  ( n14492 ) == ( bv_8_78_n590 )  ;
assign n14494 = state_in[63:56] ;
assign n14495 =  ( n14494 ) == ( bv_8_77_n593 )  ;
assign n14496 = state_in[63:56] ;
assign n14497 =  ( n14496 ) == ( bv_8_76_n596 )  ;
assign n14498 = state_in[63:56] ;
assign n14499 =  ( n14498 ) == ( bv_8_75_n503 )  ;
assign n14500 = state_in[63:56] ;
assign n14501 =  ( n14500 ) == ( bv_8_74_n237 )  ;
assign n14502 = state_in[63:56] ;
assign n14503 =  ( n14502 ) == ( bv_8_73_n275 )  ;
assign n14504 = state_in[63:56] ;
assign n14505 =  ( n14504 ) == ( bv_8_72_n330 )  ;
assign n14506 = state_in[63:56] ;
assign n14507 =  ( n14506 ) == ( bv_8_71_n252 )  ;
assign n14508 = state_in[63:56] ;
assign n14509 =  ( n14508 ) == ( bv_8_70_n609 )  ;
assign n14510 = state_in[63:56] ;
assign n14511 =  ( n14510 ) == ( bv_8_69_n612 )  ;
assign n14512 = state_in[63:56] ;
assign n14513 =  ( n14512 ) == ( bv_8_68_n390 )  ;
assign n14514 = state_in[63:56] ;
assign n14515 =  ( n14514 ) == ( bv_8_67_n318 )  ;
assign n14516 = state_in[63:56] ;
assign n14517 =  ( n14516 ) == ( bv_8_66_n466 )  ;
assign n14518 = state_in[63:56] ;
assign n14519 =  ( n14518 ) == ( bv_8_65_n623 )  ;
assign n14520 = state_in[63:56] ;
assign n14521 =  ( n14520 ) == ( bv_8_64_n573 )  ;
assign n14522 = state_in[63:56] ;
assign n14523 =  ( n14522 ) == ( bv_8_63_n489 )  ;
assign n14524 = state_in[63:56] ;
assign n14525 =  ( n14524 ) == ( bv_8_62_n205 )  ;
assign n14526 = state_in[63:56] ;
assign n14527 =  ( n14526 ) == ( bv_8_61_n634 )  ;
assign n14528 = state_in[63:56] ;
assign n14529 =  ( n14528 ) == ( bv_8_60_n93 )  ;
assign n14530 = state_in[63:56] ;
assign n14531 =  ( n14530 ) == ( bv_8_59_n382 )  ;
assign n14532 = state_in[63:56] ;
assign n14533 =  ( n14532 ) == ( bv_8_58_n136 )  ;
assign n14534 = state_in[63:56] ;
assign n14535 =  ( n14534 ) == ( bv_8_57_n312 )  ;
assign n14536 = state_in[63:56] ;
assign n14537 =  ( n14536 ) == ( bv_8_56_n230 )  ;
assign n14538 = state_in[63:56] ;
assign n14539 =  ( n14538 ) == ( bv_8_55_n650 )  ;
assign n14540 = state_in[63:56] ;
assign n14541 =  ( n14540 ) == ( bv_8_54_n616 )  ;
assign n14542 = state_in[63:56] ;
assign n14543 =  ( n14542 ) == ( bv_8_53_n436 )  ;
assign n14544 = state_in[63:56] ;
assign n14545 =  ( n14544 ) == ( bv_8_52_n619 )  ;
assign n14546 = state_in[63:56] ;
assign n14547 =  ( n14546 ) == ( bv_8_51_n101 )  ;
assign n14548 = state_in[63:56] ;
assign n14549 =  ( n14548 ) == ( bv_8_50_n408 )  ;
assign n14550 = state_in[63:56] ;
assign n14551 =  ( n14550 ) == ( bv_8_49_n309 )  ;
assign n14552 = state_in[63:56] ;
assign n14553 =  ( n14552 ) == ( bv_8_48_n660 )  ;
assign n14554 = state_in[63:56] ;
assign n14555 =  ( n14554 ) == ( bv_8_47_n652 )  ;
assign n14556 = state_in[63:56] ;
assign n14557 =  ( n14556 ) == ( bv_8_46_n429 )  ;
assign n14558 = state_in[63:56] ;
assign n14559 =  ( n14558 ) == ( bv_8_45_n97 )  ;
assign n14560 = state_in[63:56] ;
assign n14561 =  ( n14560 ) == ( bv_8_44_n5 )  ;
assign n14562 = state_in[63:56] ;
assign n14563 =  ( n14562 ) == ( bv_8_43_n121 )  ;
assign n14564 = state_in[63:56] ;
assign n14565 =  ( n14564 ) == ( bv_8_42_n672 )  ;
assign n14566 = state_in[63:56] ;
assign n14567 =  ( n14566 ) == ( bv_8_41_n29 )  ;
assign n14568 = state_in[63:56] ;
assign n14569 =  ( n14568 ) == ( bv_8_40_n366 )  ;
assign n14570 = state_in[63:56] ;
assign n14571 =  ( n14570 ) == ( bv_8_39_n132 )  ;
assign n14572 = state_in[63:56] ;
assign n14573 =  ( n14572 ) == ( bv_8_38_n444 )  ;
assign n14574 = state_in[63:56] ;
assign n14575 =  ( n14574 ) == ( bv_8_37_n506 )  ;
assign n14576 = state_in[63:56] ;
assign n14577 =  ( n14576 ) == ( bv_8_36_n645 )  ;
assign n14578 = state_in[63:56] ;
assign n14579 =  ( n14578 ) == ( bv_8_35_n696 )  ;
assign n14580 = state_in[63:56] ;
assign n14581 =  ( n14580 ) == ( bv_8_34_n117 )  ;
assign n14582 = state_in[63:56] ;
assign n14583 =  ( n14582 ) == ( bv_8_33_n486 )  ;
assign n14584 = state_in[63:56] ;
assign n14585 =  ( n14584 ) == ( bv_8_32_n463 )  ;
assign n14586 = state_in[63:56] ;
assign n14587 =  ( n14586 ) == ( bv_8_31_n705 )  ;
assign n14588 = state_in[63:56] ;
assign n14589 =  ( n14588 ) == ( bv_8_30_n21 )  ;
assign n14590 = state_in[63:56] ;
assign n14591 =  ( n14590 ) == ( bv_8_29_n625 )  ;
assign n14592 = state_in[63:56] ;
assign n14593 =  ( n14592 ) == ( bv_8_28_n162 )  ;
assign n14594 = state_in[63:56] ;
assign n14595 =  ( n14594 ) == ( bv_8_27_n642 )  ;
assign n14596 = state_in[63:56] ;
assign n14597 =  ( n14596 ) == ( bv_8_26_n53 )  ;
assign n14598 = state_in[63:56] ;
assign n14599 =  ( n14598 ) == ( bv_8_25_n399 )  ;
assign n14600 = state_in[63:56] ;
assign n14601 =  ( n14600 ) == ( bv_8_24_n448 )  ;
assign n14602 = state_in[63:56] ;
assign n14603 =  ( n14602 ) == ( bv_8_23_n144 )  ;
assign n14604 = state_in[63:56] ;
assign n14605 =  ( n14604 ) == ( bv_8_22_n357 )  ;
assign n14606 = state_in[63:56] ;
assign n14607 =  ( n14606 ) == ( bv_8_21_n89 )  ;
assign n14608 = state_in[63:56] ;
assign n14609 =  ( n14608 ) == ( bv_8_20_n341 )  ;
assign n14610 = state_in[63:56] ;
assign n14611 =  ( n14610 ) == ( bv_8_19_n588 )  ;
assign n14612 = state_in[63:56] ;
assign n14613 =  ( n14612 ) == ( bv_8_18_n628 )  ;
assign n14614 = state_in[63:56] ;
assign n14615 =  ( n14614 ) == ( bv_8_17_n525 )  ;
assign n14616 = state_in[63:56] ;
assign n14617 =  ( n14616 ) == ( bv_8_16_n248 )  ;
assign n14618 = state_in[63:56] ;
assign n14619 =  ( n14618 ) == ( bv_8_15_n190 )  ;
assign n14620 = state_in[63:56] ;
assign n14621 =  ( n14620 ) == ( bv_8_14_n648 )  ;
assign n14622 = state_in[63:56] ;
assign n14623 =  ( n14622 ) == ( bv_8_13_n194 )  ;
assign n14624 = state_in[63:56] ;
assign n14625 =  ( n14624 ) == ( bv_8_12_n333 )  ;
assign n14626 = state_in[63:56] ;
assign n14627 =  ( n14626 ) == ( bv_8_11_n379 )  ;
assign n14628 = state_in[63:56] ;
assign n14629 =  ( n14628 ) == ( bv_8_10_n655 )  ;
assign n14630 = state_in[63:56] ;
assign n14631 =  ( n14630 ) == ( bv_8_9_n57 )  ;
assign n14632 = state_in[63:56] ;
assign n14633 =  ( n14632 ) == ( bv_8_8_n669 )  ;
assign n14634 = state_in[63:56] ;
assign n14635 =  ( n14634 ) == ( bv_8_7_n105 )  ;
assign n14636 = state_in[63:56] ;
assign n14637 =  ( n14636 ) == ( bv_8_6_n169 )  ;
assign n14638 = state_in[63:56] ;
assign n14639 =  ( n14638 ) == ( bv_8_5_n492 )  ;
assign n14640 = state_in[63:56] ;
assign n14641 =  ( n14640 ) == ( bv_8_4_n516 )  ;
assign n14642 = state_in[63:56] ;
assign n14643 =  ( n14642 ) == ( bv_8_3_n65 )  ;
assign n14644 = state_in[63:56] ;
assign n14645 =  ( n14644 ) == ( bv_8_2_n751 )  ;
assign n14646 = state_in[63:56] ;
assign n14647 =  ( n14646 ) == ( bv_8_1_n287 )  ;
assign n14648 = state_in[63:56] ;
assign n14649 =  ( n14648 ) == ( bv_8_0_n580 )  ;
assign n14650 =  ( n14649 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n14651 =  ( n14647 ) ? ( bv_8_248_n31 ) : ( n14650 ) ;
assign n14652 =  ( n14645 ) ? ( bv_8_238_n71 ) : ( n14651 ) ;
assign n14653 =  ( n14643 ) ? ( bv_8_246_n39 ) : ( n14652 ) ;
assign n14654 =  ( n14641 ) ? ( bv_8_255_n3 ) : ( n14653 ) ;
assign n14655 =  ( n14639 ) ? ( bv_8_214_n164 ) : ( n14654 ) ;
assign n14656 =  ( n14637 ) ? ( bv_8_222_n134 ) : ( n14655 ) ;
assign n14657 =  ( n14635 ) ? ( bv_8_145_n397 ) : ( n14656 ) ;
assign n14658 =  ( n14633 ) ? ( bv_8_96_n542 ) : ( n14657 ) ;
assign n14659 =  ( n14631 ) ? ( bv_8_2_n751 ) : ( n14658 ) ;
assign n14660 =  ( n14629 ) ? ( bv_8_206_n192 ) : ( n14659 ) ;
assign n14661 =  ( n14627 ) ? ( bv_8_86_n567 ) : ( n14660 ) ;
assign n14662 =  ( n14625 ) ? ( bv_8_231_n99 ) : ( n14661 ) ;
assign n14663 =  ( n14623 ) ? ( bv_8_181_n281 ) : ( n14662 ) ;
assign n14664 =  ( n14621 ) ? ( bv_8_77_n593 ) : ( n14663 ) ;
assign n14665 =  ( n14619 ) ? ( bv_8_236_n79 ) : ( n14664 ) ;
assign n14666 =  ( n14617 ) ? ( bv_8_143_n403 ) : ( n14665 ) ;
assign n14667 =  ( n14615 ) ? ( bv_8_31_n705 ) : ( n14666 ) ;
assign n14668 =  ( n14613 ) ? ( bv_8_137_n421 ) : ( n14667 ) ;
assign n14669 =  ( n14611 ) ? ( bv_8_250_n23 ) : ( n14668 ) ;
assign n14670 =  ( n14609 ) ? ( bv_8_239_n67 ) : ( n14669 ) ;
assign n14671 =  ( n14607 ) ? ( bv_8_178_n292 ) : ( n14670 ) ;
assign n14672 =  ( n14605 ) ? ( bv_8_142_n406 ) : ( n14671 ) ;
assign n14673 =  ( n14603 ) ? ( bv_8_251_n19 ) : ( n14672 ) ;
assign n14674 =  ( n14601 ) ? ( bv_8_65_n623 ) : ( n14673 ) ;
assign n14675 =  ( n14599 ) ? ( bv_8_179_n289 ) : ( n14674 ) ;
assign n14676 =  ( n14597 ) ? ( bv_8_95_n545 ) : ( n14675 ) ;
assign n14677 =  ( n14595 ) ? ( bv_8_69_n612 ) : ( n14676 ) ;
assign n14678 =  ( n14593 ) ? ( bv_8_35_n696 ) : ( n14677 ) ;
assign n14679 =  ( n14591 ) ? ( bv_8_83_n575 ) : ( n14678 ) ;
assign n14680 =  ( n14589 ) ? ( bv_8_228_n111 ) : ( n14679 ) ;
assign n14681 =  ( n14587 ) ? ( bv_8_155_n364 ) : ( n14680 ) ;
assign n14682 =  ( n14585 ) ? ( bv_8_117_n484 ) : ( n14681 ) ;
assign n14683 =  ( n14583 ) ? ( bv_8_225_n123 ) : ( n14682 ) ;
assign n14684 =  ( n14581 ) ? ( bv_8_61_n634 ) : ( n14683 ) ;
assign n14685 =  ( n14579 ) ? ( bv_8_76_n596 ) : ( n14684 ) ;
assign n14686 =  ( n14577 ) ? ( bv_8_108_n510 ) : ( n14685 ) ;
assign n14687 =  ( n14575 ) ? ( bv_8_126_n456 ) : ( n14686 ) ;
assign n14688 =  ( n14573 ) ? ( bv_8_245_n43 ) : ( n14687 ) ;
assign n14689 =  ( n14571 ) ? ( bv_8_131_n440 ) : ( n14688 ) ;
assign n14690 =  ( n14569 ) ? ( bv_8_104_n520 ) : ( n14689 ) ;
assign n14691 =  ( n14567 ) ? ( bv_8_81_n582 ) : ( n14690 ) ;
assign n14692 =  ( n14565 ) ? ( bv_8_209_n182 ) : ( n14691 ) ;
assign n14693 =  ( n14563 ) ? ( bv_8_249_n27 ) : ( n14692 ) ;
assign n14694 =  ( n14561 ) ? ( bv_8_226_n119 ) : ( n14693 ) ;
assign n14695 =  ( n14559 ) ? ( bv_8_171_n314 ) : ( n14694 ) ;
assign n14696 =  ( n14557 ) ? ( bv_8_98_n536 ) : ( n14695 ) ;
assign n14697 =  ( n14555 ) ? ( bv_8_42_n672 ) : ( n14696 ) ;
assign n14698 =  ( n14553 ) ? ( bv_8_8_n669 ) : ( n14697 ) ;
assign n14699 =  ( n14551 ) ? ( bv_8_149_n384 ) : ( n14698 ) ;
assign n14700 =  ( n14549 ) ? ( bv_8_70_n609 ) : ( n14699 ) ;
assign n14701 =  ( n14547 ) ? ( bv_8_157_n359 ) : ( n14700 ) ;
assign n14702 =  ( n14545 ) ? ( bv_8_48_n660 ) : ( n14701 ) ;
assign n14703 =  ( n14543 ) ? ( bv_8_55_n650 ) : ( n14702 ) ;
assign n14704 =  ( n14541 ) ? ( bv_8_10_n655 ) : ( n14703 ) ;
assign n14705 =  ( n14539 ) ? ( bv_8_47_n652 ) : ( n14704 ) ;
assign n14706 =  ( n14537 ) ? ( bv_8_14_n648 ) : ( n14705 ) ;
assign n14707 =  ( n14535 ) ? ( bv_8_36_n645 ) : ( n14706 ) ;
assign n14708 =  ( n14533 ) ? ( bv_8_27_n642 ) : ( n14707 ) ;
assign n14709 =  ( n14531 ) ? ( bv_8_223_n130 ) : ( n14708 ) ;
assign n14710 =  ( n14529 ) ? ( bv_8_205_n196 ) : ( n14709 ) ;
assign n14711 =  ( n14527 ) ? ( bv_8_78_n590 ) : ( n14710 ) ;
assign n14712 =  ( n14525 ) ? ( bv_8_127_n453 ) : ( n14711 ) ;
assign n14713 =  ( n14523 ) ? ( bv_8_234_n87 ) : ( n14712 ) ;
assign n14714 =  ( n14521 ) ? ( bv_8_18_n628 ) : ( n14713 ) ;
assign n14715 =  ( n14519 ) ? ( bv_8_29_n625 ) : ( n14714 ) ;
assign n14716 =  ( n14517 ) ? ( bv_8_88_n562 ) : ( n14715 ) ;
assign n14717 =  ( n14515 ) ? ( bv_8_52_n619 ) : ( n14716 ) ;
assign n14718 =  ( n14513 ) ? ( bv_8_54_n616 ) : ( n14717 ) ;
assign n14719 =  ( n14511 ) ? ( bv_8_220_n142 ) : ( n14718 ) ;
assign n14720 =  ( n14509 ) ? ( bv_8_180_n285 ) : ( n14719 ) ;
assign n14721 =  ( n14507 ) ? ( bv_8_91_n555 ) : ( n14720 ) ;
assign n14722 =  ( n14505 ) ? ( bv_8_164_n335 ) : ( n14721 ) ;
assign n14723 =  ( n14503 ) ? ( bv_8_118_n480 ) : ( n14722 ) ;
assign n14724 =  ( n14501 ) ? ( bv_8_183_n273 ) : ( n14723 ) ;
assign n14725 =  ( n14499 ) ? ( bv_8_125_n459 ) : ( n14724 ) ;
assign n14726 =  ( n14497 ) ? ( bv_8_82_n578 ) : ( n14725 ) ;
assign n14727 =  ( n14495 ) ? ( bv_8_221_n138 ) : ( n14726 ) ;
assign n14728 =  ( n14493 ) ? ( bv_8_94_n548 ) : ( n14727 ) ;
assign n14729 =  ( n14491 ) ? ( bv_8_19_n588 ) : ( n14728 ) ;
assign n14730 =  ( n14489 ) ? ( bv_8_166_n328 ) : ( n14729 ) ;
assign n14731 =  ( n14487 ) ? ( bv_8_185_n266 ) : ( n14730 ) ;
assign n14732 =  ( n14485 ) ? ( bv_8_0_n580 ) : ( n14731 ) ;
assign n14733 =  ( n14483 ) ? ( bv_8_193_n239 ) : ( n14732 ) ;
assign n14734 =  ( n14481 ) ? ( bv_8_64_n573 ) : ( n14733 ) ;
assign n14735 =  ( n14479 ) ? ( bv_8_227_n115 ) : ( n14734 ) ;
assign n14736 =  ( n14477 ) ? ( bv_8_121_n470 ) : ( n14735 ) ;
assign n14737 =  ( n14475 ) ? ( bv_8_182_n277 ) : ( n14736 ) ;
assign n14738 =  ( n14473 ) ? ( bv_8_212_n171 ) : ( n14737 ) ;
assign n14739 =  ( n14471 ) ? ( bv_8_141_n410 ) : ( n14738 ) ;
assign n14740 =  ( n14469 ) ? ( bv_8_103_n523 ) : ( n14739 ) ;
assign n14741 =  ( n14467 ) ? ( bv_8_114_n494 ) : ( n14740 ) ;
assign n14742 =  ( n14465 ) ? ( bv_8_148_n388 ) : ( n14741 ) ;
assign n14743 =  ( n14463 ) ? ( bv_8_152_n374 ) : ( n14742 ) ;
assign n14744 =  ( n14461 ) ? ( bv_8_176_n299 ) : ( n14743 ) ;
assign n14745 =  ( n14459 ) ? ( bv_8_133_n434 ) : ( n14744 ) ;
assign n14746 =  ( n14457 ) ? ( bv_8_187_n260 ) : ( n14745 ) ;
assign n14747 =  ( n14455 ) ? ( bv_8_197_n224 ) : ( n14746 ) ;
assign n14748 =  ( n14453 ) ? ( bv_8_79_n538 ) : ( n14747 ) ;
assign n14749 =  ( n14451 ) ? ( bv_8_237_n75 ) : ( n14748 ) ;
assign n14750 =  ( n14449 ) ? ( bv_8_134_n431 ) : ( n14749 ) ;
assign n14751 =  ( n14447 ) ? ( bv_8_154_n368 ) : ( n14750 ) ;
assign n14752 =  ( n14445 ) ? ( bv_8_102_n527 ) : ( n14751 ) ;
assign n14753 =  ( n14443 ) ? ( bv_8_17_n525 ) : ( n14752 ) ;
assign n14754 =  ( n14441 ) ? ( bv_8_138_n418 ) : ( n14753 ) ;
assign n14755 =  ( n14439 ) ? ( bv_8_233_n91 ) : ( n14754 ) ;
assign n14756 =  ( n14437 ) ? ( bv_8_4_n516 ) : ( n14755 ) ;
assign n14757 =  ( n14435 ) ? ( bv_8_254_n7 ) : ( n14756 ) ;
assign n14758 =  ( n14433 ) ? ( bv_8_160_n350 ) : ( n14757 ) ;
assign n14759 =  ( n14431 ) ? ( bv_8_120_n474 ) : ( n14758 ) ;
assign n14760 =  ( n14429 ) ? ( bv_8_37_n506 ) : ( n14759 ) ;
assign n14761 =  ( n14427 ) ? ( bv_8_75_n503 ) : ( n14760 ) ;
assign n14762 =  ( n14425 ) ? ( bv_8_162_n343 ) : ( n14761 ) ;
assign n14763 =  ( n14423 ) ? ( bv_8_93_n498 ) : ( n14762 ) ;
assign n14764 =  ( n14421 ) ? ( bv_8_128_n450 ) : ( n14763 ) ;
assign n14765 =  ( n14419 ) ? ( bv_8_5_n492 ) : ( n14764 ) ;
assign n14766 =  ( n14417 ) ? ( bv_8_63_n489 ) : ( n14765 ) ;
assign n14767 =  ( n14415 ) ? ( bv_8_33_n486 ) : ( n14766 ) ;
assign n14768 =  ( n14413 ) ? ( bv_8_112_n482 ) : ( n14767 ) ;
assign n14769 =  ( n14411 ) ? ( bv_8_241_n59 ) : ( n14768 ) ;
assign n14770 =  ( n14409 ) ? ( bv_8_99_n476 ) : ( n14769 ) ;
assign n14771 =  ( n14407 ) ? ( bv_8_119_n472 ) : ( n14770 ) ;
assign n14772 =  ( n14405 ) ? ( bv_8_175_n302 ) : ( n14771 ) ;
assign n14773 =  ( n14403 ) ? ( bv_8_66_n466 ) : ( n14772 ) ;
assign n14774 =  ( n14401 ) ? ( bv_8_32_n463 ) : ( n14773 ) ;
assign n14775 =  ( n14399 ) ? ( bv_8_229_n107 ) : ( n14774 ) ;
assign n14776 =  ( n14397 ) ? ( bv_8_253_n11 ) : ( n14775 ) ;
assign n14777 =  ( n14395 ) ? ( bv_8_191_n246 ) : ( n14776 ) ;
assign n14778 =  ( n14393 ) ? ( bv_8_129_n446 ) : ( n14777 ) ;
assign n14779 =  ( n14391 ) ? ( bv_8_24_n448 ) : ( n14778 ) ;
assign n14780 =  ( n14389 ) ? ( bv_8_38_n444 ) : ( n14779 ) ;
assign n14781 =  ( n14387 ) ? ( bv_8_195_n232 ) : ( n14780 ) ;
assign n14782 =  ( n14385 ) ? ( bv_8_190_n250 ) : ( n14781 ) ;
assign n14783 =  ( n14383 ) ? ( bv_8_53_n436 ) : ( n14782 ) ;
assign n14784 =  ( n14381 ) ? ( bv_8_136_n425 ) : ( n14783 ) ;
assign n14785 =  ( n14379 ) ? ( bv_8_46_n429 ) : ( n14784 ) ;
assign n14786 =  ( n14377 ) ? ( bv_8_147_n392 ) : ( n14785 ) ;
assign n14787 =  ( n14375 ) ? ( bv_8_85_n423 ) : ( n14786 ) ;
assign n14788 =  ( n14373 ) ? ( bv_8_252_n15 ) : ( n14787 ) ;
assign n14789 =  ( n14371 ) ? ( bv_8_122_n416 ) : ( n14788 ) ;
assign n14790 =  ( n14369 ) ? ( bv_8_200_n213 ) : ( n14789 ) ;
assign n14791 =  ( n14367 ) ? ( bv_8_186_n263 ) : ( n14790 ) ;
assign n14792 =  ( n14365 ) ? ( bv_8_50_n408 ) : ( n14791 ) ;
assign n14793 =  ( n14363 ) ? ( bv_8_230_n103 ) : ( n14792 ) ;
assign n14794 =  ( n14361 ) ? ( bv_8_192_n242 ) : ( n14793 ) ;
assign n14795 =  ( n14359 ) ? ( bv_8_25_n399 ) : ( n14794 ) ;
assign n14796 =  ( n14357 ) ? ( bv_8_158_n355 ) : ( n14795 ) ;
assign n14797 =  ( n14355 ) ? ( bv_8_163_n339 ) : ( n14796 ) ;
assign n14798 =  ( n14353 ) ? ( bv_8_68_n390 ) : ( n14797 ) ;
assign n14799 =  ( n14351 ) ? ( bv_8_84_n386 ) : ( n14798 ) ;
assign n14800 =  ( n14349 ) ? ( bv_8_59_n382 ) : ( n14799 ) ;
assign n14801 =  ( n14347 ) ? ( bv_8_11_n379 ) : ( n14800 ) ;
assign n14802 =  ( n14345 ) ? ( bv_8_140_n376 ) : ( n14801 ) ;
assign n14803 =  ( n14343 ) ? ( bv_8_199_n216 ) : ( n14802 ) ;
assign n14804 =  ( n14341 ) ? ( bv_8_107_n370 ) : ( n14803 ) ;
assign n14805 =  ( n14339 ) ? ( bv_8_40_n366 ) : ( n14804 ) ;
assign n14806 =  ( n14337 ) ? ( bv_8_167_n325 ) : ( n14805 ) ;
assign n14807 =  ( n14335 ) ? ( bv_8_188_n257 ) : ( n14806 ) ;
assign n14808 =  ( n14333 ) ? ( bv_8_22_n357 ) : ( n14807 ) ;
assign n14809 =  ( n14331 ) ? ( bv_8_173_n307 ) : ( n14808 ) ;
assign n14810 =  ( n14329 ) ? ( bv_8_219_n146 ) : ( n14809 ) ;
assign n14811 =  ( n14327 ) ? ( bv_8_100_n348 ) : ( n14810 ) ;
assign n14812 =  ( n14325 ) ? ( bv_8_116_n345 ) : ( n14811 ) ;
assign n14813 =  ( n14323 ) ? ( bv_8_20_n341 ) : ( n14812 ) ;
assign n14814 =  ( n14321 ) ? ( bv_8_146_n337 ) : ( n14813 ) ;
assign n14815 =  ( n14319 ) ? ( bv_8_12_n333 ) : ( n14814 ) ;
assign n14816 =  ( n14317 ) ? ( bv_8_72_n330 ) : ( n14815 ) ;
assign n14817 =  ( n14315 ) ? ( bv_8_184_n270 ) : ( n14816 ) ;
assign n14818 =  ( n14313 ) ? ( bv_8_159_n323 ) : ( n14817 ) ;
assign n14819 =  ( n14311 ) ? ( bv_8_189_n254 ) : ( n14818 ) ;
assign n14820 =  ( n14309 ) ? ( bv_8_67_n318 ) : ( n14819 ) ;
assign n14821 =  ( n14307 ) ? ( bv_8_196_n228 ) : ( n14820 ) ;
assign n14822 =  ( n14305 ) ? ( bv_8_57_n312 ) : ( n14821 ) ;
assign n14823 =  ( n14303 ) ? ( bv_8_49_n309 ) : ( n14822 ) ;
assign n14824 =  ( n14301 ) ? ( bv_8_211_n175 ) : ( n14823 ) ;
assign n14825 =  ( n14299 ) ? ( bv_8_242_n55 ) : ( n14824 ) ;
assign n14826 =  ( n14297 ) ? ( bv_8_213_n167 ) : ( n14825 ) ;
assign n14827 =  ( n14295 ) ? ( bv_8_139_n297 ) : ( n14826 ) ;
assign n14828 =  ( n14293 ) ? ( bv_8_110_n294 ) : ( n14827 ) ;
assign n14829 =  ( n14291 ) ? ( bv_8_218_n150 ) : ( n14828 ) ;
assign n14830 =  ( n14289 ) ? ( bv_8_1_n287 ) : ( n14829 ) ;
assign n14831 =  ( n14287 ) ? ( bv_8_177_n283 ) : ( n14830 ) ;
assign n14832 =  ( n14285 ) ? ( bv_8_156_n279 ) : ( n14831 ) ;
assign n14833 =  ( n14283 ) ? ( bv_8_73_n275 ) : ( n14832 ) ;
assign n14834 =  ( n14281 ) ? ( bv_8_216_n157 ) : ( n14833 ) ;
assign n14835 =  ( n14279 ) ? ( bv_8_172_n268 ) : ( n14834 ) ;
assign n14836 =  ( n14277 ) ? ( bv_8_243_n51 ) : ( n14835 ) ;
assign n14837 =  ( n14275 ) ? ( bv_8_207_n188 ) : ( n14836 ) ;
assign n14838 =  ( n14273 ) ? ( bv_8_202_n207 ) : ( n14837 ) ;
assign n14839 =  ( n14271 ) ? ( bv_8_244_n47 ) : ( n14838 ) ;
assign n14840 =  ( n14269 ) ? ( bv_8_71_n252 ) : ( n14839 ) ;
assign n14841 =  ( n14267 ) ? ( bv_8_16_n248 ) : ( n14840 ) ;
assign n14842 =  ( n14265 ) ? ( bv_8_111_n244 ) : ( n14841 ) ;
assign n14843 =  ( n14263 ) ? ( bv_8_240_n63 ) : ( n14842 ) ;
assign n14844 =  ( n14261 ) ? ( bv_8_74_n237 ) : ( n14843 ) ;
assign n14845 =  ( n14259 ) ? ( bv_8_92_n234 ) : ( n14844 ) ;
assign n14846 =  ( n14257 ) ? ( bv_8_56_n230 ) : ( n14845 ) ;
assign n14847 =  ( n14255 ) ? ( bv_8_87_n226 ) : ( n14846 ) ;
assign n14848 =  ( n14253 ) ? ( bv_8_115_n222 ) : ( n14847 ) ;
assign n14849 =  ( n14251 ) ? ( bv_8_151_n218 ) : ( n14848 ) ;
assign n14850 =  ( n14249 ) ? ( bv_8_203_n203 ) : ( n14849 ) ;
assign n14851 =  ( n14247 ) ? ( bv_8_161_n211 ) : ( n14850 ) ;
assign n14852 =  ( n14245 ) ? ( bv_8_232_n95 ) : ( n14851 ) ;
assign n14853 =  ( n14243 ) ? ( bv_8_62_n205 ) : ( n14852 ) ;
assign n14854 =  ( n14241 ) ? ( bv_8_150_n201 ) : ( n14853 ) ;
assign n14855 =  ( n14239 ) ? ( bv_8_97_n198 ) : ( n14854 ) ;
assign n14856 =  ( n14237 ) ? ( bv_8_13_n194 ) : ( n14855 ) ;
assign n14857 =  ( n14235 ) ? ( bv_8_15_n190 ) : ( n14856 ) ;
assign n14858 =  ( n14233 ) ? ( bv_8_224_n126 ) : ( n14857 ) ;
assign n14859 =  ( n14231 ) ? ( bv_8_124_n184 ) : ( n14858 ) ;
assign n14860 =  ( n14229 ) ? ( bv_8_113_n180 ) : ( n14859 ) ;
assign n14861 =  ( n14227 ) ? ( bv_8_204_n177 ) : ( n14860 ) ;
assign n14862 =  ( n14225 ) ? ( bv_8_144_n173 ) : ( n14861 ) ;
assign n14863 =  ( n14223 ) ? ( bv_8_6_n169 ) : ( n14862 ) ;
assign n14864 =  ( n14221 ) ? ( bv_8_247_n35 ) : ( n14863 ) ;
assign n14865 =  ( n14219 ) ? ( bv_8_28_n162 ) : ( n14864 ) ;
assign n14866 =  ( n14217 ) ? ( bv_8_194_n159 ) : ( n14865 ) ;
assign n14867 =  ( n14215 ) ? ( bv_8_106_n155 ) : ( n14866 ) ;
assign n14868 =  ( n14213 ) ? ( bv_8_174_n152 ) : ( n14867 ) ;
assign n14869 =  ( n14211 ) ? ( bv_8_105_n148 ) : ( n14868 ) ;
assign n14870 =  ( n14209 ) ? ( bv_8_23_n144 ) : ( n14869 ) ;
assign n14871 =  ( n14207 ) ? ( bv_8_153_n140 ) : ( n14870 ) ;
assign n14872 =  ( n14205 ) ? ( bv_8_58_n136 ) : ( n14871 ) ;
assign n14873 =  ( n14203 ) ? ( bv_8_39_n132 ) : ( n14872 ) ;
assign n14874 =  ( n14201 ) ? ( bv_8_217_n128 ) : ( n14873 ) ;
assign n14875 =  ( n14199 ) ? ( bv_8_235_n83 ) : ( n14874 ) ;
assign n14876 =  ( n14197 ) ? ( bv_8_43_n121 ) : ( n14875 ) ;
assign n14877 =  ( n14195 ) ? ( bv_8_34_n117 ) : ( n14876 ) ;
assign n14878 =  ( n14193 ) ? ( bv_8_210_n113 ) : ( n14877 ) ;
assign n14879 =  ( n14191 ) ? ( bv_8_169_n109 ) : ( n14878 ) ;
assign n14880 =  ( n14189 ) ? ( bv_8_7_n105 ) : ( n14879 ) ;
assign n14881 =  ( n14187 ) ? ( bv_8_51_n101 ) : ( n14880 ) ;
assign n14882 =  ( n14185 ) ? ( bv_8_45_n97 ) : ( n14881 ) ;
assign n14883 =  ( n14183 ) ? ( bv_8_60_n93 ) : ( n14882 ) ;
assign n14884 =  ( n14181 ) ? ( bv_8_21_n89 ) : ( n14883 ) ;
assign n14885 =  ( n14179 ) ? ( bv_8_201_n85 ) : ( n14884 ) ;
assign n14886 =  ( n14177 ) ? ( bv_8_135_n81 ) : ( n14885 ) ;
assign n14887 =  ( n14175 ) ? ( bv_8_170_n77 ) : ( n14886 ) ;
assign n14888 =  ( n14173 ) ? ( bv_8_80_n73 ) : ( n14887 ) ;
assign n14889 =  ( n14171 ) ? ( bv_8_165_n69 ) : ( n14888 ) ;
assign n14890 =  ( n14169 ) ? ( bv_8_3_n65 ) : ( n14889 ) ;
assign n14891 =  ( n14167 ) ? ( bv_8_89_n61 ) : ( n14890 ) ;
assign n14892 =  ( n14165 ) ? ( bv_8_9_n57 ) : ( n14891 ) ;
assign n14893 =  ( n14163 ) ? ( bv_8_26_n53 ) : ( n14892 ) ;
assign n14894 =  ( n14161 ) ? ( bv_8_101_n49 ) : ( n14893 ) ;
assign n14895 =  ( n14159 ) ? ( bv_8_215_n45 ) : ( n14894 ) ;
assign n14896 =  ( n14157 ) ? ( bv_8_132_n41 ) : ( n14895 ) ;
assign n14897 =  ( n14155 ) ? ( bv_8_208_n37 ) : ( n14896 ) ;
assign n14898 =  ( n14153 ) ? ( bv_8_130_n33 ) : ( n14897 ) ;
assign n14899 =  ( n14151 ) ? ( bv_8_41_n29 ) : ( n14898 ) ;
assign n14900 =  ( n14149 ) ? ( bv_8_90_n25 ) : ( n14899 ) ;
assign n14901 =  ( n14147 ) ? ( bv_8_30_n21 ) : ( n14900 ) ;
assign n14902 =  ( n14145 ) ? ( bv_8_123_n17 ) : ( n14901 ) ;
assign n14903 =  ( n14143 ) ? ( bv_8_168_n13 ) : ( n14902 ) ;
assign n14904 =  ( n14141 ) ? ( bv_8_109_n9 ) : ( n14903 ) ;
assign n14905 =  ( n14139 ) ? ( bv_8_44_n5 ) : ( n14904 ) ;
assign n14906 =  ( n14137 ) ^ ( n14905 )  ;
assign n14907 = state_in[23:16] ;
assign n14908 =  ( n14907 ) == ( bv_8_255_n3 )  ;
assign n14909 = state_in[23:16] ;
assign n14910 =  ( n14909 ) == ( bv_8_254_n7 )  ;
assign n14911 = state_in[23:16] ;
assign n14912 =  ( n14911 ) == ( bv_8_253_n11 )  ;
assign n14913 = state_in[23:16] ;
assign n14914 =  ( n14913 ) == ( bv_8_252_n15 )  ;
assign n14915 = state_in[23:16] ;
assign n14916 =  ( n14915 ) == ( bv_8_251_n19 )  ;
assign n14917 = state_in[23:16] ;
assign n14918 =  ( n14917 ) == ( bv_8_250_n23 )  ;
assign n14919 = state_in[23:16] ;
assign n14920 =  ( n14919 ) == ( bv_8_249_n27 )  ;
assign n14921 = state_in[23:16] ;
assign n14922 =  ( n14921 ) == ( bv_8_248_n31 )  ;
assign n14923 = state_in[23:16] ;
assign n14924 =  ( n14923 ) == ( bv_8_247_n35 )  ;
assign n14925 = state_in[23:16] ;
assign n14926 =  ( n14925 ) == ( bv_8_246_n39 )  ;
assign n14927 = state_in[23:16] ;
assign n14928 =  ( n14927 ) == ( bv_8_245_n43 )  ;
assign n14929 = state_in[23:16] ;
assign n14930 =  ( n14929 ) == ( bv_8_244_n47 )  ;
assign n14931 = state_in[23:16] ;
assign n14932 =  ( n14931 ) == ( bv_8_243_n51 )  ;
assign n14933 = state_in[23:16] ;
assign n14934 =  ( n14933 ) == ( bv_8_242_n55 )  ;
assign n14935 = state_in[23:16] ;
assign n14936 =  ( n14935 ) == ( bv_8_241_n59 )  ;
assign n14937 = state_in[23:16] ;
assign n14938 =  ( n14937 ) == ( bv_8_240_n63 )  ;
assign n14939 = state_in[23:16] ;
assign n14940 =  ( n14939 ) == ( bv_8_239_n67 )  ;
assign n14941 = state_in[23:16] ;
assign n14942 =  ( n14941 ) == ( bv_8_238_n71 )  ;
assign n14943 = state_in[23:16] ;
assign n14944 =  ( n14943 ) == ( bv_8_237_n75 )  ;
assign n14945 = state_in[23:16] ;
assign n14946 =  ( n14945 ) == ( bv_8_236_n79 )  ;
assign n14947 = state_in[23:16] ;
assign n14948 =  ( n14947 ) == ( bv_8_235_n83 )  ;
assign n14949 = state_in[23:16] ;
assign n14950 =  ( n14949 ) == ( bv_8_234_n87 )  ;
assign n14951 = state_in[23:16] ;
assign n14952 =  ( n14951 ) == ( bv_8_233_n91 )  ;
assign n14953 = state_in[23:16] ;
assign n14954 =  ( n14953 ) == ( bv_8_232_n95 )  ;
assign n14955 = state_in[23:16] ;
assign n14956 =  ( n14955 ) == ( bv_8_231_n99 )  ;
assign n14957 = state_in[23:16] ;
assign n14958 =  ( n14957 ) == ( bv_8_230_n103 )  ;
assign n14959 = state_in[23:16] ;
assign n14960 =  ( n14959 ) == ( bv_8_229_n107 )  ;
assign n14961 = state_in[23:16] ;
assign n14962 =  ( n14961 ) == ( bv_8_228_n111 )  ;
assign n14963 = state_in[23:16] ;
assign n14964 =  ( n14963 ) == ( bv_8_227_n115 )  ;
assign n14965 = state_in[23:16] ;
assign n14966 =  ( n14965 ) == ( bv_8_226_n119 )  ;
assign n14967 = state_in[23:16] ;
assign n14968 =  ( n14967 ) == ( bv_8_225_n123 )  ;
assign n14969 = state_in[23:16] ;
assign n14970 =  ( n14969 ) == ( bv_8_224_n126 )  ;
assign n14971 = state_in[23:16] ;
assign n14972 =  ( n14971 ) == ( bv_8_223_n130 )  ;
assign n14973 = state_in[23:16] ;
assign n14974 =  ( n14973 ) == ( bv_8_222_n134 )  ;
assign n14975 = state_in[23:16] ;
assign n14976 =  ( n14975 ) == ( bv_8_221_n138 )  ;
assign n14977 = state_in[23:16] ;
assign n14978 =  ( n14977 ) == ( bv_8_220_n142 )  ;
assign n14979 = state_in[23:16] ;
assign n14980 =  ( n14979 ) == ( bv_8_219_n146 )  ;
assign n14981 = state_in[23:16] ;
assign n14982 =  ( n14981 ) == ( bv_8_218_n150 )  ;
assign n14983 = state_in[23:16] ;
assign n14984 =  ( n14983 ) == ( bv_8_217_n128 )  ;
assign n14985 = state_in[23:16] ;
assign n14986 =  ( n14985 ) == ( bv_8_216_n157 )  ;
assign n14987 = state_in[23:16] ;
assign n14988 =  ( n14987 ) == ( bv_8_215_n45 )  ;
assign n14989 = state_in[23:16] ;
assign n14990 =  ( n14989 ) == ( bv_8_214_n164 )  ;
assign n14991 = state_in[23:16] ;
assign n14992 =  ( n14991 ) == ( bv_8_213_n167 )  ;
assign n14993 = state_in[23:16] ;
assign n14994 =  ( n14993 ) == ( bv_8_212_n171 )  ;
assign n14995 = state_in[23:16] ;
assign n14996 =  ( n14995 ) == ( bv_8_211_n175 )  ;
assign n14997 = state_in[23:16] ;
assign n14998 =  ( n14997 ) == ( bv_8_210_n113 )  ;
assign n14999 = state_in[23:16] ;
assign n15000 =  ( n14999 ) == ( bv_8_209_n182 )  ;
assign n15001 = state_in[23:16] ;
assign n15002 =  ( n15001 ) == ( bv_8_208_n37 )  ;
assign n15003 = state_in[23:16] ;
assign n15004 =  ( n15003 ) == ( bv_8_207_n188 )  ;
assign n15005 = state_in[23:16] ;
assign n15006 =  ( n15005 ) == ( bv_8_206_n192 )  ;
assign n15007 = state_in[23:16] ;
assign n15008 =  ( n15007 ) == ( bv_8_205_n196 )  ;
assign n15009 = state_in[23:16] ;
assign n15010 =  ( n15009 ) == ( bv_8_204_n177 )  ;
assign n15011 = state_in[23:16] ;
assign n15012 =  ( n15011 ) == ( bv_8_203_n203 )  ;
assign n15013 = state_in[23:16] ;
assign n15014 =  ( n15013 ) == ( bv_8_202_n207 )  ;
assign n15015 = state_in[23:16] ;
assign n15016 =  ( n15015 ) == ( bv_8_201_n85 )  ;
assign n15017 = state_in[23:16] ;
assign n15018 =  ( n15017 ) == ( bv_8_200_n213 )  ;
assign n15019 = state_in[23:16] ;
assign n15020 =  ( n15019 ) == ( bv_8_199_n216 )  ;
assign n15021 = state_in[23:16] ;
assign n15022 =  ( n15021 ) == ( bv_8_198_n220 )  ;
assign n15023 = state_in[23:16] ;
assign n15024 =  ( n15023 ) == ( bv_8_197_n224 )  ;
assign n15025 = state_in[23:16] ;
assign n15026 =  ( n15025 ) == ( bv_8_196_n228 )  ;
assign n15027 = state_in[23:16] ;
assign n15028 =  ( n15027 ) == ( bv_8_195_n232 )  ;
assign n15029 = state_in[23:16] ;
assign n15030 =  ( n15029 ) == ( bv_8_194_n159 )  ;
assign n15031 = state_in[23:16] ;
assign n15032 =  ( n15031 ) == ( bv_8_193_n239 )  ;
assign n15033 = state_in[23:16] ;
assign n15034 =  ( n15033 ) == ( bv_8_192_n242 )  ;
assign n15035 = state_in[23:16] ;
assign n15036 =  ( n15035 ) == ( bv_8_191_n246 )  ;
assign n15037 = state_in[23:16] ;
assign n15038 =  ( n15037 ) == ( bv_8_190_n250 )  ;
assign n15039 = state_in[23:16] ;
assign n15040 =  ( n15039 ) == ( bv_8_189_n254 )  ;
assign n15041 = state_in[23:16] ;
assign n15042 =  ( n15041 ) == ( bv_8_188_n257 )  ;
assign n15043 = state_in[23:16] ;
assign n15044 =  ( n15043 ) == ( bv_8_187_n260 )  ;
assign n15045 = state_in[23:16] ;
assign n15046 =  ( n15045 ) == ( bv_8_186_n263 )  ;
assign n15047 = state_in[23:16] ;
assign n15048 =  ( n15047 ) == ( bv_8_185_n266 )  ;
assign n15049 = state_in[23:16] ;
assign n15050 =  ( n15049 ) == ( bv_8_184_n270 )  ;
assign n15051 = state_in[23:16] ;
assign n15052 =  ( n15051 ) == ( bv_8_183_n273 )  ;
assign n15053 = state_in[23:16] ;
assign n15054 =  ( n15053 ) == ( bv_8_182_n277 )  ;
assign n15055 = state_in[23:16] ;
assign n15056 =  ( n15055 ) == ( bv_8_181_n281 )  ;
assign n15057 = state_in[23:16] ;
assign n15058 =  ( n15057 ) == ( bv_8_180_n285 )  ;
assign n15059 = state_in[23:16] ;
assign n15060 =  ( n15059 ) == ( bv_8_179_n289 )  ;
assign n15061 = state_in[23:16] ;
assign n15062 =  ( n15061 ) == ( bv_8_178_n292 )  ;
assign n15063 = state_in[23:16] ;
assign n15064 =  ( n15063 ) == ( bv_8_177_n283 )  ;
assign n15065 = state_in[23:16] ;
assign n15066 =  ( n15065 ) == ( bv_8_176_n299 )  ;
assign n15067 = state_in[23:16] ;
assign n15068 =  ( n15067 ) == ( bv_8_175_n302 )  ;
assign n15069 = state_in[23:16] ;
assign n15070 =  ( n15069 ) == ( bv_8_174_n152 )  ;
assign n15071 = state_in[23:16] ;
assign n15072 =  ( n15071 ) == ( bv_8_173_n307 )  ;
assign n15073 = state_in[23:16] ;
assign n15074 =  ( n15073 ) == ( bv_8_172_n268 )  ;
assign n15075 = state_in[23:16] ;
assign n15076 =  ( n15075 ) == ( bv_8_171_n314 )  ;
assign n15077 = state_in[23:16] ;
assign n15078 =  ( n15077 ) == ( bv_8_170_n77 )  ;
assign n15079 = state_in[23:16] ;
assign n15080 =  ( n15079 ) == ( bv_8_169_n109 )  ;
assign n15081 = state_in[23:16] ;
assign n15082 =  ( n15081 ) == ( bv_8_168_n13 )  ;
assign n15083 = state_in[23:16] ;
assign n15084 =  ( n15083 ) == ( bv_8_167_n325 )  ;
assign n15085 = state_in[23:16] ;
assign n15086 =  ( n15085 ) == ( bv_8_166_n328 )  ;
assign n15087 = state_in[23:16] ;
assign n15088 =  ( n15087 ) == ( bv_8_165_n69 )  ;
assign n15089 = state_in[23:16] ;
assign n15090 =  ( n15089 ) == ( bv_8_164_n335 )  ;
assign n15091 = state_in[23:16] ;
assign n15092 =  ( n15091 ) == ( bv_8_163_n339 )  ;
assign n15093 = state_in[23:16] ;
assign n15094 =  ( n15093 ) == ( bv_8_162_n343 )  ;
assign n15095 = state_in[23:16] ;
assign n15096 =  ( n15095 ) == ( bv_8_161_n211 )  ;
assign n15097 = state_in[23:16] ;
assign n15098 =  ( n15097 ) == ( bv_8_160_n350 )  ;
assign n15099 = state_in[23:16] ;
assign n15100 =  ( n15099 ) == ( bv_8_159_n323 )  ;
assign n15101 = state_in[23:16] ;
assign n15102 =  ( n15101 ) == ( bv_8_158_n355 )  ;
assign n15103 = state_in[23:16] ;
assign n15104 =  ( n15103 ) == ( bv_8_157_n359 )  ;
assign n15105 = state_in[23:16] ;
assign n15106 =  ( n15105 ) == ( bv_8_156_n279 )  ;
assign n15107 = state_in[23:16] ;
assign n15108 =  ( n15107 ) == ( bv_8_155_n364 )  ;
assign n15109 = state_in[23:16] ;
assign n15110 =  ( n15109 ) == ( bv_8_154_n368 )  ;
assign n15111 = state_in[23:16] ;
assign n15112 =  ( n15111 ) == ( bv_8_153_n140 )  ;
assign n15113 = state_in[23:16] ;
assign n15114 =  ( n15113 ) == ( bv_8_152_n374 )  ;
assign n15115 = state_in[23:16] ;
assign n15116 =  ( n15115 ) == ( bv_8_151_n218 )  ;
assign n15117 = state_in[23:16] ;
assign n15118 =  ( n15117 ) == ( bv_8_150_n201 )  ;
assign n15119 = state_in[23:16] ;
assign n15120 =  ( n15119 ) == ( bv_8_149_n384 )  ;
assign n15121 = state_in[23:16] ;
assign n15122 =  ( n15121 ) == ( bv_8_148_n388 )  ;
assign n15123 = state_in[23:16] ;
assign n15124 =  ( n15123 ) == ( bv_8_147_n392 )  ;
assign n15125 = state_in[23:16] ;
assign n15126 =  ( n15125 ) == ( bv_8_146_n337 )  ;
assign n15127 = state_in[23:16] ;
assign n15128 =  ( n15127 ) == ( bv_8_145_n397 )  ;
assign n15129 = state_in[23:16] ;
assign n15130 =  ( n15129 ) == ( bv_8_144_n173 )  ;
assign n15131 = state_in[23:16] ;
assign n15132 =  ( n15131 ) == ( bv_8_143_n403 )  ;
assign n15133 = state_in[23:16] ;
assign n15134 =  ( n15133 ) == ( bv_8_142_n406 )  ;
assign n15135 = state_in[23:16] ;
assign n15136 =  ( n15135 ) == ( bv_8_141_n410 )  ;
assign n15137 = state_in[23:16] ;
assign n15138 =  ( n15137 ) == ( bv_8_140_n376 )  ;
assign n15139 = state_in[23:16] ;
assign n15140 =  ( n15139 ) == ( bv_8_139_n297 )  ;
assign n15141 = state_in[23:16] ;
assign n15142 =  ( n15141 ) == ( bv_8_138_n418 )  ;
assign n15143 = state_in[23:16] ;
assign n15144 =  ( n15143 ) == ( bv_8_137_n421 )  ;
assign n15145 = state_in[23:16] ;
assign n15146 =  ( n15145 ) == ( bv_8_136_n425 )  ;
assign n15147 = state_in[23:16] ;
assign n15148 =  ( n15147 ) == ( bv_8_135_n81 )  ;
assign n15149 = state_in[23:16] ;
assign n15150 =  ( n15149 ) == ( bv_8_134_n431 )  ;
assign n15151 = state_in[23:16] ;
assign n15152 =  ( n15151 ) == ( bv_8_133_n434 )  ;
assign n15153 = state_in[23:16] ;
assign n15154 =  ( n15153 ) == ( bv_8_132_n41 )  ;
assign n15155 = state_in[23:16] ;
assign n15156 =  ( n15155 ) == ( bv_8_131_n440 )  ;
assign n15157 = state_in[23:16] ;
assign n15158 =  ( n15157 ) == ( bv_8_130_n33 )  ;
assign n15159 = state_in[23:16] ;
assign n15160 =  ( n15159 ) == ( bv_8_129_n446 )  ;
assign n15161 = state_in[23:16] ;
assign n15162 =  ( n15161 ) == ( bv_8_128_n450 )  ;
assign n15163 = state_in[23:16] ;
assign n15164 =  ( n15163 ) == ( bv_8_127_n453 )  ;
assign n15165 = state_in[23:16] ;
assign n15166 =  ( n15165 ) == ( bv_8_126_n456 )  ;
assign n15167 = state_in[23:16] ;
assign n15168 =  ( n15167 ) == ( bv_8_125_n459 )  ;
assign n15169 = state_in[23:16] ;
assign n15170 =  ( n15169 ) == ( bv_8_124_n184 )  ;
assign n15171 = state_in[23:16] ;
assign n15172 =  ( n15171 ) == ( bv_8_123_n17 )  ;
assign n15173 = state_in[23:16] ;
assign n15174 =  ( n15173 ) == ( bv_8_122_n416 )  ;
assign n15175 = state_in[23:16] ;
assign n15176 =  ( n15175 ) == ( bv_8_121_n470 )  ;
assign n15177 = state_in[23:16] ;
assign n15178 =  ( n15177 ) == ( bv_8_120_n474 )  ;
assign n15179 = state_in[23:16] ;
assign n15180 =  ( n15179 ) == ( bv_8_119_n472 )  ;
assign n15181 = state_in[23:16] ;
assign n15182 =  ( n15181 ) == ( bv_8_118_n480 )  ;
assign n15183 = state_in[23:16] ;
assign n15184 =  ( n15183 ) == ( bv_8_117_n484 )  ;
assign n15185 = state_in[23:16] ;
assign n15186 =  ( n15185 ) == ( bv_8_116_n345 )  ;
assign n15187 = state_in[23:16] ;
assign n15188 =  ( n15187 ) == ( bv_8_115_n222 )  ;
assign n15189 = state_in[23:16] ;
assign n15190 =  ( n15189 ) == ( bv_8_114_n494 )  ;
assign n15191 = state_in[23:16] ;
assign n15192 =  ( n15191 ) == ( bv_8_113_n180 )  ;
assign n15193 = state_in[23:16] ;
assign n15194 =  ( n15193 ) == ( bv_8_112_n482 )  ;
assign n15195 = state_in[23:16] ;
assign n15196 =  ( n15195 ) == ( bv_8_111_n244 )  ;
assign n15197 = state_in[23:16] ;
assign n15198 =  ( n15197 ) == ( bv_8_110_n294 )  ;
assign n15199 = state_in[23:16] ;
assign n15200 =  ( n15199 ) == ( bv_8_109_n9 )  ;
assign n15201 = state_in[23:16] ;
assign n15202 =  ( n15201 ) == ( bv_8_108_n510 )  ;
assign n15203 = state_in[23:16] ;
assign n15204 =  ( n15203 ) == ( bv_8_107_n370 )  ;
assign n15205 = state_in[23:16] ;
assign n15206 =  ( n15205 ) == ( bv_8_106_n155 )  ;
assign n15207 = state_in[23:16] ;
assign n15208 =  ( n15207 ) == ( bv_8_105_n148 )  ;
assign n15209 = state_in[23:16] ;
assign n15210 =  ( n15209 ) == ( bv_8_104_n520 )  ;
assign n15211 = state_in[23:16] ;
assign n15212 =  ( n15211 ) == ( bv_8_103_n523 )  ;
assign n15213 = state_in[23:16] ;
assign n15214 =  ( n15213 ) == ( bv_8_102_n527 )  ;
assign n15215 = state_in[23:16] ;
assign n15216 =  ( n15215 ) == ( bv_8_101_n49 )  ;
assign n15217 = state_in[23:16] ;
assign n15218 =  ( n15217 ) == ( bv_8_100_n348 )  ;
assign n15219 = state_in[23:16] ;
assign n15220 =  ( n15219 ) == ( bv_8_99_n476 )  ;
assign n15221 = state_in[23:16] ;
assign n15222 =  ( n15221 ) == ( bv_8_98_n536 )  ;
assign n15223 = state_in[23:16] ;
assign n15224 =  ( n15223 ) == ( bv_8_97_n198 )  ;
assign n15225 = state_in[23:16] ;
assign n15226 =  ( n15225 ) == ( bv_8_96_n542 )  ;
assign n15227 = state_in[23:16] ;
assign n15228 =  ( n15227 ) == ( bv_8_95_n545 )  ;
assign n15229 = state_in[23:16] ;
assign n15230 =  ( n15229 ) == ( bv_8_94_n548 )  ;
assign n15231 = state_in[23:16] ;
assign n15232 =  ( n15231 ) == ( bv_8_93_n498 )  ;
assign n15233 = state_in[23:16] ;
assign n15234 =  ( n15233 ) == ( bv_8_92_n234 )  ;
assign n15235 = state_in[23:16] ;
assign n15236 =  ( n15235 ) == ( bv_8_91_n555 )  ;
assign n15237 = state_in[23:16] ;
assign n15238 =  ( n15237 ) == ( bv_8_90_n25 )  ;
assign n15239 = state_in[23:16] ;
assign n15240 =  ( n15239 ) == ( bv_8_89_n61 )  ;
assign n15241 = state_in[23:16] ;
assign n15242 =  ( n15241 ) == ( bv_8_88_n562 )  ;
assign n15243 = state_in[23:16] ;
assign n15244 =  ( n15243 ) == ( bv_8_87_n226 )  ;
assign n15245 = state_in[23:16] ;
assign n15246 =  ( n15245 ) == ( bv_8_86_n567 )  ;
assign n15247 = state_in[23:16] ;
assign n15248 =  ( n15247 ) == ( bv_8_85_n423 )  ;
assign n15249 = state_in[23:16] ;
assign n15250 =  ( n15249 ) == ( bv_8_84_n386 )  ;
assign n15251 = state_in[23:16] ;
assign n15252 =  ( n15251 ) == ( bv_8_83_n575 )  ;
assign n15253 = state_in[23:16] ;
assign n15254 =  ( n15253 ) == ( bv_8_82_n578 )  ;
assign n15255 = state_in[23:16] ;
assign n15256 =  ( n15255 ) == ( bv_8_81_n582 )  ;
assign n15257 = state_in[23:16] ;
assign n15258 =  ( n15257 ) == ( bv_8_80_n73 )  ;
assign n15259 = state_in[23:16] ;
assign n15260 =  ( n15259 ) == ( bv_8_79_n538 )  ;
assign n15261 = state_in[23:16] ;
assign n15262 =  ( n15261 ) == ( bv_8_78_n590 )  ;
assign n15263 = state_in[23:16] ;
assign n15264 =  ( n15263 ) == ( bv_8_77_n593 )  ;
assign n15265 = state_in[23:16] ;
assign n15266 =  ( n15265 ) == ( bv_8_76_n596 )  ;
assign n15267 = state_in[23:16] ;
assign n15268 =  ( n15267 ) == ( bv_8_75_n503 )  ;
assign n15269 = state_in[23:16] ;
assign n15270 =  ( n15269 ) == ( bv_8_74_n237 )  ;
assign n15271 = state_in[23:16] ;
assign n15272 =  ( n15271 ) == ( bv_8_73_n275 )  ;
assign n15273 = state_in[23:16] ;
assign n15274 =  ( n15273 ) == ( bv_8_72_n330 )  ;
assign n15275 = state_in[23:16] ;
assign n15276 =  ( n15275 ) == ( bv_8_71_n252 )  ;
assign n15277 = state_in[23:16] ;
assign n15278 =  ( n15277 ) == ( bv_8_70_n609 )  ;
assign n15279 = state_in[23:16] ;
assign n15280 =  ( n15279 ) == ( bv_8_69_n612 )  ;
assign n15281 = state_in[23:16] ;
assign n15282 =  ( n15281 ) == ( bv_8_68_n390 )  ;
assign n15283 = state_in[23:16] ;
assign n15284 =  ( n15283 ) == ( bv_8_67_n318 )  ;
assign n15285 = state_in[23:16] ;
assign n15286 =  ( n15285 ) == ( bv_8_66_n466 )  ;
assign n15287 = state_in[23:16] ;
assign n15288 =  ( n15287 ) == ( bv_8_65_n623 )  ;
assign n15289 = state_in[23:16] ;
assign n15290 =  ( n15289 ) == ( bv_8_64_n573 )  ;
assign n15291 = state_in[23:16] ;
assign n15292 =  ( n15291 ) == ( bv_8_63_n489 )  ;
assign n15293 = state_in[23:16] ;
assign n15294 =  ( n15293 ) == ( bv_8_62_n205 )  ;
assign n15295 = state_in[23:16] ;
assign n15296 =  ( n15295 ) == ( bv_8_61_n634 )  ;
assign n15297 = state_in[23:16] ;
assign n15298 =  ( n15297 ) == ( bv_8_60_n93 )  ;
assign n15299 = state_in[23:16] ;
assign n15300 =  ( n15299 ) == ( bv_8_59_n382 )  ;
assign n15301 = state_in[23:16] ;
assign n15302 =  ( n15301 ) == ( bv_8_58_n136 )  ;
assign n15303 = state_in[23:16] ;
assign n15304 =  ( n15303 ) == ( bv_8_57_n312 )  ;
assign n15305 = state_in[23:16] ;
assign n15306 =  ( n15305 ) == ( bv_8_56_n230 )  ;
assign n15307 = state_in[23:16] ;
assign n15308 =  ( n15307 ) == ( bv_8_55_n650 )  ;
assign n15309 = state_in[23:16] ;
assign n15310 =  ( n15309 ) == ( bv_8_54_n616 )  ;
assign n15311 = state_in[23:16] ;
assign n15312 =  ( n15311 ) == ( bv_8_53_n436 )  ;
assign n15313 = state_in[23:16] ;
assign n15314 =  ( n15313 ) == ( bv_8_52_n619 )  ;
assign n15315 = state_in[23:16] ;
assign n15316 =  ( n15315 ) == ( bv_8_51_n101 )  ;
assign n15317 = state_in[23:16] ;
assign n15318 =  ( n15317 ) == ( bv_8_50_n408 )  ;
assign n15319 = state_in[23:16] ;
assign n15320 =  ( n15319 ) == ( bv_8_49_n309 )  ;
assign n15321 = state_in[23:16] ;
assign n15322 =  ( n15321 ) == ( bv_8_48_n660 )  ;
assign n15323 = state_in[23:16] ;
assign n15324 =  ( n15323 ) == ( bv_8_47_n652 )  ;
assign n15325 = state_in[23:16] ;
assign n15326 =  ( n15325 ) == ( bv_8_46_n429 )  ;
assign n15327 = state_in[23:16] ;
assign n15328 =  ( n15327 ) == ( bv_8_45_n97 )  ;
assign n15329 = state_in[23:16] ;
assign n15330 =  ( n15329 ) == ( bv_8_44_n5 )  ;
assign n15331 = state_in[23:16] ;
assign n15332 =  ( n15331 ) == ( bv_8_43_n121 )  ;
assign n15333 = state_in[23:16] ;
assign n15334 =  ( n15333 ) == ( bv_8_42_n672 )  ;
assign n15335 = state_in[23:16] ;
assign n15336 =  ( n15335 ) == ( bv_8_41_n29 )  ;
assign n15337 = state_in[23:16] ;
assign n15338 =  ( n15337 ) == ( bv_8_40_n366 )  ;
assign n15339 = state_in[23:16] ;
assign n15340 =  ( n15339 ) == ( bv_8_39_n132 )  ;
assign n15341 = state_in[23:16] ;
assign n15342 =  ( n15341 ) == ( bv_8_38_n444 )  ;
assign n15343 = state_in[23:16] ;
assign n15344 =  ( n15343 ) == ( bv_8_37_n506 )  ;
assign n15345 = state_in[23:16] ;
assign n15346 =  ( n15345 ) == ( bv_8_36_n645 )  ;
assign n15347 = state_in[23:16] ;
assign n15348 =  ( n15347 ) == ( bv_8_35_n696 )  ;
assign n15349 = state_in[23:16] ;
assign n15350 =  ( n15349 ) == ( bv_8_34_n117 )  ;
assign n15351 = state_in[23:16] ;
assign n15352 =  ( n15351 ) == ( bv_8_33_n486 )  ;
assign n15353 = state_in[23:16] ;
assign n15354 =  ( n15353 ) == ( bv_8_32_n463 )  ;
assign n15355 = state_in[23:16] ;
assign n15356 =  ( n15355 ) == ( bv_8_31_n705 )  ;
assign n15357 = state_in[23:16] ;
assign n15358 =  ( n15357 ) == ( bv_8_30_n21 )  ;
assign n15359 = state_in[23:16] ;
assign n15360 =  ( n15359 ) == ( bv_8_29_n625 )  ;
assign n15361 = state_in[23:16] ;
assign n15362 =  ( n15361 ) == ( bv_8_28_n162 )  ;
assign n15363 = state_in[23:16] ;
assign n15364 =  ( n15363 ) == ( bv_8_27_n642 )  ;
assign n15365 = state_in[23:16] ;
assign n15366 =  ( n15365 ) == ( bv_8_26_n53 )  ;
assign n15367 = state_in[23:16] ;
assign n15368 =  ( n15367 ) == ( bv_8_25_n399 )  ;
assign n15369 = state_in[23:16] ;
assign n15370 =  ( n15369 ) == ( bv_8_24_n448 )  ;
assign n15371 = state_in[23:16] ;
assign n15372 =  ( n15371 ) == ( bv_8_23_n144 )  ;
assign n15373 = state_in[23:16] ;
assign n15374 =  ( n15373 ) == ( bv_8_22_n357 )  ;
assign n15375 = state_in[23:16] ;
assign n15376 =  ( n15375 ) == ( bv_8_21_n89 )  ;
assign n15377 = state_in[23:16] ;
assign n15378 =  ( n15377 ) == ( bv_8_20_n341 )  ;
assign n15379 = state_in[23:16] ;
assign n15380 =  ( n15379 ) == ( bv_8_19_n588 )  ;
assign n15381 = state_in[23:16] ;
assign n15382 =  ( n15381 ) == ( bv_8_18_n628 )  ;
assign n15383 = state_in[23:16] ;
assign n15384 =  ( n15383 ) == ( bv_8_17_n525 )  ;
assign n15385 = state_in[23:16] ;
assign n15386 =  ( n15385 ) == ( bv_8_16_n248 )  ;
assign n15387 = state_in[23:16] ;
assign n15388 =  ( n15387 ) == ( bv_8_15_n190 )  ;
assign n15389 = state_in[23:16] ;
assign n15390 =  ( n15389 ) == ( bv_8_14_n648 )  ;
assign n15391 = state_in[23:16] ;
assign n15392 =  ( n15391 ) == ( bv_8_13_n194 )  ;
assign n15393 = state_in[23:16] ;
assign n15394 =  ( n15393 ) == ( bv_8_12_n333 )  ;
assign n15395 = state_in[23:16] ;
assign n15396 =  ( n15395 ) == ( bv_8_11_n379 )  ;
assign n15397 = state_in[23:16] ;
assign n15398 =  ( n15397 ) == ( bv_8_10_n655 )  ;
assign n15399 = state_in[23:16] ;
assign n15400 =  ( n15399 ) == ( bv_8_9_n57 )  ;
assign n15401 = state_in[23:16] ;
assign n15402 =  ( n15401 ) == ( bv_8_8_n669 )  ;
assign n15403 = state_in[23:16] ;
assign n15404 =  ( n15403 ) == ( bv_8_7_n105 )  ;
assign n15405 = state_in[23:16] ;
assign n15406 =  ( n15405 ) == ( bv_8_6_n169 )  ;
assign n15407 = state_in[23:16] ;
assign n15408 =  ( n15407 ) == ( bv_8_5_n492 )  ;
assign n15409 = state_in[23:16] ;
assign n15410 =  ( n15409 ) == ( bv_8_4_n516 )  ;
assign n15411 = state_in[23:16] ;
assign n15412 =  ( n15411 ) == ( bv_8_3_n65 )  ;
assign n15413 = state_in[23:16] ;
assign n15414 =  ( n15413 ) == ( bv_8_2_n751 )  ;
assign n15415 = state_in[23:16] ;
assign n15416 =  ( n15415 ) == ( bv_8_1_n287 )  ;
assign n15417 = state_in[23:16] ;
assign n15418 =  ( n15417 ) == ( bv_8_0_n580 )  ;
assign n15419 =  ( n15418 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n15420 =  ( n15416 ) ? ( bv_8_124_n184 ) : ( n15419 ) ;
assign n15421 =  ( n15414 ) ? ( bv_8_119_n472 ) : ( n15420 ) ;
assign n15422 =  ( n15412 ) ? ( bv_8_123_n17 ) : ( n15421 ) ;
assign n15423 =  ( n15410 ) ? ( bv_8_242_n55 ) : ( n15422 ) ;
assign n15424 =  ( n15408 ) ? ( bv_8_107_n370 ) : ( n15423 ) ;
assign n15425 =  ( n15406 ) ? ( bv_8_111_n244 ) : ( n15424 ) ;
assign n15426 =  ( n15404 ) ? ( bv_8_197_n224 ) : ( n15425 ) ;
assign n15427 =  ( n15402 ) ? ( bv_8_48_n660 ) : ( n15426 ) ;
assign n15428 =  ( n15400 ) ? ( bv_8_1_n287 ) : ( n15427 ) ;
assign n15429 =  ( n15398 ) ? ( bv_8_103_n523 ) : ( n15428 ) ;
assign n15430 =  ( n15396 ) ? ( bv_8_43_n121 ) : ( n15429 ) ;
assign n15431 =  ( n15394 ) ? ( bv_8_254_n7 ) : ( n15430 ) ;
assign n15432 =  ( n15392 ) ? ( bv_8_215_n45 ) : ( n15431 ) ;
assign n15433 =  ( n15390 ) ? ( bv_8_171_n314 ) : ( n15432 ) ;
assign n15434 =  ( n15388 ) ? ( bv_8_118_n480 ) : ( n15433 ) ;
assign n15435 =  ( n15386 ) ? ( bv_8_202_n207 ) : ( n15434 ) ;
assign n15436 =  ( n15384 ) ? ( bv_8_130_n33 ) : ( n15435 ) ;
assign n15437 =  ( n15382 ) ? ( bv_8_201_n85 ) : ( n15436 ) ;
assign n15438 =  ( n15380 ) ? ( bv_8_125_n459 ) : ( n15437 ) ;
assign n15439 =  ( n15378 ) ? ( bv_8_250_n23 ) : ( n15438 ) ;
assign n15440 =  ( n15376 ) ? ( bv_8_89_n61 ) : ( n15439 ) ;
assign n15441 =  ( n15374 ) ? ( bv_8_71_n252 ) : ( n15440 ) ;
assign n15442 =  ( n15372 ) ? ( bv_8_240_n63 ) : ( n15441 ) ;
assign n15443 =  ( n15370 ) ? ( bv_8_173_n307 ) : ( n15442 ) ;
assign n15444 =  ( n15368 ) ? ( bv_8_212_n171 ) : ( n15443 ) ;
assign n15445 =  ( n15366 ) ? ( bv_8_162_n343 ) : ( n15444 ) ;
assign n15446 =  ( n15364 ) ? ( bv_8_175_n302 ) : ( n15445 ) ;
assign n15447 =  ( n15362 ) ? ( bv_8_156_n279 ) : ( n15446 ) ;
assign n15448 =  ( n15360 ) ? ( bv_8_164_n335 ) : ( n15447 ) ;
assign n15449 =  ( n15358 ) ? ( bv_8_114_n494 ) : ( n15448 ) ;
assign n15450 =  ( n15356 ) ? ( bv_8_192_n242 ) : ( n15449 ) ;
assign n15451 =  ( n15354 ) ? ( bv_8_183_n273 ) : ( n15450 ) ;
assign n15452 =  ( n15352 ) ? ( bv_8_253_n11 ) : ( n15451 ) ;
assign n15453 =  ( n15350 ) ? ( bv_8_147_n392 ) : ( n15452 ) ;
assign n15454 =  ( n15348 ) ? ( bv_8_38_n444 ) : ( n15453 ) ;
assign n15455 =  ( n15346 ) ? ( bv_8_54_n616 ) : ( n15454 ) ;
assign n15456 =  ( n15344 ) ? ( bv_8_63_n489 ) : ( n15455 ) ;
assign n15457 =  ( n15342 ) ? ( bv_8_247_n35 ) : ( n15456 ) ;
assign n15458 =  ( n15340 ) ? ( bv_8_204_n177 ) : ( n15457 ) ;
assign n15459 =  ( n15338 ) ? ( bv_8_52_n619 ) : ( n15458 ) ;
assign n15460 =  ( n15336 ) ? ( bv_8_165_n69 ) : ( n15459 ) ;
assign n15461 =  ( n15334 ) ? ( bv_8_229_n107 ) : ( n15460 ) ;
assign n15462 =  ( n15332 ) ? ( bv_8_241_n59 ) : ( n15461 ) ;
assign n15463 =  ( n15330 ) ? ( bv_8_113_n180 ) : ( n15462 ) ;
assign n15464 =  ( n15328 ) ? ( bv_8_216_n157 ) : ( n15463 ) ;
assign n15465 =  ( n15326 ) ? ( bv_8_49_n309 ) : ( n15464 ) ;
assign n15466 =  ( n15324 ) ? ( bv_8_21_n89 ) : ( n15465 ) ;
assign n15467 =  ( n15322 ) ? ( bv_8_4_n516 ) : ( n15466 ) ;
assign n15468 =  ( n15320 ) ? ( bv_8_199_n216 ) : ( n15467 ) ;
assign n15469 =  ( n15318 ) ? ( bv_8_35_n696 ) : ( n15468 ) ;
assign n15470 =  ( n15316 ) ? ( bv_8_195_n232 ) : ( n15469 ) ;
assign n15471 =  ( n15314 ) ? ( bv_8_24_n448 ) : ( n15470 ) ;
assign n15472 =  ( n15312 ) ? ( bv_8_150_n201 ) : ( n15471 ) ;
assign n15473 =  ( n15310 ) ? ( bv_8_5_n492 ) : ( n15472 ) ;
assign n15474 =  ( n15308 ) ? ( bv_8_154_n368 ) : ( n15473 ) ;
assign n15475 =  ( n15306 ) ? ( bv_8_7_n105 ) : ( n15474 ) ;
assign n15476 =  ( n15304 ) ? ( bv_8_18_n628 ) : ( n15475 ) ;
assign n15477 =  ( n15302 ) ? ( bv_8_128_n450 ) : ( n15476 ) ;
assign n15478 =  ( n15300 ) ? ( bv_8_226_n119 ) : ( n15477 ) ;
assign n15479 =  ( n15298 ) ? ( bv_8_235_n83 ) : ( n15478 ) ;
assign n15480 =  ( n15296 ) ? ( bv_8_39_n132 ) : ( n15479 ) ;
assign n15481 =  ( n15294 ) ? ( bv_8_178_n292 ) : ( n15480 ) ;
assign n15482 =  ( n15292 ) ? ( bv_8_117_n484 ) : ( n15481 ) ;
assign n15483 =  ( n15290 ) ? ( bv_8_9_n57 ) : ( n15482 ) ;
assign n15484 =  ( n15288 ) ? ( bv_8_131_n440 ) : ( n15483 ) ;
assign n15485 =  ( n15286 ) ? ( bv_8_44_n5 ) : ( n15484 ) ;
assign n15486 =  ( n15284 ) ? ( bv_8_26_n53 ) : ( n15485 ) ;
assign n15487 =  ( n15282 ) ? ( bv_8_27_n642 ) : ( n15486 ) ;
assign n15488 =  ( n15280 ) ? ( bv_8_110_n294 ) : ( n15487 ) ;
assign n15489 =  ( n15278 ) ? ( bv_8_90_n25 ) : ( n15488 ) ;
assign n15490 =  ( n15276 ) ? ( bv_8_160_n350 ) : ( n15489 ) ;
assign n15491 =  ( n15274 ) ? ( bv_8_82_n578 ) : ( n15490 ) ;
assign n15492 =  ( n15272 ) ? ( bv_8_59_n382 ) : ( n15491 ) ;
assign n15493 =  ( n15270 ) ? ( bv_8_214_n164 ) : ( n15492 ) ;
assign n15494 =  ( n15268 ) ? ( bv_8_179_n289 ) : ( n15493 ) ;
assign n15495 =  ( n15266 ) ? ( bv_8_41_n29 ) : ( n15494 ) ;
assign n15496 =  ( n15264 ) ? ( bv_8_227_n115 ) : ( n15495 ) ;
assign n15497 =  ( n15262 ) ? ( bv_8_47_n652 ) : ( n15496 ) ;
assign n15498 =  ( n15260 ) ? ( bv_8_132_n41 ) : ( n15497 ) ;
assign n15499 =  ( n15258 ) ? ( bv_8_83_n575 ) : ( n15498 ) ;
assign n15500 =  ( n15256 ) ? ( bv_8_209_n182 ) : ( n15499 ) ;
assign n15501 =  ( n15254 ) ? ( bv_8_0_n580 ) : ( n15500 ) ;
assign n15502 =  ( n15252 ) ? ( bv_8_237_n75 ) : ( n15501 ) ;
assign n15503 =  ( n15250 ) ? ( bv_8_32_n463 ) : ( n15502 ) ;
assign n15504 =  ( n15248 ) ? ( bv_8_252_n15 ) : ( n15503 ) ;
assign n15505 =  ( n15246 ) ? ( bv_8_177_n283 ) : ( n15504 ) ;
assign n15506 =  ( n15244 ) ? ( bv_8_91_n555 ) : ( n15505 ) ;
assign n15507 =  ( n15242 ) ? ( bv_8_106_n155 ) : ( n15506 ) ;
assign n15508 =  ( n15240 ) ? ( bv_8_203_n203 ) : ( n15507 ) ;
assign n15509 =  ( n15238 ) ? ( bv_8_190_n250 ) : ( n15508 ) ;
assign n15510 =  ( n15236 ) ? ( bv_8_57_n312 ) : ( n15509 ) ;
assign n15511 =  ( n15234 ) ? ( bv_8_74_n237 ) : ( n15510 ) ;
assign n15512 =  ( n15232 ) ? ( bv_8_76_n596 ) : ( n15511 ) ;
assign n15513 =  ( n15230 ) ? ( bv_8_88_n562 ) : ( n15512 ) ;
assign n15514 =  ( n15228 ) ? ( bv_8_207_n188 ) : ( n15513 ) ;
assign n15515 =  ( n15226 ) ? ( bv_8_208_n37 ) : ( n15514 ) ;
assign n15516 =  ( n15224 ) ? ( bv_8_239_n67 ) : ( n15515 ) ;
assign n15517 =  ( n15222 ) ? ( bv_8_170_n77 ) : ( n15516 ) ;
assign n15518 =  ( n15220 ) ? ( bv_8_251_n19 ) : ( n15517 ) ;
assign n15519 =  ( n15218 ) ? ( bv_8_67_n318 ) : ( n15518 ) ;
assign n15520 =  ( n15216 ) ? ( bv_8_77_n593 ) : ( n15519 ) ;
assign n15521 =  ( n15214 ) ? ( bv_8_51_n101 ) : ( n15520 ) ;
assign n15522 =  ( n15212 ) ? ( bv_8_133_n434 ) : ( n15521 ) ;
assign n15523 =  ( n15210 ) ? ( bv_8_69_n612 ) : ( n15522 ) ;
assign n15524 =  ( n15208 ) ? ( bv_8_249_n27 ) : ( n15523 ) ;
assign n15525 =  ( n15206 ) ? ( bv_8_2_n751 ) : ( n15524 ) ;
assign n15526 =  ( n15204 ) ? ( bv_8_127_n453 ) : ( n15525 ) ;
assign n15527 =  ( n15202 ) ? ( bv_8_80_n73 ) : ( n15526 ) ;
assign n15528 =  ( n15200 ) ? ( bv_8_60_n93 ) : ( n15527 ) ;
assign n15529 =  ( n15198 ) ? ( bv_8_159_n323 ) : ( n15528 ) ;
assign n15530 =  ( n15196 ) ? ( bv_8_168_n13 ) : ( n15529 ) ;
assign n15531 =  ( n15194 ) ? ( bv_8_81_n582 ) : ( n15530 ) ;
assign n15532 =  ( n15192 ) ? ( bv_8_163_n339 ) : ( n15531 ) ;
assign n15533 =  ( n15190 ) ? ( bv_8_64_n573 ) : ( n15532 ) ;
assign n15534 =  ( n15188 ) ? ( bv_8_143_n403 ) : ( n15533 ) ;
assign n15535 =  ( n15186 ) ? ( bv_8_146_n337 ) : ( n15534 ) ;
assign n15536 =  ( n15184 ) ? ( bv_8_157_n359 ) : ( n15535 ) ;
assign n15537 =  ( n15182 ) ? ( bv_8_56_n230 ) : ( n15536 ) ;
assign n15538 =  ( n15180 ) ? ( bv_8_245_n43 ) : ( n15537 ) ;
assign n15539 =  ( n15178 ) ? ( bv_8_188_n257 ) : ( n15538 ) ;
assign n15540 =  ( n15176 ) ? ( bv_8_182_n277 ) : ( n15539 ) ;
assign n15541 =  ( n15174 ) ? ( bv_8_218_n150 ) : ( n15540 ) ;
assign n15542 =  ( n15172 ) ? ( bv_8_33_n486 ) : ( n15541 ) ;
assign n15543 =  ( n15170 ) ? ( bv_8_16_n248 ) : ( n15542 ) ;
assign n15544 =  ( n15168 ) ? ( bv_8_255_n3 ) : ( n15543 ) ;
assign n15545 =  ( n15166 ) ? ( bv_8_243_n51 ) : ( n15544 ) ;
assign n15546 =  ( n15164 ) ? ( bv_8_210_n113 ) : ( n15545 ) ;
assign n15547 =  ( n15162 ) ? ( bv_8_205_n196 ) : ( n15546 ) ;
assign n15548 =  ( n15160 ) ? ( bv_8_12_n333 ) : ( n15547 ) ;
assign n15549 =  ( n15158 ) ? ( bv_8_19_n588 ) : ( n15548 ) ;
assign n15550 =  ( n15156 ) ? ( bv_8_236_n79 ) : ( n15549 ) ;
assign n15551 =  ( n15154 ) ? ( bv_8_95_n545 ) : ( n15550 ) ;
assign n15552 =  ( n15152 ) ? ( bv_8_151_n218 ) : ( n15551 ) ;
assign n15553 =  ( n15150 ) ? ( bv_8_68_n390 ) : ( n15552 ) ;
assign n15554 =  ( n15148 ) ? ( bv_8_23_n144 ) : ( n15553 ) ;
assign n15555 =  ( n15146 ) ? ( bv_8_196_n228 ) : ( n15554 ) ;
assign n15556 =  ( n15144 ) ? ( bv_8_167_n325 ) : ( n15555 ) ;
assign n15557 =  ( n15142 ) ? ( bv_8_126_n456 ) : ( n15556 ) ;
assign n15558 =  ( n15140 ) ? ( bv_8_61_n634 ) : ( n15557 ) ;
assign n15559 =  ( n15138 ) ? ( bv_8_100_n348 ) : ( n15558 ) ;
assign n15560 =  ( n15136 ) ? ( bv_8_93_n498 ) : ( n15559 ) ;
assign n15561 =  ( n15134 ) ? ( bv_8_25_n399 ) : ( n15560 ) ;
assign n15562 =  ( n15132 ) ? ( bv_8_115_n222 ) : ( n15561 ) ;
assign n15563 =  ( n15130 ) ? ( bv_8_96_n542 ) : ( n15562 ) ;
assign n15564 =  ( n15128 ) ? ( bv_8_129_n446 ) : ( n15563 ) ;
assign n15565 =  ( n15126 ) ? ( bv_8_79_n538 ) : ( n15564 ) ;
assign n15566 =  ( n15124 ) ? ( bv_8_220_n142 ) : ( n15565 ) ;
assign n15567 =  ( n15122 ) ? ( bv_8_34_n117 ) : ( n15566 ) ;
assign n15568 =  ( n15120 ) ? ( bv_8_42_n672 ) : ( n15567 ) ;
assign n15569 =  ( n15118 ) ? ( bv_8_144_n173 ) : ( n15568 ) ;
assign n15570 =  ( n15116 ) ? ( bv_8_136_n425 ) : ( n15569 ) ;
assign n15571 =  ( n15114 ) ? ( bv_8_70_n609 ) : ( n15570 ) ;
assign n15572 =  ( n15112 ) ? ( bv_8_238_n71 ) : ( n15571 ) ;
assign n15573 =  ( n15110 ) ? ( bv_8_184_n270 ) : ( n15572 ) ;
assign n15574 =  ( n15108 ) ? ( bv_8_20_n341 ) : ( n15573 ) ;
assign n15575 =  ( n15106 ) ? ( bv_8_222_n134 ) : ( n15574 ) ;
assign n15576 =  ( n15104 ) ? ( bv_8_94_n548 ) : ( n15575 ) ;
assign n15577 =  ( n15102 ) ? ( bv_8_11_n379 ) : ( n15576 ) ;
assign n15578 =  ( n15100 ) ? ( bv_8_219_n146 ) : ( n15577 ) ;
assign n15579 =  ( n15098 ) ? ( bv_8_224_n126 ) : ( n15578 ) ;
assign n15580 =  ( n15096 ) ? ( bv_8_50_n408 ) : ( n15579 ) ;
assign n15581 =  ( n15094 ) ? ( bv_8_58_n136 ) : ( n15580 ) ;
assign n15582 =  ( n15092 ) ? ( bv_8_10_n655 ) : ( n15581 ) ;
assign n15583 =  ( n15090 ) ? ( bv_8_73_n275 ) : ( n15582 ) ;
assign n15584 =  ( n15088 ) ? ( bv_8_6_n169 ) : ( n15583 ) ;
assign n15585 =  ( n15086 ) ? ( bv_8_36_n645 ) : ( n15584 ) ;
assign n15586 =  ( n15084 ) ? ( bv_8_92_n234 ) : ( n15585 ) ;
assign n15587 =  ( n15082 ) ? ( bv_8_194_n159 ) : ( n15586 ) ;
assign n15588 =  ( n15080 ) ? ( bv_8_211_n175 ) : ( n15587 ) ;
assign n15589 =  ( n15078 ) ? ( bv_8_172_n268 ) : ( n15588 ) ;
assign n15590 =  ( n15076 ) ? ( bv_8_98_n536 ) : ( n15589 ) ;
assign n15591 =  ( n15074 ) ? ( bv_8_145_n397 ) : ( n15590 ) ;
assign n15592 =  ( n15072 ) ? ( bv_8_149_n384 ) : ( n15591 ) ;
assign n15593 =  ( n15070 ) ? ( bv_8_228_n111 ) : ( n15592 ) ;
assign n15594 =  ( n15068 ) ? ( bv_8_121_n470 ) : ( n15593 ) ;
assign n15595 =  ( n15066 ) ? ( bv_8_231_n99 ) : ( n15594 ) ;
assign n15596 =  ( n15064 ) ? ( bv_8_200_n213 ) : ( n15595 ) ;
assign n15597 =  ( n15062 ) ? ( bv_8_55_n650 ) : ( n15596 ) ;
assign n15598 =  ( n15060 ) ? ( bv_8_109_n9 ) : ( n15597 ) ;
assign n15599 =  ( n15058 ) ? ( bv_8_141_n410 ) : ( n15598 ) ;
assign n15600 =  ( n15056 ) ? ( bv_8_213_n167 ) : ( n15599 ) ;
assign n15601 =  ( n15054 ) ? ( bv_8_78_n590 ) : ( n15600 ) ;
assign n15602 =  ( n15052 ) ? ( bv_8_169_n109 ) : ( n15601 ) ;
assign n15603 =  ( n15050 ) ? ( bv_8_108_n510 ) : ( n15602 ) ;
assign n15604 =  ( n15048 ) ? ( bv_8_86_n567 ) : ( n15603 ) ;
assign n15605 =  ( n15046 ) ? ( bv_8_244_n47 ) : ( n15604 ) ;
assign n15606 =  ( n15044 ) ? ( bv_8_234_n87 ) : ( n15605 ) ;
assign n15607 =  ( n15042 ) ? ( bv_8_101_n49 ) : ( n15606 ) ;
assign n15608 =  ( n15040 ) ? ( bv_8_122_n416 ) : ( n15607 ) ;
assign n15609 =  ( n15038 ) ? ( bv_8_174_n152 ) : ( n15608 ) ;
assign n15610 =  ( n15036 ) ? ( bv_8_8_n669 ) : ( n15609 ) ;
assign n15611 =  ( n15034 ) ? ( bv_8_186_n263 ) : ( n15610 ) ;
assign n15612 =  ( n15032 ) ? ( bv_8_120_n474 ) : ( n15611 ) ;
assign n15613 =  ( n15030 ) ? ( bv_8_37_n506 ) : ( n15612 ) ;
assign n15614 =  ( n15028 ) ? ( bv_8_46_n429 ) : ( n15613 ) ;
assign n15615 =  ( n15026 ) ? ( bv_8_28_n162 ) : ( n15614 ) ;
assign n15616 =  ( n15024 ) ? ( bv_8_166_n328 ) : ( n15615 ) ;
assign n15617 =  ( n15022 ) ? ( bv_8_180_n285 ) : ( n15616 ) ;
assign n15618 =  ( n15020 ) ? ( bv_8_198_n220 ) : ( n15617 ) ;
assign n15619 =  ( n15018 ) ? ( bv_8_232_n95 ) : ( n15618 ) ;
assign n15620 =  ( n15016 ) ? ( bv_8_221_n138 ) : ( n15619 ) ;
assign n15621 =  ( n15014 ) ? ( bv_8_116_n345 ) : ( n15620 ) ;
assign n15622 =  ( n15012 ) ? ( bv_8_31_n705 ) : ( n15621 ) ;
assign n15623 =  ( n15010 ) ? ( bv_8_75_n503 ) : ( n15622 ) ;
assign n15624 =  ( n15008 ) ? ( bv_8_189_n254 ) : ( n15623 ) ;
assign n15625 =  ( n15006 ) ? ( bv_8_139_n297 ) : ( n15624 ) ;
assign n15626 =  ( n15004 ) ? ( bv_8_138_n418 ) : ( n15625 ) ;
assign n15627 =  ( n15002 ) ? ( bv_8_112_n482 ) : ( n15626 ) ;
assign n15628 =  ( n15000 ) ? ( bv_8_62_n205 ) : ( n15627 ) ;
assign n15629 =  ( n14998 ) ? ( bv_8_181_n281 ) : ( n15628 ) ;
assign n15630 =  ( n14996 ) ? ( bv_8_102_n527 ) : ( n15629 ) ;
assign n15631 =  ( n14994 ) ? ( bv_8_72_n330 ) : ( n15630 ) ;
assign n15632 =  ( n14992 ) ? ( bv_8_3_n65 ) : ( n15631 ) ;
assign n15633 =  ( n14990 ) ? ( bv_8_246_n39 ) : ( n15632 ) ;
assign n15634 =  ( n14988 ) ? ( bv_8_14_n648 ) : ( n15633 ) ;
assign n15635 =  ( n14986 ) ? ( bv_8_97_n198 ) : ( n15634 ) ;
assign n15636 =  ( n14984 ) ? ( bv_8_53_n436 ) : ( n15635 ) ;
assign n15637 =  ( n14982 ) ? ( bv_8_87_n226 ) : ( n15636 ) ;
assign n15638 =  ( n14980 ) ? ( bv_8_185_n266 ) : ( n15637 ) ;
assign n15639 =  ( n14978 ) ? ( bv_8_134_n431 ) : ( n15638 ) ;
assign n15640 =  ( n14976 ) ? ( bv_8_193_n239 ) : ( n15639 ) ;
assign n15641 =  ( n14974 ) ? ( bv_8_29_n625 ) : ( n15640 ) ;
assign n15642 =  ( n14972 ) ? ( bv_8_158_n355 ) : ( n15641 ) ;
assign n15643 =  ( n14970 ) ? ( bv_8_225_n123 ) : ( n15642 ) ;
assign n15644 =  ( n14968 ) ? ( bv_8_248_n31 ) : ( n15643 ) ;
assign n15645 =  ( n14966 ) ? ( bv_8_152_n374 ) : ( n15644 ) ;
assign n15646 =  ( n14964 ) ? ( bv_8_17_n525 ) : ( n15645 ) ;
assign n15647 =  ( n14962 ) ? ( bv_8_105_n148 ) : ( n15646 ) ;
assign n15648 =  ( n14960 ) ? ( bv_8_217_n128 ) : ( n15647 ) ;
assign n15649 =  ( n14958 ) ? ( bv_8_142_n406 ) : ( n15648 ) ;
assign n15650 =  ( n14956 ) ? ( bv_8_148_n388 ) : ( n15649 ) ;
assign n15651 =  ( n14954 ) ? ( bv_8_155_n364 ) : ( n15650 ) ;
assign n15652 =  ( n14952 ) ? ( bv_8_30_n21 ) : ( n15651 ) ;
assign n15653 =  ( n14950 ) ? ( bv_8_135_n81 ) : ( n15652 ) ;
assign n15654 =  ( n14948 ) ? ( bv_8_233_n91 ) : ( n15653 ) ;
assign n15655 =  ( n14946 ) ? ( bv_8_206_n192 ) : ( n15654 ) ;
assign n15656 =  ( n14944 ) ? ( bv_8_85_n423 ) : ( n15655 ) ;
assign n15657 =  ( n14942 ) ? ( bv_8_40_n366 ) : ( n15656 ) ;
assign n15658 =  ( n14940 ) ? ( bv_8_223_n130 ) : ( n15657 ) ;
assign n15659 =  ( n14938 ) ? ( bv_8_140_n376 ) : ( n15658 ) ;
assign n15660 =  ( n14936 ) ? ( bv_8_161_n211 ) : ( n15659 ) ;
assign n15661 =  ( n14934 ) ? ( bv_8_137_n421 ) : ( n15660 ) ;
assign n15662 =  ( n14932 ) ? ( bv_8_13_n194 ) : ( n15661 ) ;
assign n15663 =  ( n14930 ) ? ( bv_8_191_n246 ) : ( n15662 ) ;
assign n15664 =  ( n14928 ) ? ( bv_8_230_n103 ) : ( n15663 ) ;
assign n15665 =  ( n14926 ) ? ( bv_8_66_n466 ) : ( n15664 ) ;
assign n15666 =  ( n14924 ) ? ( bv_8_104_n520 ) : ( n15665 ) ;
assign n15667 =  ( n14922 ) ? ( bv_8_65_n623 ) : ( n15666 ) ;
assign n15668 =  ( n14920 ) ? ( bv_8_153_n140 ) : ( n15667 ) ;
assign n15669 =  ( n14918 ) ? ( bv_8_45_n97 ) : ( n15668 ) ;
assign n15670 =  ( n14916 ) ? ( bv_8_15_n190 ) : ( n15669 ) ;
assign n15671 =  ( n14914 ) ? ( bv_8_176_n299 ) : ( n15670 ) ;
assign n15672 =  ( n14912 ) ? ( bv_8_84_n386 ) : ( n15671 ) ;
assign n15673 =  ( n14910 ) ? ( bv_8_187_n260 ) : ( n15672 ) ;
assign n15674 =  ( n14908 ) ? ( bv_8_22_n357 ) : ( n15673 ) ;
assign n15675 =  ( n14906 ) ^ ( n15674 )  ;
assign n15676 = state_in[23:16] ;
assign n15677 =  ( n15676 ) == ( bv_8_255_n3 )  ;
assign n15678 = state_in[23:16] ;
assign n15679 =  ( n15678 ) == ( bv_8_254_n7 )  ;
assign n15680 = state_in[23:16] ;
assign n15681 =  ( n15680 ) == ( bv_8_253_n11 )  ;
assign n15682 = state_in[23:16] ;
assign n15683 =  ( n15682 ) == ( bv_8_252_n15 )  ;
assign n15684 = state_in[23:16] ;
assign n15685 =  ( n15684 ) == ( bv_8_251_n19 )  ;
assign n15686 = state_in[23:16] ;
assign n15687 =  ( n15686 ) == ( bv_8_250_n23 )  ;
assign n15688 = state_in[23:16] ;
assign n15689 =  ( n15688 ) == ( bv_8_249_n27 )  ;
assign n15690 = state_in[23:16] ;
assign n15691 =  ( n15690 ) == ( bv_8_248_n31 )  ;
assign n15692 = state_in[23:16] ;
assign n15693 =  ( n15692 ) == ( bv_8_247_n35 )  ;
assign n15694 = state_in[23:16] ;
assign n15695 =  ( n15694 ) == ( bv_8_246_n39 )  ;
assign n15696 = state_in[23:16] ;
assign n15697 =  ( n15696 ) == ( bv_8_245_n43 )  ;
assign n15698 = state_in[23:16] ;
assign n15699 =  ( n15698 ) == ( bv_8_244_n47 )  ;
assign n15700 = state_in[23:16] ;
assign n15701 =  ( n15700 ) == ( bv_8_243_n51 )  ;
assign n15702 = state_in[23:16] ;
assign n15703 =  ( n15702 ) == ( bv_8_242_n55 )  ;
assign n15704 = state_in[23:16] ;
assign n15705 =  ( n15704 ) == ( bv_8_241_n59 )  ;
assign n15706 = state_in[23:16] ;
assign n15707 =  ( n15706 ) == ( bv_8_240_n63 )  ;
assign n15708 = state_in[23:16] ;
assign n15709 =  ( n15708 ) == ( bv_8_239_n67 )  ;
assign n15710 = state_in[23:16] ;
assign n15711 =  ( n15710 ) == ( bv_8_238_n71 )  ;
assign n15712 = state_in[23:16] ;
assign n15713 =  ( n15712 ) == ( bv_8_237_n75 )  ;
assign n15714 = state_in[23:16] ;
assign n15715 =  ( n15714 ) == ( bv_8_236_n79 )  ;
assign n15716 = state_in[23:16] ;
assign n15717 =  ( n15716 ) == ( bv_8_235_n83 )  ;
assign n15718 = state_in[23:16] ;
assign n15719 =  ( n15718 ) == ( bv_8_234_n87 )  ;
assign n15720 = state_in[23:16] ;
assign n15721 =  ( n15720 ) == ( bv_8_233_n91 )  ;
assign n15722 = state_in[23:16] ;
assign n15723 =  ( n15722 ) == ( bv_8_232_n95 )  ;
assign n15724 = state_in[23:16] ;
assign n15725 =  ( n15724 ) == ( bv_8_231_n99 )  ;
assign n15726 = state_in[23:16] ;
assign n15727 =  ( n15726 ) == ( bv_8_230_n103 )  ;
assign n15728 = state_in[23:16] ;
assign n15729 =  ( n15728 ) == ( bv_8_229_n107 )  ;
assign n15730 = state_in[23:16] ;
assign n15731 =  ( n15730 ) == ( bv_8_228_n111 )  ;
assign n15732 = state_in[23:16] ;
assign n15733 =  ( n15732 ) == ( bv_8_227_n115 )  ;
assign n15734 = state_in[23:16] ;
assign n15735 =  ( n15734 ) == ( bv_8_226_n119 )  ;
assign n15736 = state_in[23:16] ;
assign n15737 =  ( n15736 ) == ( bv_8_225_n123 )  ;
assign n15738 = state_in[23:16] ;
assign n15739 =  ( n15738 ) == ( bv_8_224_n126 )  ;
assign n15740 = state_in[23:16] ;
assign n15741 =  ( n15740 ) == ( bv_8_223_n130 )  ;
assign n15742 = state_in[23:16] ;
assign n15743 =  ( n15742 ) == ( bv_8_222_n134 )  ;
assign n15744 = state_in[23:16] ;
assign n15745 =  ( n15744 ) == ( bv_8_221_n138 )  ;
assign n15746 = state_in[23:16] ;
assign n15747 =  ( n15746 ) == ( bv_8_220_n142 )  ;
assign n15748 = state_in[23:16] ;
assign n15749 =  ( n15748 ) == ( bv_8_219_n146 )  ;
assign n15750 = state_in[23:16] ;
assign n15751 =  ( n15750 ) == ( bv_8_218_n150 )  ;
assign n15752 = state_in[23:16] ;
assign n15753 =  ( n15752 ) == ( bv_8_217_n128 )  ;
assign n15754 = state_in[23:16] ;
assign n15755 =  ( n15754 ) == ( bv_8_216_n157 )  ;
assign n15756 = state_in[23:16] ;
assign n15757 =  ( n15756 ) == ( bv_8_215_n45 )  ;
assign n15758 = state_in[23:16] ;
assign n15759 =  ( n15758 ) == ( bv_8_214_n164 )  ;
assign n15760 = state_in[23:16] ;
assign n15761 =  ( n15760 ) == ( bv_8_213_n167 )  ;
assign n15762 = state_in[23:16] ;
assign n15763 =  ( n15762 ) == ( bv_8_212_n171 )  ;
assign n15764 = state_in[23:16] ;
assign n15765 =  ( n15764 ) == ( bv_8_211_n175 )  ;
assign n15766 = state_in[23:16] ;
assign n15767 =  ( n15766 ) == ( bv_8_210_n113 )  ;
assign n15768 = state_in[23:16] ;
assign n15769 =  ( n15768 ) == ( bv_8_209_n182 )  ;
assign n15770 = state_in[23:16] ;
assign n15771 =  ( n15770 ) == ( bv_8_208_n37 )  ;
assign n15772 = state_in[23:16] ;
assign n15773 =  ( n15772 ) == ( bv_8_207_n188 )  ;
assign n15774 = state_in[23:16] ;
assign n15775 =  ( n15774 ) == ( bv_8_206_n192 )  ;
assign n15776 = state_in[23:16] ;
assign n15777 =  ( n15776 ) == ( bv_8_205_n196 )  ;
assign n15778 = state_in[23:16] ;
assign n15779 =  ( n15778 ) == ( bv_8_204_n177 )  ;
assign n15780 = state_in[23:16] ;
assign n15781 =  ( n15780 ) == ( bv_8_203_n203 )  ;
assign n15782 = state_in[23:16] ;
assign n15783 =  ( n15782 ) == ( bv_8_202_n207 )  ;
assign n15784 = state_in[23:16] ;
assign n15785 =  ( n15784 ) == ( bv_8_201_n85 )  ;
assign n15786 = state_in[23:16] ;
assign n15787 =  ( n15786 ) == ( bv_8_200_n213 )  ;
assign n15788 = state_in[23:16] ;
assign n15789 =  ( n15788 ) == ( bv_8_199_n216 )  ;
assign n15790 = state_in[23:16] ;
assign n15791 =  ( n15790 ) == ( bv_8_198_n220 )  ;
assign n15792 = state_in[23:16] ;
assign n15793 =  ( n15792 ) == ( bv_8_197_n224 )  ;
assign n15794 = state_in[23:16] ;
assign n15795 =  ( n15794 ) == ( bv_8_196_n228 )  ;
assign n15796 = state_in[23:16] ;
assign n15797 =  ( n15796 ) == ( bv_8_195_n232 )  ;
assign n15798 = state_in[23:16] ;
assign n15799 =  ( n15798 ) == ( bv_8_194_n159 )  ;
assign n15800 = state_in[23:16] ;
assign n15801 =  ( n15800 ) == ( bv_8_193_n239 )  ;
assign n15802 = state_in[23:16] ;
assign n15803 =  ( n15802 ) == ( bv_8_192_n242 )  ;
assign n15804 = state_in[23:16] ;
assign n15805 =  ( n15804 ) == ( bv_8_191_n246 )  ;
assign n15806 = state_in[23:16] ;
assign n15807 =  ( n15806 ) == ( bv_8_190_n250 )  ;
assign n15808 = state_in[23:16] ;
assign n15809 =  ( n15808 ) == ( bv_8_189_n254 )  ;
assign n15810 = state_in[23:16] ;
assign n15811 =  ( n15810 ) == ( bv_8_188_n257 )  ;
assign n15812 = state_in[23:16] ;
assign n15813 =  ( n15812 ) == ( bv_8_187_n260 )  ;
assign n15814 = state_in[23:16] ;
assign n15815 =  ( n15814 ) == ( bv_8_186_n263 )  ;
assign n15816 = state_in[23:16] ;
assign n15817 =  ( n15816 ) == ( bv_8_185_n266 )  ;
assign n15818 = state_in[23:16] ;
assign n15819 =  ( n15818 ) == ( bv_8_184_n270 )  ;
assign n15820 = state_in[23:16] ;
assign n15821 =  ( n15820 ) == ( bv_8_183_n273 )  ;
assign n15822 = state_in[23:16] ;
assign n15823 =  ( n15822 ) == ( bv_8_182_n277 )  ;
assign n15824 = state_in[23:16] ;
assign n15825 =  ( n15824 ) == ( bv_8_181_n281 )  ;
assign n15826 = state_in[23:16] ;
assign n15827 =  ( n15826 ) == ( bv_8_180_n285 )  ;
assign n15828 = state_in[23:16] ;
assign n15829 =  ( n15828 ) == ( bv_8_179_n289 )  ;
assign n15830 = state_in[23:16] ;
assign n15831 =  ( n15830 ) == ( bv_8_178_n292 )  ;
assign n15832 = state_in[23:16] ;
assign n15833 =  ( n15832 ) == ( bv_8_177_n283 )  ;
assign n15834 = state_in[23:16] ;
assign n15835 =  ( n15834 ) == ( bv_8_176_n299 )  ;
assign n15836 = state_in[23:16] ;
assign n15837 =  ( n15836 ) == ( bv_8_175_n302 )  ;
assign n15838 = state_in[23:16] ;
assign n15839 =  ( n15838 ) == ( bv_8_174_n152 )  ;
assign n15840 = state_in[23:16] ;
assign n15841 =  ( n15840 ) == ( bv_8_173_n307 )  ;
assign n15842 = state_in[23:16] ;
assign n15843 =  ( n15842 ) == ( bv_8_172_n268 )  ;
assign n15844 = state_in[23:16] ;
assign n15845 =  ( n15844 ) == ( bv_8_171_n314 )  ;
assign n15846 = state_in[23:16] ;
assign n15847 =  ( n15846 ) == ( bv_8_170_n77 )  ;
assign n15848 = state_in[23:16] ;
assign n15849 =  ( n15848 ) == ( bv_8_169_n109 )  ;
assign n15850 = state_in[23:16] ;
assign n15851 =  ( n15850 ) == ( bv_8_168_n13 )  ;
assign n15852 = state_in[23:16] ;
assign n15853 =  ( n15852 ) == ( bv_8_167_n325 )  ;
assign n15854 = state_in[23:16] ;
assign n15855 =  ( n15854 ) == ( bv_8_166_n328 )  ;
assign n15856 = state_in[23:16] ;
assign n15857 =  ( n15856 ) == ( bv_8_165_n69 )  ;
assign n15858 = state_in[23:16] ;
assign n15859 =  ( n15858 ) == ( bv_8_164_n335 )  ;
assign n15860 = state_in[23:16] ;
assign n15861 =  ( n15860 ) == ( bv_8_163_n339 )  ;
assign n15862 = state_in[23:16] ;
assign n15863 =  ( n15862 ) == ( bv_8_162_n343 )  ;
assign n15864 = state_in[23:16] ;
assign n15865 =  ( n15864 ) == ( bv_8_161_n211 )  ;
assign n15866 = state_in[23:16] ;
assign n15867 =  ( n15866 ) == ( bv_8_160_n350 )  ;
assign n15868 = state_in[23:16] ;
assign n15869 =  ( n15868 ) == ( bv_8_159_n323 )  ;
assign n15870 = state_in[23:16] ;
assign n15871 =  ( n15870 ) == ( bv_8_158_n355 )  ;
assign n15872 = state_in[23:16] ;
assign n15873 =  ( n15872 ) == ( bv_8_157_n359 )  ;
assign n15874 = state_in[23:16] ;
assign n15875 =  ( n15874 ) == ( bv_8_156_n279 )  ;
assign n15876 = state_in[23:16] ;
assign n15877 =  ( n15876 ) == ( bv_8_155_n364 )  ;
assign n15878 = state_in[23:16] ;
assign n15879 =  ( n15878 ) == ( bv_8_154_n368 )  ;
assign n15880 = state_in[23:16] ;
assign n15881 =  ( n15880 ) == ( bv_8_153_n140 )  ;
assign n15882 = state_in[23:16] ;
assign n15883 =  ( n15882 ) == ( bv_8_152_n374 )  ;
assign n15884 = state_in[23:16] ;
assign n15885 =  ( n15884 ) == ( bv_8_151_n218 )  ;
assign n15886 = state_in[23:16] ;
assign n15887 =  ( n15886 ) == ( bv_8_150_n201 )  ;
assign n15888 = state_in[23:16] ;
assign n15889 =  ( n15888 ) == ( bv_8_149_n384 )  ;
assign n15890 = state_in[23:16] ;
assign n15891 =  ( n15890 ) == ( bv_8_148_n388 )  ;
assign n15892 = state_in[23:16] ;
assign n15893 =  ( n15892 ) == ( bv_8_147_n392 )  ;
assign n15894 = state_in[23:16] ;
assign n15895 =  ( n15894 ) == ( bv_8_146_n337 )  ;
assign n15896 = state_in[23:16] ;
assign n15897 =  ( n15896 ) == ( bv_8_145_n397 )  ;
assign n15898 = state_in[23:16] ;
assign n15899 =  ( n15898 ) == ( bv_8_144_n173 )  ;
assign n15900 = state_in[23:16] ;
assign n15901 =  ( n15900 ) == ( bv_8_143_n403 )  ;
assign n15902 = state_in[23:16] ;
assign n15903 =  ( n15902 ) == ( bv_8_142_n406 )  ;
assign n15904 = state_in[23:16] ;
assign n15905 =  ( n15904 ) == ( bv_8_141_n410 )  ;
assign n15906 = state_in[23:16] ;
assign n15907 =  ( n15906 ) == ( bv_8_140_n376 )  ;
assign n15908 = state_in[23:16] ;
assign n15909 =  ( n15908 ) == ( bv_8_139_n297 )  ;
assign n15910 = state_in[23:16] ;
assign n15911 =  ( n15910 ) == ( bv_8_138_n418 )  ;
assign n15912 = state_in[23:16] ;
assign n15913 =  ( n15912 ) == ( bv_8_137_n421 )  ;
assign n15914 = state_in[23:16] ;
assign n15915 =  ( n15914 ) == ( bv_8_136_n425 )  ;
assign n15916 = state_in[23:16] ;
assign n15917 =  ( n15916 ) == ( bv_8_135_n81 )  ;
assign n15918 = state_in[23:16] ;
assign n15919 =  ( n15918 ) == ( bv_8_134_n431 )  ;
assign n15920 = state_in[23:16] ;
assign n15921 =  ( n15920 ) == ( bv_8_133_n434 )  ;
assign n15922 = state_in[23:16] ;
assign n15923 =  ( n15922 ) == ( bv_8_132_n41 )  ;
assign n15924 = state_in[23:16] ;
assign n15925 =  ( n15924 ) == ( bv_8_131_n440 )  ;
assign n15926 = state_in[23:16] ;
assign n15927 =  ( n15926 ) == ( bv_8_130_n33 )  ;
assign n15928 = state_in[23:16] ;
assign n15929 =  ( n15928 ) == ( bv_8_129_n446 )  ;
assign n15930 = state_in[23:16] ;
assign n15931 =  ( n15930 ) == ( bv_8_128_n450 )  ;
assign n15932 = state_in[23:16] ;
assign n15933 =  ( n15932 ) == ( bv_8_127_n453 )  ;
assign n15934 = state_in[23:16] ;
assign n15935 =  ( n15934 ) == ( bv_8_126_n456 )  ;
assign n15936 = state_in[23:16] ;
assign n15937 =  ( n15936 ) == ( bv_8_125_n459 )  ;
assign n15938 = state_in[23:16] ;
assign n15939 =  ( n15938 ) == ( bv_8_124_n184 )  ;
assign n15940 = state_in[23:16] ;
assign n15941 =  ( n15940 ) == ( bv_8_123_n17 )  ;
assign n15942 = state_in[23:16] ;
assign n15943 =  ( n15942 ) == ( bv_8_122_n416 )  ;
assign n15944 = state_in[23:16] ;
assign n15945 =  ( n15944 ) == ( bv_8_121_n470 )  ;
assign n15946 = state_in[23:16] ;
assign n15947 =  ( n15946 ) == ( bv_8_120_n474 )  ;
assign n15948 = state_in[23:16] ;
assign n15949 =  ( n15948 ) == ( bv_8_119_n472 )  ;
assign n15950 = state_in[23:16] ;
assign n15951 =  ( n15950 ) == ( bv_8_118_n480 )  ;
assign n15952 = state_in[23:16] ;
assign n15953 =  ( n15952 ) == ( bv_8_117_n484 )  ;
assign n15954 = state_in[23:16] ;
assign n15955 =  ( n15954 ) == ( bv_8_116_n345 )  ;
assign n15956 = state_in[23:16] ;
assign n15957 =  ( n15956 ) == ( bv_8_115_n222 )  ;
assign n15958 = state_in[23:16] ;
assign n15959 =  ( n15958 ) == ( bv_8_114_n494 )  ;
assign n15960 = state_in[23:16] ;
assign n15961 =  ( n15960 ) == ( bv_8_113_n180 )  ;
assign n15962 = state_in[23:16] ;
assign n15963 =  ( n15962 ) == ( bv_8_112_n482 )  ;
assign n15964 = state_in[23:16] ;
assign n15965 =  ( n15964 ) == ( bv_8_111_n244 )  ;
assign n15966 = state_in[23:16] ;
assign n15967 =  ( n15966 ) == ( bv_8_110_n294 )  ;
assign n15968 = state_in[23:16] ;
assign n15969 =  ( n15968 ) == ( bv_8_109_n9 )  ;
assign n15970 = state_in[23:16] ;
assign n15971 =  ( n15970 ) == ( bv_8_108_n510 )  ;
assign n15972 = state_in[23:16] ;
assign n15973 =  ( n15972 ) == ( bv_8_107_n370 )  ;
assign n15974 = state_in[23:16] ;
assign n15975 =  ( n15974 ) == ( bv_8_106_n155 )  ;
assign n15976 = state_in[23:16] ;
assign n15977 =  ( n15976 ) == ( bv_8_105_n148 )  ;
assign n15978 = state_in[23:16] ;
assign n15979 =  ( n15978 ) == ( bv_8_104_n520 )  ;
assign n15980 = state_in[23:16] ;
assign n15981 =  ( n15980 ) == ( bv_8_103_n523 )  ;
assign n15982 = state_in[23:16] ;
assign n15983 =  ( n15982 ) == ( bv_8_102_n527 )  ;
assign n15984 = state_in[23:16] ;
assign n15985 =  ( n15984 ) == ( bv_8_101_n49 )  ;
assign n15986 = state_in[23:16] ;
assign n15987 =  ( n15986 ) == ( bv_8_100_n348 )  ;
assign n15988 = state_in[23:16] ;
assign n15989 =  ( n15988 ) == ( bv_8_99_n476 )  ;
assign n15990 = state_in[23:16] ;
assign n15991 =  ( n15990 ) == ( bv_8_98_n536 )  ;
assign n15992 = state_in[23:16] ;
assign n15993 =  ( n15992 ) == ( bv_8_97_n198 )  ;
assign n15994 = state_in[23:16] ;
assign n15995 =  ( n15994 ) == ( bv_8_96_n542 )  ;
assign n15996 = state_in[23:16] ;
assign n15997 =  ( n15996 ) == ( bv_8_95_n545 )  ;
assign n15998 = state_in[23:16] ;
assign n15999 =  ( n15998 ) == ( bv_8_94_n548 )  ;
assign n16000 = state_in[23:16] ;
assign n16001 =  ( n16000 ) == ( bv_8_93_n498 )  ;
assign n16002 = state_in[23:16] ;
assign n16003 =  ( n16002 ) == ( bv_8_92_n234 )  ;
assign n16004 = state_in[23:16] ;
assign n16005 =  ( n16004 ) == ( bv_8_91_n555 )  ;
assign n16006 = state_in[23:16] ;
assign n16007 =  ( n16006 ) == ( bv_8_90_n25 )  ;
assign n16008 = state_in[23:16] ;
assign n16009 =  ( n16008 ) == ( bv_8_89_n61 )  ;
assign n16010 = state_in[23:16] ;
assign n16011 =  ( n16010 ) == ( bv_8_88_n562 )  ;
assign n16012 = state_in[23:16] ;
assign n16013 =  ( n16012 ) == ( bv_8_87_n226 )  ;
assign n16014 = state_in[23:16] ;
assign n16015 =  ( n16014 ) == ( bv_8_86_n567 )  ;
assign n16016 = state_in[23:16] ;
assign n16017 =  ( n16016 ) == ( bv_8_85_n423 )  ;
assign n16018 = state_in[23:16] ;
assign n16019 =  ( n16018 ) == ( bv_8_84_n386 )  ;
assign n16020 = state_in[23:16] ;
assign n16021 =  ( n16020 ) == ( bv_8_83_n575 )  ;
assign n16022 = state_in[23:16] ;
assign n16023 =  ( n16022 ) == ( bv_8_82_n578 )  ;
assign n16024 = state_in[23:16] ;
assign n16025 =  ( n16024 ) == ( bv_8_81_n582 )  ;
assign n16026 = state_in[23:16] ;
assign n16027 =  ( n16026 ) == ( bv_8_80_n73 )  ;
assign n16028 = state_in[23:16] ;
assign n16029 =  ( n16028 ) == ( bv_8_79_n538 )  ;
assign n16030 = state_in[23:16] ;
assign n16031 =  ( n16030 ) == ( bv_8_78_n590 )  ;
assign n16032 = state_in[23:16] ;
assign n16033 =  ( n16032 ) == ( bv_8_77_n593 )  ;
assign n16034 = state_in[23:16] ;
assign n16035 =  ( n16034 ) == ( bv_8_76_n596 )  ;
assign n16036 = state_in[23:16] ;
assign n16037 =  ( n16036 ) == ( bv_8_75_n503 )  ;
assign n16038 = state_in[23:16] ;
assign n16039 =  ( n16038 ) == ( bv_8_74_n237 )  ;
assign n16040 = state_in[23:16] ;
assign n16041 =  ( n16040 ) == ( bv_8_73_n275 )  ;
assign n16042 = state_in[23:16] ;
assign n16043 =  ( n16042 ) == ( bv_8_72_n330 )  ;
assign n16044 = state_in[23:16] ;
assign n16045 =  ( n16044 ) == ( bv_8_71_n252 )  ;
assign n16046 = state_in[23:16] ;
assign n16047 =  ( n16046 ) == ( bv_8_70_n609 )  ;
assign n16048 = state_in[23:16] ;
assign n16049 =  ( n16048 ) == ( bv_8_69_n612 )  ;
assign n16050 = state_in[23:16] ;
assign n16051 =  ( n16050 ) == ( bv_8_68_n390 )  ;
assign n16052 = state_in[23:16] ;
assign n16053 =  ( n16052 ) == ( bv_8_67_n318 )  ;
assign n16054 = state_in[23:16] ;
assign n16055 =  ( n16054 ) == ( bv_8_66_n466 )  ;
assign n16056 = state_in[23:16] ;
assign n16057 =  ( n16056 ) == ( bv_8_65_n623 )  ;
assign n16058 = state_in[23:16] ;
assign n16059 =  ( n16058 ) == ( bv_8_64_n573 )  ;
assign n16060 = state_in[23:16] ;
assign n16061 =  ( n16060 ) == ( bv_8_63_n489 )  ;
assign n16062 = state_in[23:16] ;
assign n16063 =  ( n16062 ) == ( bv_8_62_n205 )  ;
assign n16064 = state_in[23:16] ;
assign n16065 =  ( n16064 ) == ( bv_8_61_n634 )  ;
assign n16066 = state_in[23:16] ;
assign n16067 =  ( n16066 ) == ( bv_8_60_n93 )  ;
assign n16068 = state_in[23:16] ;
assign n16069 =  ( n16068 ) == ( bv_8_59_n382 )  ;
assign n16070 = state_in[23:16] ;
assign n16071 =  ( n16070 ) == ( bv_8_58_n136 )  ;
assign n16072 = state_in[23:16] ;
assign n16073 =  ( n16072 ) == ( bv_8_57_n312 )  ;
assign n16074 = state_in[23:16] ;
assign n16075 =  ( n16074 ) == ( bv_8_56_n230 )  ;
assign n16076 = state_in[23:16] ;
assign n16077 =  ( n16076 ) == ( bv_8_55_n650 )  ;
assign n16078 = state_in[23:16] ;
assign n16079 =  ( n16078 ) == ( bv_8_54_n616 )  ;
assign n16080 = state_in[23:16] ;
assign n16081 =  ( n16080 ) == ( bv_8_53_n436 )  ;
assign n16082 = state_in[23:16] ;
assign n16083 =  ( n16082 ) == ( bv_8_52_n619 )  ;
assign n16084 = state_in[23:16] ;
assign n16085 =  ( n16084 ) == ( bv_8_51_n101 )  ;
assign n16086 = state_in[23:16] ;
assign n16087 =  ( n16086 ) == ( bv_8_50_n408 )  ;
assign n16088 = state_in[23:16] ;
assign n16089 =  ( n16088 ) == ( bv_8_49_n309 )  ;
assign n16090 = state_in[23:16] ;
assign n16091 =  ( n16090 ) == ( bv_8_48_n660 )  ;
assign n16092 = state_in[23:16] ;
assign n16093 =  ( n16092 ) == ( bv_8_47_n652 )  ;
assign n16094 = state_in[23:16] ;
assign n16095 =  ( n16094 ) == ( bv_8_46_n429 )  ;
assign n16096 = state_in[23:16] ;
assign n16097 =  ( n16096 ) == ( bv_8_45_n97 )  ;
assign n16098 = state_in[23:16] ;
assign n16099 =  ( n16098 ) == ( bv_8_44_n5 )  ;
assign n16100 = state_in[23:16] ;
assign n16101 =  ( n16100 ) == ( bv_8_43_n121 )  ;
assign n16102 = state_in[23:16] ;
assign n16103 =  ( n16102 ) == ( bv_8_42_n672 )  ;
assign n16104 = state_in[23:16] ;
assign n16105 =  ( n16104 ) == ( bv_8_41_n29 )  ;
assign n16106 = state_in[23:16] ;
assign n16107 =  ( n16106 ) == ( bv_8_40_n366 )  ;
assign n16108 = state_in[23:16] ;
assign n16109 =  ( n16108 ) == ( bv_8_39_n132 )  ;
assign n16110 = state_in[23:16] ;
assign n16111 =  ( n16110 ) == ( bv_8_38_n444 )  ;
assign n16112 = state_in[23:16] ;
assign n16113 =  ( n16112 ) == ( bv_8_37_n506 )  ;
assign n16114 = state_in[23:16] ;
assign n16115 =  ( n16114 ) == ( bv_8_36_n645 )  ;
assign n16116 = state_in[23:16] ;
assign n16117 =  ( n16116 ) == ( bv_8_35_n696 )  ;
assign n16118 = state_in[23:16] ;
assign n16119 =  ( n16118 ) == ( bv_8_34_n117 )  ;
assign n16120 = state_in[23:16] ;
assign n16121 =  ( n16120 ) == ( bv_8_33_n486 )  ;
assign n16122 = state_in[23:16] ;
assign n16123 =  ( n16122 ) == ( bv_8_32_n463 )  ;
assign n16124 = state_in[23:16] ;
assign n16125 =  ( n16124 ) == ( bv_8_31_n705 )  ;
assign n16126 = state_in[23:16] ;
assign n16127 =  ( n16126 ) == ( bv_8_30_n21 )  ;
assign n16128 = state_in[23:16] ;
assign n16129 =  ( n16128 ) == ( bv_8_29_n625 )  ;
assign n16130 = state_in[23:16] ;
assign n16131 =  ( n16130 ) == ( bv_8_28_n162 )  ;
assign n16132 = state_in[23:16] ;
assign n16133 =  ( n16132 ) == ( bv_8_27_n642 )  ;
assign n16134 = state_in[23:16] ;
assign n16135 =  ( n16134 ) == ( bv_8_26_n53 )  ;
assign n16136 = state_in[23:16] ;
assign n16137 =  ( n16136 ) == ( bv_8_25_n399 )  ;
assign n16138 = state_in[23:16] ;
assign n16139 =  ( n16138 ) == ( bv_8_24_n448 )  ;
assign n16140 = state_in[23:16] ;
assign n16141 =  ( n16140 ) == ( bv_8_23_n144 )  ;
assign n16142 = state_in[23:16] ;
assign n16143 =  ( n16142 ) == ( bv_8_22_n357 )  ;
assign n16144 = state_in[23:16] ;
assign n16145 =  ( n16144 ) == ( bv_8_21_n89 )  ;
assign n16146 = state_in[23:16] ;
assign n16147 =  ( n16146 ) == ( bv_8_20_n341 )  ;
assign n16148 = state_in[23:16] ;
assign n16149 =  ( n16148 ) == ( bv_8_19_n588 )  ;
assign n16150 = state_in[23:16] ;
assign n16151 =  ( n16150 ) == ( bv_8_18_n628 )  ;
assign n16152 = state_in[23:16] ;
assign n16153 =  ( n16152 ) == ( bv_8_17_n525 )  ;
assign n16154 = state_in[23:16] ;
assign n16155 =  ( n16154 ) == ( bv_8_16_n248 )  ;
assign n16156 = state_in[23:16] ;
assign n16157 =  ( n16156 ) == ( bv_8_15_n190 )  ;
assign n16158 = state_in[23:16] ;
assign n16159 =  ( n16158 ) == ( bv_8_14_n648 )  ;
assign n16160 = state_in[23:16] ;
assign n16161 =  ( n16160 ) == ( bv_8_13_n194 )  ;
assign n16162 = state_in[23:16] ;
assign n16163 =  ( n16162 ) == ( bv_8_12_n333 )  ;
assign n16164 = state_in[23:16] ;
assign n16165 =  ( n16164 ) == ( bv_8_11_n379 )  ;
assign n16166 = state_in[23:16] ;
assign n16167 =  ( n16166 ) == ( bv_8_10_n655 )  ;
assign n16168 = state_in[23:16] ;
assign n16169 =  ( n16168 ) == ( bv_8_9_n57 )  ;
assign n16170 = state_in[23:16] ;
assign n16171 =  ( n16170 ) == ( bv_8_8_n669 )  ;
assign n16172 = state_in[23:16] ;
assign n16173 =  ( n16172 ) == ( bv_8_7_n105 )  ;
assign n16174 = state_in[23:16] ;
assign n16175 =  ( n16174 ) == ( bv_8_6_n169 )  ;
assign n16176 = state_in[23:16] ;
assign n16177 =  ( n16176 ) == ( bv_8_5_n492 )  ;
assign n16178 = state_in[23:16] ;
assign n16179 =  ( n16178 ) == ( bv_8_4_n516 )  ;
assign n16180 = state_in[23:16] ;
assign n16181 =  ( n16180 ) == ( bv_8_3_n65 )  ;
assign n16182 = state_in[23:16] ;
assign n16183 =  ( n16182 ) == ( bv_8_2_n751 )  ;
assign n16184 = state_in[23:16] ;
assign n16185 =  ( n16184 ) == ( bv_8_1_n287 )  ;
assign n16186 = state_in[23:16] ;
assign n16187 =  ( n16186 ) == ( bv_8_0_n580 )  ;
assign n16188 =  ( n16187 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n16189 =  ( n16185 ) ? ( bv_8_248_n31 ) : ( n16188 ) ;
assign n16190 =  ( n16183 ) ? ( bv_8_238_n71 ) : ( n16189 ) ;
assign n16191 =  ( n16181 ) ? ( bv_8_246_n39 ) : ( n16190 ) ;
assign n16192 =  ( n16179 ) ? ( bv_8_255_n3 ) : ( n16191 ) ;
assign n16193 =  ( n16177 ) ? ( bv_8_214_n164 ) : ( n16192 ) ;
assign n16194 =  ( n16175 ) ? ( bv_8_222_n134 ) : ( n16193 ) ;
assign n16195 =  ( n16173 ) ? ( bv_8_145_n397 ) : ( n16194 ) ;
assign n16196 =  ( n16171 ) ? ( bv_8_96_n542 ) : ( n16195 ) ;
assign n16197 =  ( n16169 ) ? ( bv_8_2_n751 ) : ( n16196 ) ;
assign n16198 =  ( n16167 ) ? ( bv_8_206_n192 ) : ( n16197 ) ;
assign n16199 =  ( n16165 ) ? ( bv_8_86_n567 ) : ( n16198 ) ;
assign n16200 =  ( n16163 ) ? ( bv_8_231_n99 ) : ( n16199 ) ;
assign n16201 =  ( n16161 ) ? ( bv_8_181_n281 ) : ( n16200 ) ;
assign n16202 =  ( n16159 ) ? ( bv_8_77_n593 ) : ( n16201 ) ;
assign n16203 =  ( n16157 ) ? ( bv_8_236_n79 ) : ( n16202 ) ;
assign n16204 =  ( n16155 ) ? ( bv_8_143_n403 ) : ( n16203 ) ;
assign n16205 =  ( n16153 ) ? ( bv_8_31_n705 ) : ( n16204 ) ;
assign n16206 =  ( n16151 ) ? ( bv_8_137_n421 ) : ( n16205 ) ;
assign n16207 =  ( n16149 ) ? ( bv_8_250_n23 ) : ( n16206 ) ;
assign n16208 =  ( n16147 ) ? ( bv_8_239_n67 ) : ( n16207 ) ;
assign n16209 =  ( n16145 ) ? ( bv_8_178_n292 ) : ( n16208 ) ;
assign n16210 =  ( n16143 ) ? ( bv_8_142_n406 ) : ( n16209 ) ;
assign n16211 =  ( n16141 ) ? ( bv_8_251_n19 ) : ( n16210 ) ;
assign n16212 =  ( n16139 ) ? ( bv_8_65_n623 ) : ( n16211 ) ;
assign n16213 =  ( n16137 ) ? ( bv_8_179_n289 ) : ( n16212 ) ;
assign n16214 =  ( n16135 ) ? ( bv_8_95_n545 ) : ( n16213 ) ;
assign n16215 =  ( n16133 ) ? ( bv_8_69_n612 ) : ( n16214 ) ;
assign n16216 =  ( n16131 ) ? ( bv_8_35_n696 ) : ( n16215 ) ;
assign n16217 =  ( n16129 ) ? ( bv_8_83_n575 ) : ( n16216 ) ;
assign n16218 =  ( n16127 ) ? ( bv_8_228_n111 ) : ( n16217 ) ;
assign n16219 =  ( n16125 ) ? ( bv_8_155_n364 ) : ( n16218 ) ;
assign n16220 =  ( n16123 ) ? ( bv_8_117_n484 ) : ( n16219 ) ;
assign n16221 =  ( n16121 ) ? ( bv_8_225_n123 ) : ( n16220 ) ;
assign n16222 =  ( n16119 ) ? ( bv_8_61_n634 ) : ( n16221 ) ;
assign n16223 =  ( n16117 ) ? ( bv_8_76_n596 ) : ( n16222 ) ;
assign n16224 =  ( n16115 ) ? ( bv_8_108_n510 ) : ( n16223 ) ;
assign n16225 =  ( n16113 ) ? ( bv_8_126_n456 ) : ( n16224 ) ;
assign n16226 =  ( n16111 ) ? ( bv_8_245_n43 ) : ( n16225 ) ;
assign n16227 =  ( n16109 ) ? ( bv_8_131_n440 ) : ( n16226 ) ;
assign n16228 =  ( n16107 ) ? ( bv_8_104_n520 ) : ( n16227 ) ;
assign n16229 =  ( n16105 ) ? ( bv_8_81_n582 ) : ( n16228 ) ;
assign n16230 =  ( n16103 ) ? ( bv_8_209_n182 ) : ( n16229 ) ;
assign n16231 =  ( n16101 ) ? ( bv_8_249_n27 ) : ( n16230 ) ;
assign n16232 =  ( n16099 ) ? ( bv_8_226_n119 ) : ( n16231 ) ;
assign n16233 =  ( n16097 ) ? ( bv_8_171_n314 ) : ( n16232 ) ;
assign n16234 =  ( n16095 ) ? ( bv_8_98_n536 ) : ( n16233 ) ;
assign n16235 =  ( n16093 ) ? ( bv_8_42_n672 ) : ( n16234 ) ;
assign n16236 =  ( n16091 ) ? ( bv_8_8_n669 ) : ( n16235 ) ;
assign n16237 =  ( n16089 ) ? ( bv_8_149_n384 ) : ( n16236 ) ;
assign n16238 =  ( n16087 ) ? ( bv_8_70_n609 ) : ( n16237 ) ;
assign n16239 =  ( n16085 ) ? ( bv_8_157_n359 ) : ( n16238 ) ;
assign n16240 =  ( n16083 ) ? ( bv_8_48_n660 ) : ( n16239 ) ;
assign n16241 =  ( n16081 ) ? ( bv_8_55_n650 ) : ( n16240 ) ;
assign n16242 =  ( n16079 ) ? ( bv_8_10_n655 ) : ( n16241 ) ;
assign n16243 =  ( n16077 ) ? ( bv_8_47_n652 ) : ( n16242 ) ;
assign n16244 =  ( n16075 ) ? ( bv_8_14_n648 ) : ( n16243 ) ;
assign n16245 =  ( n16073 ) ? ( bv_8_36_n645 ) : ( n16244 ) ;
assign n16246 =  ( n16071 ) ? ( bv_8_27_n642 ) : ( n16245 ) ;
assign n16247 =  ( n16069 ) ? ( bv_8_223_n130 ) : ( n16246 ) ;
assign n16248 =  ( n16067 ) ? ( bv_8_205_n196 ) : ( n16247 ) ;
assign n16249 =  ( n16065 ) ? ( bv_8_78_n590 ) : ( n16248 ) ;
assign n16250 =  ( n16063 ) ? ( bv_8_127_n453 ) : ( n16249 ) ;
assign n16251 =  ( n16061 ) ? ( bv_8_234_n87 ) : ( n16250 ) ;
assign n16252 =  ( n16059 ) ? ( bv_8_18_n628 ) : ( n16251 ) ;
assign n16253 =  ( n16057 ) ? ( bv_8_29_n625 ) : ( n16252 ) ;
assign n16254 =  ( n16055 ) ? ( bv_8_88_n562 ) : ( n16253 ) ;
assign n16255 =  ( n16053 ) ? ( bv_8_52_n619 ) : ( n16254 ) ;
assign n16256 =  ( n16051 ) ? ( bv_8_54_n616 ) : ( n16255 ) ;
assign n16257 =  ( n16049 ) ? ( bv_8_220_n142 ) : ( n16256 ) ;
assign n16258 =  ( n16047 ) ? ( bv_8_180_n285 ) : ( n16257 ) ;
assign n16259 =  ( n16045 ) ? ( bv_8_91_n555 ) : ( n16258 ) ;
assign n16260 =  ( n16043 ) ? ( bv_8_164_n335 ) : ( n16259 ) ;
assign n16261 =  ( n16041 ) ? ( bv_8_118_n480 ) : ( n16260 ) ;
assign n16262 =  ( n16039 ) ? ( bv_8_183_n273 ) : ( n16261 ) ;
assign n16263 =  ( n16037 ) ? ( bv_8_125_n459 ) : ( n16262 ) ;
assign n16264 =  ( n16035 ) ? ( bv_8_82_n578 ) : ( n16263 ) ;
assign n16265 =  ( n16033 ) ? ( bv_8_221_n138 ) : ( n16264 ) ;
assign n16266 =  ( n16031 ) ? ( bv_8_94_n548 ) : ( n16265 ) ;
assign n16267 =  ( n16029 ) ? ( bv_8_19_n588 ) : ( n16266 ) ;
assign n16268 =  ( n16027 ) ? ( bv_8_166_n328 ) : ( n16267 ) ;
assign n16269 =  ( n16025 ) ? ( bv_8_185_n266 ) : ( n16268 ) ;
assign n16270 =  ( n16023 ) ? ( bv_8_0_n580 ) : ( n16269 ) ;
assign n16271 =  ( n16021 ) ? ( bv_8_193_n239 ) : ( n16270 ) ;
assign n16272 =  ( n16019 ) ? ( bv_8_64_n573 ) : ( n16271 ) ;
assign n16273 =  ( n16017 ) ? ( bv_8_227_n115 ) : ( n16272 ) ;
assign n16274 =  ( n16015 ) ? ( bv_8_121_n470 ) : ( n16273 ) ;
assign n16275 =  ( n16013 ) ? ( bv_8_182_n277 ) : ( n16274 ) ;
assign n16276 =  ( n16011 ) ? ( bv_8_212_n171 ) : ( n16275 ) ;
assign n16277 =  ( n16009 ) ? ( bv_8_141_n410 ) : ( n16276 ) ;
assign n16278 =  ( n16007 ) ? ( bv_8_103_n523 ) : ( n16277 ) ;
assign n16279 =  ( n16005 ) ? ( bv_8_114_n494 ) : ( n16278 ) ;
assign n16280 =  ( n16003 ) ? ( bv_8_148_n388 ) : ( n16279 ) ;
assign n16281 =  ( n16001 ) ? ( bv_8_152_n374 ) : ( n16280 ) ;
assign n16282 =  ( n15999 ) ? ( bv_8_176_n299 ) : ( n16281 ) ;
assign n16283 =  ( n15997 ) ? ( bv_8_133_n434 ) : ( n16282 ) ;
assign n16284 =  ( n15995 ) ? ( bv_8_187_n260 ) : ( n16283 ) ;
assign n16285 =  ( n15993 ) ? ( bv_8_197_n224 ) : ( n16284 ) ;
assign n16286 =  ( n15991 ) ? ( bv_8_79_n538 ) : ( n16285 ) ;
assign n16287 =  ( n15989 ) ? ( bv_8_237_n75 ) : ( n16286 ) ;
assign n16288 =  ( n15987 ) ? ( bv_8_134_n431 ) : ( n16287 ) ;
assign n16289 =  ( n15985 ) ? ( bv_8_154_n368 ) : ( n16288 ) ;
assign n16290 =  ( n15983 ) ? ( bv_8_102_n527 ) : ( n16289 ) ;
assign n16291 =  ( n15981 ) ? ( bv_8_17_n525 ) : ( n16290 ) ;
assign n16292 =  ( n15979 ) ? ( bv_8_138_n418 ) : ( n16291 ) ;
assign n16293 =  ( n15977 ) ? ( bv_8_233_n91 ) : ( n16292 ) ;
assign n16294 =  ( n15975 ) ? ( bv_8_4_n516 ) : ( n16293 ) ;
assign n16295 =  ( n15973 ) ? ( bv_8_254_n7 ) : ( n16294 ) ;
assign n16296 =  ( n15971 ) ? ( bv_8_160_n350 ) : ( n16295 ) ;
assign n16297 =  ( n15969 ) ? ( bv_8_120_n474 ) : ( n16296 ) ;
assign n16298 =  ( n15967 ) ? ( bv_8_37_n506 ) : ( n16297 ) ;
assign n16299 =  ( n15965 ) ? ( bv_8_75_n503 ) : ( n16298 ) ;
assign n16300 =  ( n15963 ) ? ( bv_8_162_n343 ) : ( n16299 ) ;
assign n16301 =  ( n15961 ) ? ( bv_8_93_n498 ) : ( n16300 ) ;
assign n16302 =  ( n15959 ) ? ( bv_8_128_n450 ) : ( n16301 ) ;
assign n16303 =  ( n15957 ) ? ( bv_8_5_n492 ) : ( n16302 ) ;
assign n16304 =  ( n15955 ) ? ( bv_8_63_n489 ) : ( n16303 ) ;
assign n16305 =  ( n15953 ) ? ( bv_8_33_n486 ) : ( n16304 ) ;
assign n16306 =  ( n15951 ) ? ( bv_8_112_n482 ) : ( n16305 ) ;
assign n16307 =  ( n15949 ) ? ( bv_8_241_n59 ) : ( n16306 ) ;
assign n16308 =  ( n15947 ) ? ( bv_8_99_n476 ) : ( n16307 ) ;
assign n16309 =  ( n15945 ) ? ( bv_8_119_n472 ) : ( n16308 ) ;
assign n16310 =  ( n15943 ) ? ( bv_8_175_n302 ) : ( n16309 ) ;
assign n16311 =  ( n15941 ) ? ( bv_8_66_n466 ) : ( n16310 ) ;
assign n16312 =  ( n15939 ) ? ( bv_8_32_n463 ) : ( n16311 ) ;
assign n16313 =  ( n15937 ) ? ( bv_8_229_n107 ) : ( n16312 ) ;
assign n16314 =  ( n15935 ) ? ( bv_8_253_n11 ) : ( n16313 ) ;
assign n16315 =  ( n15933 ) ? ( bv_8_191_n246 ) : ( n16314 ) ;
assign n16316 =  ( n15931 ) ? ( bv_8_129_n446 ) : ( n16315 ) ;
assign n16317 =  ( n15929 ) ? ( bv_8_24_n448 ) : ( n16316 ) ;
assign n16318 =  ( n15927 ) ? ( bv_8_38_n444 ) : ( n16317 ) ;
assign n16319 =  ( n15925 ) ? ( bv_8_195_n232 ) : ( n16318 ) ;
assign n16320 =  ( n15923 ) ? ( bv_8_190_n250 ) : ( n16319 ) ;
assign n16321 =  ( n15921 ) ? ( bv_8_53_n436 ) : ( n16320 ) ;
assign n16322 =  ( n15919 ) ? ( bv_8_136_n425 ) : ( n16321 ) ;
assign n16323 =  ( n15917 ) ? ( bv_8_46_n429 ) : ( n16322 ) ;
assign n16324 =  ( n15915 ) ? ( bv_8_147_n392 ) : ( n16323 ) ;
assign n16325 =  ( n15913 ) ? ( bv_8_85_n423 ) : ( n16324 ) ;
assign n16326 =  ( n15911 ) ? ( bv_8_252_n15 ) : ( n16325 ) ;
assign n16327 =  ( n15909 ) ? ( bv_8_122_n416 ) : ( n16326 ) ;
assign n16328 =  ( n15907 ) ? ( bv_8_200_n213 ) : ( n16327 ) ;
assign n16329 =  ( n15905 ) ? ( bv_8_186_n263 ) : ( n16328 ) ;
assign n16330 =  ( n15903 ) ? ( bv_8_50_n408 ) : ( n16329 ) ;
assign n16331 =  ( n15901 ) ? ( bv_8_230_n103 ) : ( n16330 ) ;
assign n16332 =  ( n15899 ) ? ( bv_8_192_n242 ) : ( n16331 ) ;
assign n16333 =  ( n15897 ) ? ( bv_8_25_n399 ) : ( n16332 ) ;
assign n16334 =  ( n15895 ) ? ( bv_8_158_n355 ) : ( n16333 ) ;
assign n16335 =  ( n15893 ) ? ( bv_8_163_n339 ) : ( n16334 ) ;
assign n16336 =  ( n15891 ) ? ( bv_8_68_n390 ) : ( n16335 ) ;
assign n16337 =  ( n15889 ) ? ( bv_8_84_n386 ) : ( n16336 ) ;
assign n16338 =  ( n15887 ) ? ( bv_8_59_n382 ) : ( n16337 ) ;
assign n16339 =  ( n15885 ) ? ( bv_8_11_n379 ) : ( n16338 ) ;
assign n16340 =  ( n15883 ) ? ( bv_8_140_n376 ) : ( n16339 ) ;
assign n16341 =  ( n15881 ) ? ( bv_8_199_n216 ) : ( n16340 ) ;
assign n16342 =  ( n15879 ) ? ( bv_8_107_n370 ) : ( n16341 ) ;
assign n16343 =  ( n15877 ) ? ( bv_8_40_n366 ) : ( n16342 ) ;
assign n16344 =  ( n15875 ) ? ( bv_8_167_n325 ) : ( n16343 ) ;
assign n16345 =  ( n15873 ) ? ( bv_8_188_n257 ) : ( n16344 ) ;
assign n16346 =  ( n15871 ) ? ( bv_8_22_n357 ) : ( n16345 ) ;
assign n16347 =  ( n15869 ) ? ( bv_8_173_n307 ) : ( n16346 ) ;
assign n16348 =  ( n15867 ) ? ( bv_8_219_n146 ) : ( n16347 ) ;
assign n16349 =  ( n15865 ) ? ( bv_8_100_n348 ) : ( n16348 ) ;
assign n16350 =  ( n15863 ) ? ( bv_8_116_n345 ) : ( n16349 ) ;
assign n16351 =  ( n15861 ) ? ( bv_8_20_n341 ) : ( n16350 ) ;
assign n16352 =  ( n15859 ) ? ( bv_8_146_n337 ) : ( n16351 ) ;
assign n16353 =  ( n15857 ) ? ( bv_8_12_n333 ) : ( n16352 ) ;
assign n16354 =  ( n15855 ) ? ( bv_8_72_n330 ) : ( n16353 ) ;
assign n16355 =  ( n15853 ) ? ( bv_8_184_n270 ) : ( n16354 ) ;
assign n16356 =  ( n15851 ) ? ( bv_8_159_n323 ) : ( n16355 ) ;
assign n16357 =  ( n15849 ) ? ( bv_8_189_n254 ) : ( n16356 ) ;
assign n16358 =  ( n15847 ) ? ( bv_8_67_n318 ) : ( n16357 ) ;
assign n16359 =  ( n15845 ) ? ( bv_8_196_n228 ) : ( n16358 ) ;
assign n16360 =  ( n15843 ) ? ( bv_8_57_n312 ) : ( n16359 ) ;
assign n16361 =  ( n15841 ) ? ( bv_8_49_n309 ) : ( n16360 ) ;
assign n16362 =  ( n15839 ) ? ( bv_8_211_n175 ) : ( n16361 ) ;
assign n16363 =  ( n15837 ) ? ( bv_8_242_n55 ) : ( n16362 ) ;
assign n16364 =  ( n15835 ) ? ( bv_8_213_n167 ) : ( n16363 ) ;
assign n16365 =  ( n15833 ) ? ( bv_8_139_n297 ) : ( n16364 ) ;
assign n16366 =  ( n15831 ) ? ( bv_8_110_n294 ) : ( n16365 ) ;
assign n16367 =  ( n15829 ) ? ( bv_8_218_n150 ) : ( n16366 ) ;
assign n16368 =  ( n15827 ) ? ( bv_8_1_n287 ) : ( n16367 ) ;
assign n16369 =  ( n15825 ) ? ( bv_8_177_n283 ) : ( n16368 ) ;
assign n16370 =  ( n15823 ) ? ( bv_8_156_n279 ) : ( n16369 ) ;
assign n16371 =  ( n15821 ) ? ( bv_8_73_n275 ) : ( n16370 ) ;
assign n16372 =  ( n15819 ) ? ( bv_8_216_n157 ) : ( n16371 ) ;
assign n16373 =  ( n15817 ) ? ( bv_8_172_n268 ) : ( n16372 ) ;
assign n16374 =  ( n15815 ) ? ( bv_8_243_n51 ) : ( n16373 ) ;
assign n16375 =  ( n15813 ) ? ( bv_8_207_n188 ) : ( n16374 ) ;
assign n16376 =  ( n15811 ) ? ( bv_8_202_n207 ) : ( n16375 ) ;
assign n16377 =  ( n15809 ) ? ( bv_8_244_n47 ) : ( n16376 ) ;
assign n16378 =  ( n15807 ) ? ( bv_8_71_n252 ) : ( n16377 ) ;
assign n16379 =  ( n15805 ) ? ( bv_8_16_n248 ) : ( n16378 ) ;
assign n16380 =  ( n15803 ) ? ( bv_8_111_n244 ) : ( n16379 ) ;
assign n16381 =  ( n15801 ) ? ( bv_8_240_n63 ) : ( n16380 ) ;
assign n16382 =  ( n15799 ) ? ( bv_8_74_n237 ) : ( n16381 ) ;
assign n16383 =  ( n15797 ) ? ( bv_8_92_n234 ) : ( n16382 ) ;
assign n16384 =  ( n15795 ) ? ( bv_8_56_n230 ) : ( n16383 ) ;
assign n16385 =  ( n15793 ) ? ( bv_8_87_n226 ) : ( n16384 ) ;
assign n16386 =  ( n15791 ) ? ( bv_8_115_n222 ) : ( n16385 ) ;
assign n16387 =  ( n15789 ) ? ( bv_8_151_n218 ) : ( n16386 ) ;
assign n16388 =  ( n15787 ) ? ( bv_8_203_n203 ) : ( n16387 ) ;
assign n16389 =  ( n15785 ) ? ( bv_8_161_n211 ) : ( n16388 ) ;
assign n16390 =  ( n15783 ) ? ( bv_8_232_n95 ) : ( n16389 ) ;
assign n16391 =  ( n15781 ) ? ( bv_8_62_n205 ) : ( n16390 ) ;
assign n16392 =  ( n15779 ) ? ( bv_8_150_n201 ) : ( n16391 ) ;
assign n16393 =  ( n15777 ) ? ( bv_8_97_n198 ) : ( n16392 ) ;
assign n16394 =  ( n15775 ) ? ( bv_8_13_n194 ) : ( n16393 ) ;
assign n16395 =  ( n15773 ) ? ( bv_8_15_n190 ) : ( n16394 ) ;
assign n16396 =  ( n15771 ) ? ( bv_8_224_n126 ) : ( n16395 ) ;
assign n16397 =  ( n15769 ) ? ( bv_8_124_n184 ) : ( n16396 ) ;
assign n16398 =  ( n15767 ) ? ( bv_8_113_n180 ) : ( n16397 ) ;
assign n16399 =  ( n15765 ) ? ( bv_8_204_n177 ) : ( n16398 ) ;
assign n16400 =  ( n15763 ) ? ( bv_8_144_n173 ) : ( n16399 ) ;
assign n16401 =  ( n15761 ) ? ( bv_8_6_n169 ) : ( n16400 ) ;
assign n16402 =  ( n15759 ) ? ( bv_8_247_n35 ) : ( n16401 ) ;
assign n16403 =  ( n15757 ) ? ( bv_8_28_n162 ) : ( n16402 ) ;
assign n16404 =  ( n15755 ) ? ( bv_8_194_n159 ) : ( n16403 ) ;
assign n16405 =  ( n15753 ) ? ( bv_8_106_n155 ) : ( n16404 ) ;
assign n16406 =  ( n15751 ) ? ( bv_8_174_n152 ) : ( n16405 ) ;
assign n16407 =  ( n15749 ) ? ( bv_8_105_n148 ) : ( n16406 ) ;
assign n16408 =  ( n15747 ) ? ( bv_8_23_n144 ) : ( n16407 ) ;
assign n16409 =  ( n15745 ) ? ( bv_8_153_n140 ) : ( n16408 ) ;
assign n16410 =  ( n15743 ) ? ( bv_8_58_n136 ) : ( n16409 ) ;
assign n16411 =  ( n15741 ) ? ( bv_8_39_n132 ) : ( n16410 ) ;
assign n16412 =  ( n15739 ) ? ( bv_8_217_n128 ) : ( n16411 ) ;
assign n16413 =  ( n15737 ) ? ( bv_8_235_n83 ) : ( n16412 ) ;
assign n16414 =  ( n15735 ) ? ( bv_8_43_n121 ) : ( n16413 ) ;
assign n16415 =  ( n15733 ) ? ( bv_8_34_n117 ) : ( n16414 ) ;
assign n16416 =  ( n15731 ) ? ( bv_8_210_n113 ) : ( n16415 ) ;
assign n16417 =  ( n15729 ) ? ( bv_8_169_n109 ) : ( n16416 ) ;
assign n16418 =  ( n15727 ) ? ( bv_8_7_n105 ) : ( n16417 ) ;
assign n16419 =  ( n15725 ) ? ( bv_8_51_n101 ) : ( n16418 ) ;
assign n16420 =  ( n15723 ) ? ( bv_8_45_n97 ) : ( n16419 ) ;
assign n16421 =  ( n15721 ) ? ( bv_8_60_n93 ) : ( n16420 ) ;
assign n16422 =  ( n15719 ) ? ( bv_8_21_n89 ) : ( n16421 ) ;
assign n16423 =  ( n15717 ) ? ( bv_8_201_n85 ) : ( n16422 ) ;
assign n16424 =  ( n15715 ) ? ( bv_8_135_n81 ) : ( n16423 ) ;
assign n16425 =  ( n15713 ) ? ( bv_8_170_n77 ) : ( n16424 ) ;
assign n16426 =  ( n15711 ) ? ( bv_8_80_n73 ) : ( n16425 ) ;
assign n16427 =  ( n15709 ) ? ( bv_8_165_n69 ) : ( n16426 ) ;
assign n16428 =  ( n15707 ) ? ( bv_8_3_n65 ) : ( n16427 ) ;
assign n16429 =  ( n15705 ) ? ( bv_8_89_n61 ) : ( n16428 ) ;
assign n16430 =  ( n15703 ) ? ( bv_8_9_n57 ) : ( n16429 ) ;
assign n16431 =  ( n15701 ) ? ( bv_8_26_n53 ) : ( n16430 ) ;
assign n16432 =  ( n15699 ) ? ( bv_8_101_n49 ) : ( n16431 ) ;
assign n16433 =  ( n15697 ) ? ( bv_8_215_n45 ) : ( n16432 ) ;
assign n16434 =  ( n15695 ) ? ( bv_8_132_n41 ) : ( n16433 ) ;
assign n16435 =  ( n15693 ) ? ( bv_8_208_n37 ) : ( n16434 ) ;
assign n16436 =  ( n15691 ) ? ( bv_8_130_n33 ) : ( n16435 ) ;
assign n16437 =  ( n15689 ) ? ( bv_8_41_n29 ) : ( n16436 ) ;
assign n16438 =  ( n15687 ) ? ( bv_8_90_n25 ) : ( n16437 ) ;
assign n16439 =  ( n15685 ) ? ( bv_8_30_n21 ) : ( n16438 ) ;
assign n16440 =  ( n15683 ) ? ( bv_8_123_n17 ) : ( n16439 ) ;
assign n16441 =  ( n15681 ) ? ( bv_8_168_n13 ) : ( n16440 ) ;
assign n16442 =  ( n15679 ) ? ( bv_8_109_n9 ) : ( n16441 ) ;
assign n16443 =  ( n15677 ) ? ( bv_8_44_n5 ) : ( n16442 ) ;
assign n16444 =  ( n15675 ) ^ ( n16443 )  ;
assign n16445 = key[63:56] ;
assign n16446 =  ( n16444 ) ^ ( n16445 )  ;
assign n16447 =  { ( n12600 ) , ( n16446 ) }  ;
assign n16448 = state_in[111:104] ;
assign n16449 =  ( n16448 ) == ( bv_8_255_n3 )  ;
assign n16450 = state_in[111:104] ;
assign n16451 =  ( n16450 ) == ( bv_8_254_n7 )  ;
assign n16452 = state_in[111:104] ;
assign n16453 =  ( n16452 ) == ( bv_8_253_n11 )  ;
assign n16454 = state_in[111:104] ;
assign n16455 =  ( n16454 ) == ( bv_8_252_n15 )  ;
assign n16456 = state_in[111:104] ;
assign n16457 =  ( n16456 ) == ( bv_8_251_n19 )  ;
assign n16458 = state_in[111:104] ;
assign n16459 =  ( n16458 ) == ( bv_8_250_n23 )  ;
assign n16460 = state_in[111:104] ;
assign n16461 =  ( n16460 ) == ( bv_8_249_n27 )  ;
assign n16462 = state_in[111:104] ;
assign n16463 =  ( n16462 ) == ( bv_8_248_n31 )  ;
assign n16464 = state_in[111:104] ;
assign n16465 =  ( n16464 ) == ( bv_8_247_n35 )  ;
assign n16466 = state_in[111:104] ;
assign n16467 =  ( n16466 ) == ( bv_8_246_n39 )  ;
assign n16468 = state_in[111:104] ;
assign n16469 =  ( n16468 ) == ( bv_8_245_n43 )  ;
assign n16470 = state_in[111:104] ;
assign n16471 =  ( n16470 ) == ( bv_8_244_n47 )  ;
assign n16472 = state_in[111:104] ;
assign n16473 =  ( n16472 ) == ( bv_8_243_n51 )  ;
assign n16474 = state_in[111:104] ;
assign n16475 =  ( n16474 ) == ( bv_8_242_n55 )  ;
assign n16476 = state_in[111:104] ;
assign n16477 =  ( n16476 ) == ( bv_8_241_n59 )  ;
assign n16478 = state_in[111:104] ;
assign n16479 =  ( n16478 ) == ( bv_8_240_n63 )  ;
assign n16480 = state_in[111:104] ;
assign n16481 =  ( n16480 ) == ( bv_8_239_n67 )  ;
assign n16482 = state_in[111:104] ;
assign n16483 =  ( n16482 ) == ( bv_8_238_n71 )  ;
assign n16484 = state_in[111:104] ;
assign n16485 =  ( n16484 ) == ( bv_8_237_n75 )  ;
assign n16486 = state_in[111:104] ;
assign n16487 =  ( n16486 ) == ( bv_8_236_n79 )  ;
assign n16488 = state_in[111:104] ;
assign n16489 =  ( n16488 ) == ( bv_8_235_n83 )  ;
assign n16490 = state_in[111:104] ;
assign n16491 =  ( n16490 ) == ( bv_8_234_n87 )  ;
assign n16492 = state_in[111:104] ;
assign n16493 =  ( n16492 ) == ( bv_8_233_n91 )  ;
assign n16494 = state_in[111:104] ;
assign n16495 =  ( n16494 ) == ( bv_8_232_n95 )  ;
assign n16496 = state_in[111:104] ;
assign n16497 =  ( n16496 ) == ( bv_8_231_n99 )  ;
assign n16498 = state_in[111:104] ;
assign n16499 =  ( n16498 ) == ( bv_8_230_n103 )  ;
assign n16500 = state_in[111:104] ;
assign n16501 =  ( n16500 ) == ( bv_8_229_n107 )  ;
assign n16502 = state_in[111:104] ;
assign n16503 =  ( n16502 ) == ( bv_8_228_n111 )  ;
assign n16504 = state_in[111:104] ;
assign n16505 =  ( n16504 ) == ( bv_8_227_n115 )  ;
assign n16506 = state_in[111:104] ;
assign n16507 =  ( n16506 ) == ( bv_8_226_n119 )  ;
assign n16508 = state_in[111:104] ;
assign n16509 =  ( n16508 ) == ( bv_8_225_n123 )  ;
assign n16510 = state_in[111:104] ;
assign n16511 =  ( n16510 ) == ( bv_8_224_n126 )  ;
assign n16512 = state_in[111:104] ;
assign n16513 =  ( n16512 ) == ( bv_8_223_n130 )  ;
assign n16514 = state_in[111:104] ;
assign n16515 =  ( n16514 ) == ( bv_8_222_n134 )  ;
assign n16516 = state_in[111:104] ;
assign n16517 =  ( n16516 ) == ( bv_8_221_n138 )  ;
assign n16518 = state_in[111:104] ;
assign n16519 =  ( n16518 ) == ( bv_8_220_n142 )  ;
assign n16520 = state_in[111:104] ;
assign n16521 =  ( n16520 ) == ( bv_8_219_n146 )  ;
assign n16522 = state_in[111:104] ;
assign n16523 =  ( n16522 ) == ( bv_8_218_n150 )  ;
assign n16524 = state_in[111:104] ;
assign n16525 =  ( n16524 ) == ( bv_8_217_n128 )  ;
assign n16526 = state_in[111:104] ;
assign n16527 =  ( n16526 ) == ( bv_8_216_n157 )  ;
assign n16528 = state_in[111:104] ;
assign n16529 =  ( n16528 ) == ( bv_8_215_n45 )  ;
assign n16530 = state_in[111:104] ;
assign n16531 =  ( n16530 ) == ( bv_8_214_n164 )  ;
assign n16532 = state_in[111:104] ;
assign n16533 =  ( n16532 ) == ( bv_8_213_n167 )  ;
assign n16534 = state_in[111:104] ;
assign n16535 =  ( n16534 ) == ( bv_8_212_n171 )  ;
assign n16536 = state_in[111:104] ;
assign n16537 =  ( n16536 ) == ( bv_8_211_n175 )  ;
assign n16538 = state_in[111:104] ;
assign n16539 =  ( n16538 ) == ( bv_8_210_n113 )  ;
assign n16540 = state_in[111:104] ;
assign n16541 =  ( n16540 ) == ( bv_8_209_n182 )  ;
assign n16542 = state_in[111:104] ;
assign n16543 =  ( n16542 ) == ( bv_8_208_n37 )  ;
assign n16544 = state_in[111:104] ;
assign n16545 =  ( n16544 ) == ( bv_8_207_n188 )  ;
assign n16546 = state_in[111:104] ;
assign n16547 =  ( n16546 ) == ( bv_8_206_n192 )  ;
assign n16548 = state_in[111:104] ;
assign n16549 =  ( n16548 ) == ( bv_8_205_n196 )  ;
assign n16550 = state_in[111:104] ;
assign n16551 =  ( n16550 ) == ( bv_8_204_n177 )  ;
assign n16552 = state_in[111:104] ;
assign n16553 =  ( n16552 ) == ( bv_8_203_n203 )  ;
assign n16554 = state_in[111:104] ;
assign n16555 =  ( n16554 ) == ( bv_8_202_n207 )  ;
assign n16556 = state_in[111:104] ;
assign n16557 =  ( n16556 ) == ( bv_8_201_n85 )  ;
assign n16558 = state_in[111:104] ;
assign n16559 =  ( n16558 ) == ( bv_8_200_n213 )  ;
assign n16560 = state_in[111:104] ;
assign n16561 =  ( n16560 ) == ( bv_8_199_n216 )  ;
assign n16562 = state_in[111:104] ;
assign n16563 =  ( n16562 ) == ( bv_8_198_n220 )  ;
assign n16564 = state_in[111:104] ;
assign n16565 =  ( n16564 ) == ( bv_8_197_n224 )  ;
assign n16566 = state_in[111:104] ;
assign n16567 =  ( n16566 ) == ( bv_8_196_n228 )  ;
assign n16568 = state_in[111:104] ;
assign n16569 =  ( n16568 ) == ( bv_8_195_n232 )  ;
assign n16570 = state_in[111:104] ;
assign n16571 =  ( n16570 ) == ( bv_8_194_n159 )  ;
assign n16572 = state_in[111:104] ;
assign n16573 =  ( n16572 ) == ( bv_8_193_n239 )  ;
assign n16574 = state_in[111:104] ;
assign n16575 =  ( n16574 ) == ( bv_8_192_n242 )  ;
assign n16576 = state_in[111:104] ;
assign n16577 =  ( n16576 ) == ( bv_8_191_n246 )  ;
assign n16578 = state_in[111:104] ;
assign n16579 =  ( n16578 ) == ( bv_8_190_n250 )  ;
assign n16580 = state_in[111:104] ;
assign n16581 =  ( n16580 ) == ( bv_8_189_n254 )  ;
assign n16582 = state_in[111:104] ;
assign n16583 =  ( n16582 ) == ( bv_8_188_n257 )  ;
assign n16584 = state_in[111:104] ;
assign n16585 =  ( n16584 ) == ( bv_8_187_n260 )  ;
assign n16586 = state_in[111:104] ;
assign n16587 =  ( n16586 ) == ( bv_8_186_n263 )  ;
assign n16588 = state_in[111:104] ;
assign n16589 =  ( n16588 ) == ( bv_8_185_n266 )  ;
assign n16590 = state_in[111:104] ;
assign n16591 =  ( n16590 ) == ( bv_8_184_n270 )  ;
assign n16592 = state_in[111:104] ;
assign n16593 =  ( n16592 ) == ( bv_8_183_n273 )  ;
assign n16594 = state_in[111:104] ;
assign n16595 =  ( n16594 ) == ( bv_8_182_n277 )  ;
assign n16596 = state_in[111:104] ;
assign n16597 =  ( n16596 ) == ( bv_8_181_n281 )  ;
assign n16598 = state_in[111:104] ;
assign n16599 =  ( n16598 ) == ( bv_8_180_n285 )  ;
assign n16600 = state_in[111:104] ;
assign n16601 =  ( n16600 ) == ( bv_8_179_n289 )  ;
assign n16602 = state_in[111:104] ;
assign n16603 =  ( n16602 ) == ( bv_8_178_n292 )  ;
assign n16604 = state_in[111:104] ;
assign n16605 =  ( n16604 ) == ( bv_8_177_n283 )  ;
assign n16606 = state_in[111:104] ;
assign n16607 =  ( n16606 ) == ( bv_8_176_n299 )  ;
assign n16608 = state_in[111:104] ;
assign n16609 =  ( n16608 ) == ( bv_8_175_n302 )  ;
assign n16610 = state_in[111:104] ;
assign n16611 =  ( n16610 ) == ( bv_8_174_n152 )  ;
assign n16612 = state_in[111:104] ;
assign n16613 =  ( n16612 ) == ( bv_8_173_n307 )  ;
assign n16614 = state_in[111:104] ;
assign n16615 =  ( n16614 ) == ( bv_8_172_n268 )  ;
assign n16616 = state_in[111:104] ;
assign n16617 =  ( n16616 ) == ( bv_8_171_n314 )  ;
assign n16618 = state_in[111:104] ;
assign n16619 =  ( n16618 ) == ( bv_8_170_n77 )  ;
assign n16620 = state_in[111:104] ;
assign n16621 =  ( n16620 ) == ( bv_8_169_n109 )  ;
assign n16622 = state_in[111:104] ;
assign n16623 =  ( n16622 ) == ( bv_8_168_n13 )  ;
assign n16624 = state_in[111:104] ;
assign n16625 =  ( n16624 ) == ( bv_8_167_n325 )  ;
assign n16626 = state_in[111:104] ;
assign n16627 =  ( n16626 ) == ( bv_8_166_n328 )  ;
assign n16628 = state_in[111:104] ;
assign n16629 =  ( n16628 ) == ( bv_8_165_n69 )  ;
assign n16630 = state_in[111:104] ;
assign n16631 =  ( n16630 ) == ( bv_8_164_n335 )  ;
assign n16632 = state_in[111:104] ;
assign n16633 =  ( n16632 ) == ( bv_8_163_n339 )  ;
assign n16634 = state_in[111:104] ;
assign n16635 =  ( n16634 ) == ( bv_8_162_n343 )  ;
assign n16636 = state_in[111:104] ;
assign n16637 =  ( n16636 ) == ( bv_8_161_n211 )  ;
assign n16638 = state_in[111:104] ;
assign n16639 =  ( n16638 ) == ( bv_8_160_n350 )  ;
assign n16640 = state_in[111:104] ;
assign n16641 =  ( n16640 ) == ( bv_8_159_n323 )  ;
assign n16642 = state_in[111:104] ;
assign n16643 =  ( n16642 ) == ( bv_8_158_n355 )  ;
assign n16644 = state_in[111:104] ;
assign n16645 =  ( n16644 ) == ( bv_8_157_n359 )  ;
assign n16646 = state_in[111:104] ;
assign n16647 =  ( n16646 ) == ( bv_8_156_n279 )  ;
assign n16648 = state_in[111:104] ;
assign n16649 =  ( n16648 ) == ( bv_8_155_n364 )  ;
assign n16650 = state_in[111:104] ;
assign n16651 =  ( n16650 ) == ( bv_8_154_n368 )  ;
assign n16652 = state_in[111:104] ;
assign n16653 =  ( n16652 ) == ( bv_8_153_n140 )  ;
assign n16654 = state_in[111:104] ;
assign n16655 =  ( n16654 ) == ( bv_8_152_n374 )  ;
assign n16656 = state_in[111:104] ;
assign n16657 =  ( n16656 ) == ( bv_8_151_n218 )  ;
assign n16658 = state_in[111:104] ;
assign n16659 =  ( n16658 ) == ( bv_8_150_n201 )  ;
assign n16660 = state_in[111:104] ;
assign n16661 =  ( n16660 ) == ( bv_8_149_n384 )  ;
assign n16662 = state_in[111:104] ;
assign n16663 =  ( n16662 ) == ( bv_8_148_n388 )  ;
assign n16664 = state_in[111:104] ;
assign n16665 =  ( n16664 ) == ( bv_8_147_n392 )  ;
assign n16666 = state_in[111:104] ;
assign n16667 =  ( n16666 ) == ( bv_8_146_n337 )  ;
assign n16668 = state_in[111:104] ;
assign n16669 =  ( n16668 ) == ( bv_8_145_n397 )  ;
assign n16670 = state_in[111:104] ;
assign n16671 =  ( n16670 ) == ( bv_8_144_n173 )  ;
assign n16672 = state_in[111:104] ;
assign n16673 =  ( n16672 ) == ( bv_8_143_n403 )  ;
assign n16674 = state_in[111:104] ;
assign n16675 =  ( n16674 ) == ( bv_8_142_n406 )  ;
assign n16676 = state_in[111:104] ;
assign n16677 =  ( n16676 ) == ( bv_8_141_n410 )  ;
assign n16678 = state_in[111:104] ;
assign n16679 =  ( n16678 ) == ( bv_8_140_n376 )  ;
assign n16680 = state_in[111:104] ;
assign n16681 =  ( n16680 ) == ( bv_8_139_n297 )  ;
assign n16682 = state_in[111:104] ;
assign n16683 =  ( n16682 ) == ( bv_8_138_n418 )  ;
assign n16684 = state_in[111:104] ;
assign n16685 =  ( n16684 ) == ( bv_8_137_n421 )  ;
assign n16686 = state_in[111:104] ;
assign n16687 =  ( n16686 ) == ( bv_8_136_n425 )  ;
assign n16688 = state_in[111:104] ;
assign n16689 =  ( n16688 ) == ( bv_8_135_n81 )  ;
assign n16690 = state_in[111:104] ;
assign n16691 =  ( n16690 ) == ( bv_8_134_n431 )  ;
assign n16692 = state_in[111:104] ;
assign n16693 =  ( n16692 ) == ( bv_8_133_n434 )  ;
assign n16694 = state_in[111:104] ;
assign n16695 =  ( n16694 ) == ( bv_8_132_n41 )  ;
assign n16696 = state_in[111:104] ;
assign n16697 =  ( n16696 ) == ( bv_8_131_n440 )  ;
assign n16698 = state_in[111:104] ;
assign n16699 =  ( n16698 ) == ( bv_8_130_n33 )  ;
assign n16700 = state_in[111:104] ;
assign n16701 =  ( n16700 ) == ( bv_8_129_n446 )  ;
assign n16702 = state_in[111:104] ;
assign n16703 =  ( n16702 ) == ( bv_8_128_n450 )  ;
assign n16704 = state_in[111:104] ;
assign n16705 =  ( n16704 ) == ( bv_8_127_n453 )  ;
assign n16706 = state_in[111:104] ;
assign n16707 =  ( n16706 ) == ( bv_8_126_n456 )  ;
assign n16708 = state_in[111:104] ;
assign n16709 =  ( n16708 ) == ( bv_8_125_n459 )  ;
assign n16710 = state_in[111:104] ;
assign n16711 =  ( n16710 ) == ( bv_8_124_n184 )  ;
assign n16712 = state_in[111:104] ;
assign n16713 =  ( n16712 ) == ( bv_8_123_n17 )  ;
assign n16714 = state_in[111:104] ;
assign n16715 =  ( n16714 ) == ( bv_8_122_n416 )  ;
assign n16716 = state_in[111:104] ;
assign n16717 =  ( n16716 ) == ( bv_8_121_n470 )  ;
assign n16718 = state_in[111:104] ;
assign n16719 =  ( n16718 ) == ( bv_8_120_n474 )  ;
assign n16720 = state_in[111:104] ;
assign n16721 =  ( n16720 ) == ( bv_8_119_n472 )  ;
assign n16722 = state_in[111:104] ;
assign n16723 =  ( n16722 ) == ( bv_8_118_n480 )  ;
assign n16724 = state_in[111:104] ;
assign n16725 =  ( n16724 ) == ( bv_8_117_n484 )  ;
assign n16726 = state_in[111:104] ;
assign n16727 =  ( n16726 ) == ( bv_8_116_n345 )  ;
assign n16728 = state_in[111:104] ;
assign n16729 =  ( n16728 ) == ( bv_8_115_n222 )  ;
assign n16730 = state_in[111:104] ;
assign n16731 =  ( n16730 ) == ( bv_8_114_n494 )  ;
assign n16732 = state_in[111:104] ;
assign n16733 =  ( n16732 ) == ( bv_8_113_n180 )  ;
assign n16734 = state_in[111:104] ;
assign n16735 =  ( n16734 ) == ( bv_8_112_n482 )  ;
assign n16736 = state_in[111:104] ;
assign n16737 =  ( n16736 ) == ( bv_8_111_n244 )  ;
assign n16738 = state_in[111:104] ;
assign n16739 =  ( n16738 ) == ( bv_8_110_n294 )  ;
assign n16740 = state_in[111:104] ;
assign n16741 =  ( n16740 ) == ( bv_8_109_n9 )  ;
assign n16742 = state_in[111:104] ;
assign n16743 =  ( n16742 ) == ( bv_8_108_n510 )  ;
assign n16744 = state_in[111:104] ;
assign n16745 =  ( n16744 ) == ( bv_8_107_n370 )  ;
assign n16746 = state_in[111:104] ;
assign n16747 =  ( n16746 ) == ( bv_8_106_n155 )  ;
assign n16748 = state_in[111:104] ;
assign n16749 =  ( n16748 ) == ( bv_8_105_n148 )  ;
assign n16750 = state_in[111:104] ;
assign n16751 =  ( n16750 ) == ( bv_8_104_n520 )  ;
assign n16752 = state_in[111:104] ;
assign n16753 =  ( n16752 ) == ( bv_8_103_n523 )  ;
assign n16754 = state_in[111:104] ;
assign n16755 =  ( n16754 ) == ( bv_8_102_n527 )  ;
assign n16756 = state_in[111:104] ;
assign n16757 =  ( n16756 ) == ( bv_8_101_n49 )  ;
assign n16758 = state_in[111:104] ;
assign n16759 =  ( n16758 ) == ( bv_8_100_n348 )  ;
assign n16760 = state_in[111:104] ;
assign n16761 =  ( n16760 ) == ( bv_8_99_n476 )  ;
assign n16762 = state_in[111:104] ;
assign n16763 =  ( n16762 ) == ( bv_8_98_n536 )  ;
assign n16764 = state_in[111:104] ;
assign n16765 =  ( n16764 ) == ( bv_8_97_n198 )  ;
assign n16766 = state_in[111:104] ;
assign n16767 =  ( n16766 ) == ( bv_8_96_n542 )  ;
assign n16768 = state_in[111:104] ;
assign n16769 =  ( n16768 ) == ( bv_8_95_n545 )  ;
assign n16770 = state_in[111:104] ;
assign n16771 =  ( n16770 ) == ( bv_8_94_n548 )  ;
assign n16772 = state_in[111:104] ;
assign n16773 =  ( n16772 ) == ( bv_8_93_n498 )  ;
assign n16774 = state_in[111:104] ;
assign n16775 =  ( n16774 ) == ( bv_8_92_n234 )  ;
assign n16776 = state_in[111:104] ;
assign n16777 =  ( n16776 ) == ( bv_8_91_n555 )  ;
assign n16778 = state_in[111:104] ;
assign n16779 =  ( n16778 ) == ( bv_8_90_n25 )  ;
assign n16780 = state_in[111:104] ;
assign n16781 =  ( n16780 ) == ( bv_8_89_n61 )  ;
assign n16782 = state_in[111:104] ;
assign n16783 =  ( n16782 ) == ( bv_8_88_n562 )  ;
assign n16784 = state_in[111:104] ;
assign n16785 =  ( n16784 ) == ( bv_8_87_n226 )  ;
assign n16786 = state_in[111:104] ;
assign n16787 =  ( n16786 ) == ( bv_8_86_n567 )  ;
assign n16788 = state_in[111:104] ;
assign n16789 =  ( n16788 ) == ( bv_8_85_n423 )  ;
assign n16790 = state_in[111:104] ;
assign n16791 =  ( n16790 ) == ( bv_8_84_n386 )  ;
assign n16792 = state_in[111:104] ;
assign n16793 =  ( n16792 ) == ( bv_8_83_n575 )  ;
assign n16794 = state_in[111:104] ;
assign n16795 =  ( n16794 ) == ( bv_8_82_n578 )  ;
assign n16796 = state_in[111:104] ;
assign n16797 =  ( n16796 ) == ( bv_8_81_n582 )  ;
assign n16798 = state_in[111:104] ;
assign n16799 =  ( n16798 ) == ( bv_8_80_n73 )  ;
assign n16800 = state_in[111:104] ;
assign n16801 =  ( n16800 ) == ( bv_8_79_n538 )  ;
assign n16802 = state_in[111:104] ;
assign n16803 =  ( n16802 ) == ( bv_8_78_n590 )  ;
assign n16804 = state_in[111:104] ;
assign n16805 =  ( n16804 ) == ( bv_8_77_n593 )  ;
assign n16806 = state_in[111:104] ;
assign n16807 =  ( n16806 ) == ( bv_8_76_n596 )  ;
assign n16808 = state_in[111:104] ;
assign n16809 =  ( n16808 ) == ( bv_8_75_n503 )  ;
assign n16810 = state_in[111:104] ;
assign n16811 =  ( n16810 ) == ( bv_8_74_n237 )  ;
assign n16812 = state_in[111:104] ;
assign n16813 =  ( n16812 ) == ( bv_8_73_n275 )  ;
assign n16814 = state_in[111:104] ;
assign n16815 =  ( n16814 ) == ( bv_8_72_n330 )  ;
assign n16816 = state_in[111:104] ;
assign n16817 =  ( n16816 ) == ( bv_8_71_n252 )  ;
assign n16818 = state_in[111:104] ;
assign n16819 =  ( n16818 ) == ( bv_8_70_n609 )  ;
assign n16820 = state_in[111:104] ;
assign n16821 =  ( n16820 ) == ( bv_8_69_n612 )  ;
assign n16822 = state_in[111:104] ;
assign n16823 =  ( n16822 ) == ( bv_8_68_n390 )  ;
assign n16824 = state_in[111:104] ;
assign n16825 =  ( n16824 ) == ( bv_8_67_n318 )  ;
assign n16826 = state_in[111:104] ;
assign n16827 =  ( n16826 ) == ( bv_8_66_n466 )  ;
assign n16828 = state_in[111:104] ;
assign n16829 =  ( n16828 ) == ( bv_8_65_n623 )  ;
assign n16830 = state_in[111:104] ;
assign n16831 =  ( n16830 ) == ( bv_8_64_n573 )  ;
assign n16832 = state_in[111:104] ;
assign n16833 =  ( n16832 ) == ( bv_8_63_n489 )  ;
assign n16834 = state_in[111:104] ;
assign n16835 =  ( n16834 ) == ( bv_8_62_n205 )  ;
assign n16836 = state_in[111:104] ;
assign n16837 =  ( n16836 ) == ( bv_8_61_n634 )  ;
assign n16838 = state_in[111:104] ;
assign n16839 =  ( n16838 ) == ( bv_8_60_n93 )  ;
assign n16840 = state_in[111:104] ;
assign n16841 =  ( n16840 ) == ( bv_8_59_n382 )  ;
assign n16842 = state_in[111:104] ;
assign n16843 =  ( n16842 ) == ( bv_8_58_n136 )  ;
assign n16844 = state_in[111:104] ;
assign n16845 =  ( n16844 ) == ( bv_8_57_n312 )  ;
assign n16846 = state_in[111:104] ;
assign n16847 =  ( n16846 ) == ( bv_8_56_n230 )  ;
assign n16848 = state_in[111:104] ;
assign n16849 =  ( n16848 ) == ( bv_8_55_n650 )  ;
assign n16850 = state_in[111:104] ;
assign n16851 =  ( n16850 ) == ( bv_8_54_n616 )  ;
assign n16852 = state_in[111:104] ;
assign n16853 =  ( n16852 ) == ( bv_8_53_n436 )  ;
assign n16854 = state_in[111:104] ;
assign n16855 =  ( n16854 ) == ( bv_8_52_n619 )  ;
assign n16856 = state_in[111:104] ;
assign n16857 =  ( n16856 ) == ( bv_8_51_n101 )  ;
assign n16858 = state_in[111:104] ;
assign n16859 =  ( n16858 ) == ( bv_8_50_n408 )  ;
assign n16860 = state_in[111:104] ;
assign n16861 =  ( n16860 ) == ( bv_8_49_n309 )  ;
assign n16862 = state_in[111:104] ;
assign n16863 =  ( n16862 ) == ( bv_8_48_n660 )  ;
assign n16864 = state_in[111:104] ;
assign n16865 =  ( n16864 ) == ( bv_8_47_n652 )  ;
assign n16866 = state_in[111:104] ;
assign n16867 =  ( n16866 ) == ( bv_8_46_n429 )  ;
assign n16868 = state_in[111:104] ;
assign n16869 =  ( n16868 ) == ( bv_8_45_n97 )  ;
assign n16870 = state_in[111:104] ;
assign n16871 =  ( n16870 ) == ( bv_8_44_n5 )  ;
assign n16872 = state_in[111:104] ;
assign n16873 =  ( n16872 ) == ( bv_8_43_n121 )  ;
assign n16874 = state_in[111:104] ;
assign n16875 =  ( n16874 ) == ( bv_8_42_n672 )  ;
assign n16876 = state_in[111:104] ;
assign n16877 =  ( n16876 ) == ( bv_8_41_n29 )  ;
assign n16878 = state_in[111:104] ;
assign n16879 =  ( n16878 ) == ( bv_8_40_n366 )  ;
assign n16880 = state_in[111:104] ;
assign n16881 =  ( n16880 ) == ( bv_8_39_n132 )  ;
assign n16882 = state_in[111:104] ;
assign n16883 =  ( n16882 ) == ( bv_8_38_n444 )  ;
assign n16884 = state_in[111:104] ;
assign n16885 =  ( n16884 ) == ( bv_8_37_n506 )  ;
assign n16886 = state_in[111:104] ;
assign n16887 =  ( n16886 ) == ( bv_8_36_n645 )  ;
assign n16888 = state_in[111:104] ;
assign n16889 =  ( n16888 ) == ( bv_8_35_n696 )  ;
assign n16890 = state_in[111:104] ;
assign n16891 =  ( n16890 ) == ( bv_8_34_n117 )  ;
assign n16892 = state_in[111:104] ;
assign n16893 =  ( n16892 ) == ( bv_8_33_n486 )  ;
assign n16894 = state_in[111:104] ;
assign n16895 =  ( n16894 ) == ( bv_8_32_n463 )  ;
assign n16896 = state_in[111:104] ;
assign n16897 =  ( n16896 ) == ( bv_8_31_n705 )  ;
assign n16898 = state_in[111:104] ;
assign n16899 =  ( n16898 ) == ( bv_8_30_n21 )  ;
assign n16900 = state_in[111:104] ;
assign n16901 =  ( n16900 ) == ( bv_8_29_n625 )  ;
assign n16902 = state_in[111:104] ;
assign n16903 =  ( n16902 ) == ( bv_8_28_n162 )  ;
assign n16904 = state_in[111:104] ;
assign n16905 =  ( n16904 ) == ( bv_8_27_n642 )  ;
assign n16906 = state_in[111:104] ;
assign n16907 =  ( n16906 ) == ( bv_8_26_n53 )  ;
assign n16908 = state_in[111:104] ;
assign n16909 =  ( n16908 ) == ( bv_8_25_n399 )  ;
assign n16910 = state_in[111:104] ;
assign n16911 =  ( n16910 ) == ( bv_8_24_n448 )  ;
assign n16912 = state_in[111:104] ;
assign n16913 =  ( n16912 ) == ( bv_8_23_n144 )  ;
assign n16914 = state_in[111:104] ;
assign n16915 =  ( n16914 ) == ( bv_8_22_n357 )  ;
assign n16916 = state_in[111:104] ;
assign n16917 =  ( n16916 ) == ( bv_8_21_n89 )  ;
assign n16918 = state_in[111:104] ;
assign n16919 =  ( n16918 ) == ( bv_8_20_n341 )  ;
assign n16920 = state_in[111:104] ;
assign n16921 =  ( n16920 ) == ( bv_8_19_n588 )  ;
assign n16922 = state_in[111:104] ;
assign n16923 =  ( n16922 ) == ( bv_8_18_n628 )  ;
assign n16924 = state_in[111:104] ;
assign n16925 =  ( n16924 ) == ( bv_8_17_n525 )  ;
assign n16926 = state_in[111:104] ;
assign n16927 =  ( n16926 ) == ( bv_8_16_n248 )  ;
assign n16928 = state_in[111:104] ;
assign n16929 =  ( n16928 ) == ( bv_8_15_n190 )  ;
assign n16930 = state_in[111:104] ;
assign n16931 =  ( n16930 ) == ( bv_8_14_n648 )  ;
assign n16932 = state_in[111:104] ;
assign n16933 =  ( n16932 ) == ( bv_8_13_n194 )  ;
assign n16934 = state_in[111:104] ;
assign n16935 =  ( n16934 ) == ( bv_8_12_n333 )  ;
assign n16936 = state_in[111:104] ;
assign n16937 =  ( n16936 ) == ( bv_8_11_n379 )  ;
assign n16938 = state_in[111:104] ;
assign n16939 =  ( n16938 ) == ( bv_8_10_n655 )  ;
assign n16940 = state_in[111:104] ;
assign n16941 =  ( n16940 ) == ( bv_8_9_n57 )  ;
assign n16942 = state_in[111:104] ;
assign n16943 =  ( n16942 ) == ( bv_8_8_n669 )  ;
assign n16944 = state_in[111:104] ;
assign n16945 =  ( n16944 ) == ( bv_8_7_n105 )  ;
assign n16946 = state_in[111:104] ;
assign n16947 =  ( n16946 ) == ( bv_8_6_n169 )  ;
assign n16948 = state_in[111:104] ;
assign n16949 =  ( n16948 ) == ( bv_8_5_n492 )  ;
assign n16950 = state_in[111:104] ;
assign n16951 =  ( n16950 ) == ( bv_8_4_n516 )  ;
assign n16952 = state_in[111:104] ;
assign n16953 =  ( n16952 ) == ( bv_8_3_n65 )  ;
assign n16954 = state_in[111:104] ;
assign n16955 =  ( n16954 ) == ( bv_8_2_n751 )  ;
assign n16956 = state_in[111:104] ;
assign n16957 =  ( n16956 ) == ( bv_8_1_n287 )  ;
assign n16958 = state_in[111:104] ;
assign n16959 =  ( n16958 ) == ( bv_8_0_n580 )  ;
assign n16960 =  ( n16959 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n16961 =  ( n16957 ) ? ( bv_8_248_n31 ) : ( n16960 ) ;
assign n16962 =  ( n16955 ) ? ( bv_8_238_n71 ) : ( n16961 ) ;
assign n16963 =  ( n16953 ) ? ( bv_8_246_n39 ) : ( n16962 ) ;
assign n16964 =  ( n16951 ) ? ( bv_8_255_n3 ) : ( n16963 ) ;
assign n16965 =  ( n16949 ) ? ( bv_8_214_n164 ) : ( n16964 ) ;
assign n16966 =  ( n16947 ) ? ( bv_8_222_n134 ) : ( n16965 ) ;
assign n16967 =  ( n16945 ) ? ( bv_8_145_n397 ) : ( n16966 ) ;
assign n16968 =  ( n16943 ) ? ( bv_8_96_n542 ) : ( n16967 ) ;
assign n16969 =  ( n16941 ) ? ( bv_8_2_n751 ) : ( n16968 ) ;
assign n16970 =  ( n16939 ) ? ( bv_8_206_n192 ) : ( n16969 ) ;
assign n16971 =  ( n16937 ) ? ( bv_8_86_n567 ) : ( n16970 ) ;
assign n16972 =  ( n16935 ) ? ( bv_8_231_n99 ) : ( n16971 ) ;
assign n16973 =  ( n16933 ) ? ( bv_8_181_n281 ) : ( n16972 ) ;
assign n16974 =  ( n16931 ) ? ( bv_8_77_n593 ) : ( n16973 ) ;
assign n16975 =  ( n16929 ) ? ( bv_8_236_n79 ) : ( n16974 ) ;
assign n16976 =  ( n16927 ) ? ( bv_8_143_n403 ) : ( n16975 ) ;
assign n16977 =  ( n16925 ) ? ( bv_8_31_n705 ) : ( n16976 ) ;
assign n16978 =  ( n16923 ) ? ( bv_8_137_n421 ) : ( n16977 ) ;
assign n16979 =  ( n16921 ) ? ( bv_8_250_n23 ) : ( n16978 ) ;
assign n16980 =  ( n16919 ) ? ( bv_8_239_n67 ) : ( n16979 ) ;
assign n16981 =  ( n16917 ) ? ( bv_8_178_n292 ) : ( n16980 ) ;
assign n16982 =  ( n16915 ) ? ( bv_8_142_n406 ) : ( n16981 ) ;
assign n16983 =  ( n16913 ) ? ( bv_8_251_n19 ) : ( n16982 ) ;
assign n16984 =  ( n16911 ) ? ( bv_8_65_n623 ) : ( n16983 ) ;
assign n16985 =  ( n16909 ) ? ( bv_8_179_n289 ) : ( n16984 ) ;
assign n16986 =  ( n16907 ) ? ( bv_8_95_n545 ) : ( n16985 ) ;
assign n16987 =  ( n16905 ) ? ( bv_8_69_n612 ) : ( n16986 ) ;
assign n16988 =  ( n16903 ) ? ( bv_8_35_n696 ) : ( n16987 ) ;
assign n16989 =  ( n16901 ) ? ( bv_8_83_n575 ) : ( n16988 ) ;
assign n16990 =  ( n16899 ) ? ( bv_8_228_n111 ) : ( n16989 ) ;
assign n16991 =  ( n16897 ) ? ( bv_8_155_n364 ) : ( n16990 ) ;
assign n16992 =  ( n16895 ) ? ( bv_8_117_n484 ) : ( n16991 ) ;
assign n16993 =  ( n16893 ) ? ( bv_8_225_n123 ) : ( n16992 ) ;
assign n16994 =  ( n16891 ) ? ( bv_8_61_n634 ) : ( n16993 ) ;
assign n16995 =  ( n16889 ) ? ( bv_8_76_n596 ) : ( n16994 ) ;
assign n16996 =  ( n16887 ) ? ( bv_8_108_n510 ) : ( n16995 ) ;
assign n16997 =  ( n16885 ) ? ( bv_8_126_n456 ) : ( n16996 ) ;
assign n16998 =  ( n16883 ) ? ( bv_8_245_n43 ) : ( n16997 ) ;
assign n16999 =  ( n16881 ) ? ( bv_8_131_n440 ) : ( n16998 ) ;
assign n17000 =  ( n16879 ) ? ( bv_8_104_n520 ) : ( n16999 ) ;
assign n17001 =  ( n16877 ) ? ( bv_8_81_n582 ) : ( n17000 ) ;
assign n17002 =  ( n16875 ) ? ( bv_8_209_n182 ) : ( n17001 ) ;
assign n17003 =  ( n16873 ) ? ( bv_8_249_n27 ) : ( n17002 ) ;
assign n17004 =  ( n16871 ) ? ( bv_8_226_n119 ) : ( n17003 ) ;
assign n17005 =  ( n16869 ) ? ( bv_8_171_n314 ) : ( n17004 ) ;
assign n17006 =  ( n16867 ) ? ( bv_8_98_n536 ) : ( n17005 ) ;
assign n17007 =  ( n16865 ) ? ( bv_8_42_n672 ) : ( n17006 ) ;
assign n17008 =  ( n16863 ) ? ( bv_8_8_n669 ) : ( n17007 ) ;
assign n17009 =  ( n16861 ) ? ( bv_8_149_n384 ) : ( n17008 ) ;
assign n17010 =  ( n16859 ) ? ( bv_8_70_n609 ) : ( n17009 ) ;
assign n17011 =  ( n16857 ) ? ( bv_8_157_n359 ) : ( n17010 ) ;
assign n17012 =  ( n16855 ) ? ( bv_8_48_n660 ) : ( n17011 ) ;
assign n17013 =  ( n16853 ) ? ( bv_8_55_n650 ) : ( n17012 ) ;
assign n17014 =  ( n16851 ) ? ( bv_8_10_n655 ) : ( n17013 ) ;
assign n17015 =  ( n16849 ) ? ( bv_8_47_n652 ) : ( n17014 ) ;
assign n17016 =  ( n16847 ) ? ( bv_8_14_n648 ) : ( n17015 ) ;
assign n17017 =  ( n16845 ) ? ( bv_8_36_n645 ) : ( n17016 ) ;
assign n17018 =  ( n16843 ) ? ( bv_8_27_n642 ) : ( n17017 ) ;
assign n17019 =  ( n16841 ) ? ( bv_8_223_n130 ) : ( n17018 ) ;
assign n17020 =  ( n16839 ) ? ( bv_8_205_n196 ) : ( n17019 ) ;
assign n17021 =  ( n16837 ) ? ( bv_8_78_n590 ) : ( n17020 ) ;
assign n17022 =  ( n16835 ) ? ( bv_8_127_n453 ) : ( n17021 ) ;
assign n17023 =  ( n16833 ) ? ( bv_8_234_n87 ) : ( n17022 ) ;
assign n17024 =  ( n16831 ) ? ( bv_8_18_n628 ) : ( n17023 ) ;
assign n17025 =  ( n16829 ) ? ( bv_8_29_n625 ) : ( n17024 ) ;
assign n17026 =  ( n16827 ) ? ( bv_8_88_n562 ) : ( n17025 ) ;
assign n17027 =  ( n16825 ) ? ( bv_8_52_n619 ) : ( n17026 ) ;
assign n17028 =  ( n16823 ) ? ( bv_8_54_n616 ) : ( n17027 ) ;
assign n17029 =  ( n16821 ) ? ( bv_8_220_n142 ) : ( n17028 ) ;
assign n17030 =  ( n16819 ) ? ( bv_8_180_n285 ) : ( n17029 ) ;
assign n17031 =  ( n16817 ) ? ( bv_8_91_n555 ) : ( n17030 ) ;
assign n17032 =  ( n16815 ) ? ( bv_8_164_n335 ) : ( n17031 ) ;
assign n17033 =  ( n16813 ) ? ( bv_8_118_n480 ) : ( n17032 ) ;
assign n17034 =  ( n16811 ) ? ( bv_8_183_n273 ) : ( n17033 ) ;
assign n17035 =  ( n16809 ) ? ( bv_8_125_n459 ) : ( n17034 ) ;
assign n17036 =  ( n16807 ) ? ( bv_8_82_n578 ) : ( n17035 ) ;
assign n17037 =  ( n16805 ) ? ( bv_8_221_n138 ) : ( n17036 ) ;
assign n17038 =  ( n16803 ) ? ( bv_8_94_n548 ) : ( n17037 ) ;
assign n17039 =  ( n16801 ) ? ( bv_8_19_n588 ) : ( n17038 ) ;
assign n17040 =  ( n16799 ) ? ( bv_8_166_n328 ) : ( n17039 ) ;
assign n17041 =  ( n16797 ) ? ( bv_8_185_n266 ) : ( n17040 ) ;
assign n17042 =  ( n16795 ) ? ( bv_8_0_n580 ) : ( n17041 ) ;
assign n17043 =  ( n16793 ) ? ( bv_8_193_n239 ) : ( n17042 ) ;
assign n17044 =  ( n16791 ) ? ( bv_8_64_n573 ) : ( n17043 ) ;
assign n17045 =  ( n16789 ) ? ( bv_8_227_n115 ) : ( n17044 ) ;
assign n17046 =  ( n16787 ) ? ( bv_8_121_n470 ) : ( n17045 ) ;
assign n17047 =  ( n16785 ) ? ( bv_8_182_n277 ) : ( n17046 ) ;
assign n17048 =  ( n16783 ) ? ( bv_8_212_n171 ) : ( n17047 ) ;
assign n17049 =  ( n16781 ) ? ( bv_8_141_n410 ) : ( n17048 ) ;
assign n17050 =  ( n16779 ) ? ( bv_8_103_n523 ) : ( n17049 ) ;
assign n17051 =  ( n16777 ) ? ( bv_8_114_n494 ) : ( n17050 ) ;
assign n17052 =  ( n16775 ) ? ( bv_8_148_n388 ) : ( n17051 ) ;
assign n17053 =  ( n16773 ) ? ( bv_8_152_n374 ) : ( n17052 ) ;
assign n17054 =  ( n16771 ) ? ( bv_8_176_n299 ) : ( n17053 ) ;
assign n17055 =  ( n16769 ) ? ( bv_8_133_n434 ) : ( n17054 ) ;
assign n17056 =  ( n16767 ) ? ( bv_8_187_n260 ) : ( n17055 ) ;
assign n17057 =  ( n16765 ) ? ( bv_8_197_n224 ) : ( n17056 ) ;
assign n17058 =  ( n16763 ) ? ( bv_8_79_n538 ) : ( n17057 ) ;
assign n17059 =  ( n16761 ) ? ( bv_8_237_n75 ) : ( n17058 ) ;
assign n17060 =  ( n16759 ) ? ( bv_8_134_n431 ) : ( n17059 ) ;
assign n17061 =  ( n16757 ) ? ( bv_8_154_n368 ) : ( n17060 ) ;
assign n17062 =  ( n16755 ) ? ( bv_8_102_n527 ) : ( n17061 ) ;
assign n17063 =  ( n16753 ) ? ( bv_8_17_n525 ) : ( n17062 ) ;
assign n17064 =  ( n16751 ) ? ( bv_8_138_n418 ) : ( n17063 ) ;
assign n17065 =  ( n16749 ) ? ( bv_8_233_n91 ) : ( n17064 ) ;
assign n17066 =  ( n16747 ) ? ( bv_8_4_n516 ) : ( n17065 ) ;
assign n17067 =  ( n16745 ) ? ( bv_8_254_n7 ) : ( n17066 ) ;
assign n17068 =  ( n16743 ) ? ( bv_8_160_n350 ) : ( n17067 ) ;
assign n17069 =  ( n16741 ) ? ( bv_8_120_n474 ) : ( n17068 ) ;
assign n17070 =  ( n16739 ) ? ( bv_8_37_n506 ) : ( n17069 ) ;
assign n17071 =  ( n16737 ) ? ( bv_8_75_n503 ) : ( n17070 ) ;
assign n17072 =  ( n16735 ) ? ( bv_8_162_n343 ) : ( n17071 ) ;
assign n17073 =  ( n16733 ) ? ( bv_8_93_n498 ) : ( n17072 ) ;
assign n17074 =  ( n16731 ) ? ( bv_8_128_n450 ) : ( n17073 ) ;
assign n17075 =  ( n16729 ) ? ( bv_8_5_n492 ) : ( n17074 ) ;
assign n17076 =  ( n16727 ) ? ( bv_8_63_n489 ) : ( n17075 ) ;
assign n17077 =  ( n16725 ) ? ( bv_8_33_n486 ) : ( n17076 ) ;
assign n17078 =  ( n16723 ) ? ( bv_8_112_n482 ) : ( n17077 ) ;
assign n17079 =  ( n16721 ) ? ( bv_8_241_n59 ) : ( n17078 ) ;
assign n17080 =  ( n16719 ) ? ( bv_8_99_n476 ) : ( n17079 ) ;
assign n17081 =  ( n16717 ) ? ( bv_8_119_n472 ) : ( n17080 ) ;
assign n17082 =  ( n16715 ) ? ( bv_8_175_n302 ) : ( n17081 ) ;
assign n17083 =  ( n16713 ) ? ( bv_8_66_n466 ) : ( n17082 ) ;
assign n17084 =  ( n16711 ) ? ( bv_8_32_n463 ) : ( n17083 ) ;
assign n17085 =  ( n16709 ) ? ( bv_8_229_n107 ) : ( n17084 ) ;
assign n17086 =  ( n16707 ) ? ( bv_8_253_n11 ) : ( n17085 ) ;
assign n17087 =  ( n16705 ) ? ( bv_8_191_n246 ) : ( n17086 ) ;
assign n17088 =  ( n16703 ) ? ( bv_8_129_n446 ) : ( n17087 ) ;
assign n17089 =  ( n16701 ) ? ( bv_8_24_n448 ) : ( n17088 ) ;
assign n17090 =  ( n16699 ) ? ( bv_8_38_n444 ) : ( n17089 ) ;
assign n17091 =  ( n16697 ) ? ( bv_8_195_n232 ) : ( n17090 ) ;
assign n17092 =  ( n16695 ) ? ( bv_8_190_n250 ) : ( n17091 ) ;
assign n17093 =  ( n16693 ) ? ( bv_8_53_n436 ) : ( n17092 ) ;
assign n17094 =  ( n16691 ) ? ( bv_8_136_n425 ) : ( n17093 ) ;
assign n17095 =  ( n16689 ) ? ( bv_8_46_n429 ) : ( n17094 ) ;
assign n17096 =  ( n16687 ) ? ( bv_8_147_n392 ) : ( n17095 ) ;
assign n17097 =  ( n16685 ) ? ( bv_8_85_n423 ) : ( n17096 ) ;
assign n17098 =  ( n16683 ) ? ( bv_8_252_n15 ) : ( n17097 ) ;
assign n17099 =  ( n16681 ) ? ( bv_8_122_n416 ) : ( n17098 ) ;
assign n17100 =  ( n16679 ) ? ( bv_8_200_n213 ) : ( n17099 ) ;
assign n17101 =  ( n16677 ) ? ( bv_8_186_n263 ) : ( n17100 ) ;
assign n17102 =  ( n16675 ) ? ( bv_8_50_n408 ) : ( n17101 ) ;
assign n17103 =  ( n16673 ) ? ( bv_8_230_n103 ) : ( n17102 ) ;
assign n17104 =  ( n16671 ) ? ( bv_8_192_n242 ) : ( n17103 ) ;
assign n17105 =  ( n16669 ) ? ( bv_8_25_n399 ) : ( n17104 ) ;
assign n17106 =  ( n16667 ) ? ( bv_8_158_n355 ) : ( n17105 ) ;
assign n17107 =  ( n16665 ) ? ( bv_8_163_n339 ) : ( n17106 ) ;
assign n17108 =  ( n16663 ) ? ( bv_8_68_n390 ) : ( n17107 ) ;
assign n17109 =  ( n16661 ) ? ( bv_8_84_n386 ) : ( n17108 ) ;
assign n17110 =  ( n16659 ) ? ( bv_8_59_n382 ) : ( n17109 ) ;
assign n17111 =  ( n16657 ) ? ( bv_8_11_n379 ) : ( n17110 ) ;
assign n17112 =  ( n16655 ) ? ( bv_8_140_n376 ) : ( n17111 ) ;
assign n17113 =  ( n16653 ) ? ( bv_8_199_n216 ) : ( n17112 ) ;
assign n17114 =  ( n16651 ) ? ( bv_8_107_n370 ) : ( n17113 ) ;
assign n17115 =  ( n16649 ) ? ( bv_8_40_n366 ) : ( n17114 ) ;
assign n17116 =  ( n16647 ) ? ( bv_8_167_n325 ) : ( n17115 ) ;
assign n17117 =  ( n16645 ) ? ( bv_8_188_n257 ) : ( n17116 ) ;
assign n17118 =  ( n16643 ) ? ( bv_8_22_n357 ) : ( n17117 ) ;
assign n17119 =  ( n16641 ) ? ( bv_8_173_n307 ) : ( n17118 ) ;
assign n17120 =  ( n16639 ) ? ( bv_8_219_n146 ) : ( n17119 ) ;
assign n17121 =  ( n16637 ) ? ( bv_8_100_n348 ) : ( n17120 ) ;
assign n17122 =  ( n16635 ) ? ( bv_8_116_n345 ) : ( n17121 ) ;
assign n17123 =  ( n16633 ) ? ( bv_8_20_n341 ) : ( n17122 ) ;
assign n17124 =  ( n16631 ) ? ( bv_8_146_n337 ) : ( n17123 ) ;
assign n17125 =  ( n16629 ) ? ( bv_8_12_n333 ) : ( n17124 ) ;
assign n17126 =  ( n16627 ) ? ( bv_8_72_n330 ) : ( n17125 ) ;
assign n17127 =  ( n16625 ) ? ( bv_8_184_n270 ) : ( n17126 ) ;
assign n17128 =  ( n16623 ) ? ( bv_8_159_n323 ) : ( n17127 ) ;
assign n17129 =  ( n16621 ) ? ( bv_8_189_n254 ) : ( n17128 ) ;
assign n17130 =  ( n16619 ) ? ( bv_8_67_n318 ) : ( n17129 ) ;
assign n17131 =  ( n16617 ) ? ( bv_8_196_n228 ) : ( n17130 ) ;
assign n17132 =  ( n16615 ) ? ( bv_8_57_n312 ) : ( n17131 ) ;
assign n17133 =  ( n16613 ) ? ( bv_8_49_n309 ) : ( n17132 ) ;
assign n17134 =  ( n16611 ) ? ( bv_8_211_n175 ) : ( n17133 ) ;
assign n17135 =  ( n16609 ) ? ( bv_8_242_n55 ) : ( n17134 ) ;
assign n17136 =  ( n16607 ) ? ( bv_8_213_n167 ) : ( n17135 ) ;
assign n17137 =  ( n16605 ) ? ( bv_8_139_n297 ) : ( n17136 ) ;
assign n17138 =  ( n16603 ) ? ( bv_8_110_n294 ) : ( n17137 ) ;
assign n17139 =  ( n16601 ) ? ( bv_8_218_n150 ) : ( n17138 ) ;
assign n17140 =  ( n16599 ) ? ( bv_8_1_n287 ) : ( n17139 ) ;
assign n17141 =  ( n16597 ) ? ( bv_8_177_n283 ) : ( n17140 ) ;
assign n17142 =  ( n16595 ) ? ( bv_8_156_n279 ) : ( n17141 ) ;
assign n17143 =  ( n16593 ) ? ( bv_8_73_n275 ) : ( n17142 ) ;
assign n17144 =  ( n16591 ) ? ( bv_8_216_n157 ) : ( n17143 ) ;
assign n17145 =  ( n16589 ) ? ( bv_8_172_n268 ) : ( n17144 ) ;
assign n17146 =  ( n16587 ) ? ( bv_8_243_n51 ) : ( n17145 ) ;
assign n17147 =  ( n16585 ) ? ( bv_8_207_n188 ) : ( n17146 ) ;
assign n17148 =  ( n16583 ) ? ( bv_8_202_n207 ) : ( n17147 ) ;
assign n17149 =  ( n16581 ) ? ( bv_8_244_n47 ) : ( n17148 ) ;
assign n17150 =  ( n16579 ) ? ( bv_8_71_n252 ) : ( n17149 ) ;
assign n17151 =  ( n16577 ) ? ( bv_8_16_n248 ) : ( n17150 ) ;
assign n17152 =  ( n16575 ) ? ( bv_8_111_n244 ) : ( n17151 ) ;
assign n17153 =  ( n16573 ) ? ( bv_8_240_n63 ) : ( n17152 ) ;
assign n17154 =  ( n16571 ) ? ( bv_8_74_n237 ) : ( n17153 ) ;
assign n17155 =  ( n16569 ) ? ( bv_8_92_n234 ) : ( n17154 ) ;
assign n17156 =  ( n16567 ) ? ( bv_8_56_n230 ) : ( n17155 ) ;
assign n17157 =  ( n16565 ) ? ( bv_8_87_n226 ) : ( n17156 ) ;
assign n17158 =  ( n16563 ) ? ( bv_8_115_n222 ) : ( n17157 ) ;
assign n17159 =  ( n16561 ) ? ( bv_8_151_n218 ) : ( n17158 ) ;
assign n17160 =  ( n16559 ) ? ( bv_8_203_n203 ) : ( n17159 ) ;
assign n17161 =  ( n16557 ) ? ( bv_8_161_n211 ) : ( n17160 ) ;
assign n17162 =  ( n16555 ) ? ( bv_8_232_n95 ) : ( n17161 ) ;
assign n17163 =  ( n16553 ) ? ( bv_8_62_n205 ) : ( n17162 ) ;
assign n17164 =  ( n16551 ) ? ( bv_8_150_n201 ) : ( n17163 ) ;
assign n17165 =  ( n16549 ) ? ( bv_8_97_n198 ) : ( n17164 ) ;
assign n17166 =  ( n16547 ) ? ( bv_8_13_n194 ) : ( n17165 ) ;
assign n17167 =  ( n16545 ) ? ( bv_8_15_n190 ) : ( n17166 ) ;
assign n17168 =  ( n16543 ) ? ( bv_8_224_n126 ) : ( n17167 ) ;
assign n17169 =  ( n16541 ) ? ( bv_8_124_n184 ) : ( n17168 ) ;
assign n17170 =  ( n16539 ) ? ( bv_8_113_n180 ) : ( n17169 ) ;
assign n17171 =  ( n16537 ) ? ( bv_8_204_n177 ) : ( n17170 ) ;
assign n17172 =  ( n16535 ) ? ( bv_8_144_n173 ) : ( n17171 ) ;
assign n17173 =  ( n16533 ) ? ( bv_8_6_n169 ) : ( n17172 ) ;
assign n17174 =  ( n16531 ) ? ( bv_8_247_n35 ) : ( n17173 ) ;
assign n17175 =  ( n16529 ) ? ( bv_8_28_n162 ) : ( n17174 ) ;
assign n17176 =  ( n16527 ) ? ( bv_8_194_n159 ) : ( n17175 ) ;
assign n17177 =  ( n16525 ) ? ( bv_8_106_n155 ) : ( n17176 ) ;
assign n17178 =  ( n16523 ) ? ( bv_8_174_n152 ) : ( n17177 ) ;
assign n17179 =  ( n16521 ) ? ( bv_8_105_n148 ) : ( n17178 ) ;
assign n17180 =  ( n16519 ) ? ( bv_8_23_n144 ) : ( n17179 ) ;
assign n17181 =  ( n16517 ) ? ( bv_8_153_n140 ) : ( n17180 ) ;
assign n17182 =  ( n16515 ) ? ( bv_8_58_n136 ) : ( n17181 ) ;
assign n17183 =  ( n16513 ) ? ( bv_8_39_n132 ) : ( n17182 ) ;
assign n17184 =  ( n16511 ) ? ( bv_8_217_n128 ) : ( n17183 ) ;
assign n17185 =  ( n16509 ) ? ( bv_8_235_n83 ) : ( n17184 ) ;
assign n17186 =  ( n16507 ) ? ( bv_8_43_n121 ) : ( n17185 ) ;
assign n17187 =  ( n16505 ) ? ( bv_8_34_n117 ) : ( n17186 ) ;
assign n17188 =  ( n16503 ) ? ( bv_8_210_n113 ) : ( n17187 ) ;
assign n17189 =  ( n16501 ) ? ( bv_8_169_n109 ) : ( n17188 ) ;
assign n17190 =  ( n16499 ) ? ( bv_8_7_n105 ) : ( n17189 ) ;
assign n17191 =  ( n16497 ) ? ( bv_8_51_n101 ) : ( n17190 ) ;
assign n17192 =  ( n16495 ) ? ( bv_8_45_n97 ) : ( n17191 ) ;
assign n17193 =  ( n16493 ) ? ( bv_8_60_n93 ) : ( n17192 ) ;
assign n17194 =  ( n16491 ) ? ( bv_8_21_n89 ) : ( n17193 ) ;
assign n17195 =  ( n16489 ) ? ( bv_8_201_n85 ) : ( n17194 ) ;
assign n17196 =  ( n16487 ) ? ( bv_8_135_n81 ) : ( n17195 ) ;
assign n17197 =  ( n16485 ) ? ( bv_8_170_n77 ) : ( n17196 ) ;
assign n17198 =  ( n16483 ) ? ( bv_8_80_n73 ) : ( n17197 ) ;
assign n17199 =  ( n16481 ) ? ( bv_8_165_n69 ) : ( n17198 ) ;
assign n17200 =  ( n16479 ) ? ( bv_8_3_n65 ) : ( n17199 ) ;
assign n17201 =  ( n16477 ) ? ( bv_8_89_n61 ) : ( n17200 ) ;
assign n17202 =  ( n16475 ) ? ( bv_8_9_n57 ) : ( n17201 ) ;
assign n17203 =  ( n16473 ) ? ( bv_8_26_n53 ) : ( n17202 ) ;
assign n17204 =  ( n16471 ) ? ( bv_8_101_n49 ) : ( n17203 ) ;
assign n17205 =  ( n16469 ) ? ( bv_8_215_n45 ) : ( n17204 ) ;
assign n17206 =  ( n16467 ) ? ( bv_8_132_n41 ) : ( n17205 ) ;
assign n17207 =  ( n16465 ) ? ( bv_8_208_n37 ) : ( n17206 ) ;
assign n17208 =  ( n16463 ) ? ( bv_8_130_n33 ) : ( n17207 ) ;
assign n17209 =  ( n16461 ) ? ( bv_8_41_n29 ) : ( n17208 ) ;
assign n17210 =  ( n16459 ) ? ( bv_8_90_n25 ) : ( n17209 ) ;
assign n17211 =  ( n16457 ) ? ( bv_8_30_n21 ) : ( n17210 ) ;
assign n17212 =  ( n16455 ) ? ( bv_8_123_n17 ) : ( n17211 ) ;
assign n17213 =  ( n16453 ) ? ( bv_8_168_n13 ) : ( n17212 ) ;
assign n17214 =  ( n16451 ) ? ( bv_8_109_n9 ) : ( n17213 ) ;
assign n17215 =  ( n16449 ) ? ( bv_8_44_n5 ) : ( n17214 ) ;
assign n17216 =  ( n13368 ) ^ ( n17215 )  ;
assign n17217 =  ( n17216 ) ^ ( n14136 )  ;
assign n17218 = state_in[63:56] ;
assign n17219 =  ( n17218 ) == ( bv_8_255_n3 )  ;
assign n17220 = state_in[63:56] ;
assign n17221 =  ( n17220 ) == ( bv_8_254_n7 )  ;
assign n17222 = state_in[63:56] ;
assign n17223 =  ( n17222 ) == ( bv_8_253_n11 )  ;
assign n17224 = state_in[63:56] ;
assign n17225 =  ( n17224 ) == ( bv_8_252_n15 )  ;
assign n17226 = state_in[63:56] ;
assign n17227 =  ( n17226 ) == ( bv_8_251_n19 )  ;
assign n17228 = state_in[63:56] ;
assign n17229 =  ( n17228 ) == ( bv_8_250_n23 )  ;
assign n17230 = state_in[63:56] ;
assign n17231 =  ( n17230 ) == ( bv_8_249_n27 )  ;
assign n17232 = state_in[63:56] ;
assign n17233 =  ( n17232 ) == ( bv_8_248_n31 )  ;
assign n17234 = state_in[63:56] ;
assign n17235 =  ( n17234 ) == ( bv_8_247_n35 )  ;
assign n17236 = state_in[63:56] ;
assign n17237 =  ( n17236 ) == ( bv_8_246_n39 )  ;
assign n17238 = state_in[63:56] ;
assign n17239 =  ( n17238 ) == ( bv_8_245_n43 )  ;
assign n17240 = state_in[63:56] ;
assign n17241 =  ( n17240 ) == ( bv_8_244_n47 )  ;
assign n17242 = state_in[63:56] ;
assign n17243 =  ( n17242 ) == ( bv_8_243_n51 )  ;
assign n17244 = state_in[63:56] ;
assign n17245 =  ( n17244 ) == ( bv_8_242_n55 )  ;
assign n17246 = state_in[63:56] ;
assign n17247 =  ( n17246 ) == ( bv_8_241_n59 )  ;
assign n17248 = state_in[63:56] ;
assign n17249 =  ( n17248 ) == ( bv_8_240_n63 )  ;
assign n17250 = state_in[63:56] ;
assign n17251 =  ( n17250 ) == ( bv_8_239_n67 )  ;
assign n17252 = state_in[63:56] ;
assign n17253 =  ( n17252 ) == ( bv_8_238_n71 )  ;
assign n17254 = state_in[63:56] ;
assign n17255 =  ( n17254 ) == ( bv_8_237_n75 )  ;
assign n17256 = state_in[63:56] ;
assign n17257 =  ( n17256 ) == ( bv_8_236_n79 )  ;
assign n17258 = state_in[63:56] ;
assign n17259 =  ( n17258 ) == ( bv_8_235_n83 )  ;
assign n17260 = state_in[63:56] ;
assign n17261 =  ( n17260 ) == ( bv_8_234_n87 )  ;
assign n17262 = state_in[63:56] ;
assign n17263 =  ( n17262 ) == ( bv_8_233_n91 )  ;
assign n17264 = state_in[63:56] ;
assign n17265 =  ( n17264 ) == ( bv_8_232_n95 )  ;
assign n17266 = state_in[63:56] ;
assign n17267 =  ( n17266 ) == ( bv_8_231_n99 )  ;
assign n17268 = state_in[63:56] ;
assign n17269 =  ( n17268 ) == ( bv_8_230_n103 )  ;
assign n17270 = state_in[63:56] ;
assign n17271 =  ( n17270 ) == ( bv_8_229_n107 )  ;
assign n17272 = state_in[63:56] ;
assign n17273 =  ( n17272 ) == ( bv_8_228_n111 )  ;
assign n17274 = state_in[63:56] ;
assign n17275 =  ( n17274 ) == ( bv_8_227_n115 )  ;
assign n17276 = state_in[63:56] ;
assign n17277 =  ( n17276 ) == ( bv_8_226_n119 )  ;
assign n17278 = state_in[63:56] ;
assign n17279 =  ( n17278 ) == ( bv_8_225_n123 )  ;
assign n17280 = state_in[63:56] ;
assign n17281 =  ( n17280 ) == ( bv_8_224_n126 )  ;
assign n17282 = state_in[63:56] ;
assign n17283 =  ( n17282 ) == ( bv_8_223_n130 )  ;
assign n17284 = state_in[63:56] ;
assign n17285 =  ( n17284 ) == ( bv_8_222_n134 )  ;
assign n17286 = state_in[63:56] ;
assign n17287 =  ( n17286 ) == ( bv_8_221_n138 )  ;
assign n17288 = state_in[63:56] ;
assign n17289 =  ( n17288 ) == ( bv_8_220_n142 )  ;
assign n17290 = state_in[63:56] ;
assign n17291 =  ( n17290 ) == ( bv_8_219_n146 )  ;
assign n17292 = state_in[63:56] ;
assign n17293 =  ( n17292 ) == ( bv_8_218_n150 )  ;
assign n17294 = state_in[63:56] ;
assign n17295 =  ( n17294 ) == ( bv_8_217_n128 )  ;
assign n17296 = state_in[63:56] ;
assign n17297 =  ( n17296 ) == ( bv_8_216_n157 )  ;
assign n17298 = state_in[63:56] ;
assign n17299 =  ( n17298 ) == ( bv_8_215_n45 )  ;
assign n17300 = state_in[63:56] ;
assign n17301 =  ( n17300 ) == ( bv_8_214_n164 )  ;
assign n17302 = state_in[63:56] ;
assign n17303 =  ( n17302 ) == ( bv_8_213_n167 )  ;
assign n17304 = state_in[63:56] ;
assign n17305 =  ( n17304 ) == ( bv_8_212_n171 )  ;
assign n17306 = state_in[63:56] ;
assign n17307 =  ( n17306 ) == ( bv_8_211_n175 )  ;
assign n17308 = state_in[63:56] ;
assign n17309 =  ( n17308 ) == ( bv_8_210_n113 )  ;
assign n17310 = state_in[63:56] ;
assign n17311 =  ( n17310 ) == ( bv_8_209_n182 )  ;
assign n17312 = state_in[63:56] ;
assign n17313 =  ( n17312 ) == ( bv_8_208_n37 )  ;
assign n17314 = state_in[63:56] ;
assign n17315 =  ( n17314 ) == ( bv_8_207_n188 )  ;
assign n17316 = state_in[63:56] ;
assign n17317 =  ( n17316 ) == ( bv_8_206_n192 )  ;
assign n17318 = state_in[63:56] ;
assign n17319 =  ( n17318 ) == ( bv_8_205_n196 )  ;
assign n17320 = state_in[63:56] ;
assign n17321 =  ( n17320 ) == ( bv_8_204_n177 )  ;
assign n17322 = state_in[63:56] ;
assign n17323 =  ( n17322 ) == ( bv_8_203_n203 )  ;
assign n17324 = state_in[63:56] ;
assign n17325 =  ( n17324 ) == ( bv_8_202_n207 )  ;
assign n17326 = state_in[63:56] ;
assign n17327 =  ( n17326 ) == ( bv_8_201_n85 )  ;
assign n17328 = state_in[63:56] ;
assign n17329 =  ( n17328 ) == ( bv_8_200_n213 )  ;
assign n17330 = state_in[63:56] ;
assign n17331 =  ( n17330 ) == ( bv_8_199_n216 )  ;
assign n17332 = state_in[63:56] ;
assign n17333 =  ( n17332 ) == ( bv_8_198_n220 )  ;
assign n17334 = state_in[63:56] ;
assign n17335 =  ( n17334 ) == ( bv_8_197_n224 )  ;
assign n17336 = state_in[63:56] ;
assign n17337 =  ( n17336 ) == ( bv_8_196_n228 )  ;
assign n17338 = state_in[63:56] ;
assign n17339 =  ( n17338 ) == ( bv_8_195_n232 )  ;
assign n17340 = state_in[63:56] ;
assign n17341 =  ( n17340 ) == ( bv_8_194_n159 )  ;
assign n17342 = state_in[63:56] ;
assign n17343 =  ( n17342 ) == ( bv_8_193_n239 )  ;
assign n17344 = state_in[63:56] ;
assign n17345 =  ( n17344 ) == ( bv_8_192_n242 )  ;
assign n17346 = state_in[63:56] ;
assign n17347 =  ( n17346 ) == ( bv_8_191_n246 )  ;
assign n17348 = state_in[63:56] ;
assign n17349 =  ( n17348 ) == ( bv_8_190_n250 )  ;
assign n17350 = state_in[63:56] ;
assign n17351 =  ( n17350 ) == ( bv_8_189_n254 )  ;
assign n17352 = state_in[63:56] ;
assign n17353 =  ( n17352 ) == ( bv_8_188_n257 )  ;
assign n17354 = state_in[63:56] ;
assign n17355 =  ( n17354 ) == ( bv_8_187_n260 )  ;
assign n17356 = state_in[63:56] ;
assign n17357 =  ( n17356 ) == ( bv_8_186_n263 )  ;
assign n17358 = state_in[63:56] ;
assign n17359 =  ( n17358 ) == ( bv_8_185_n266 )  ;
assign n17360 = state_in[63:56] ;
assign n17361 =  ( n17360 ) == ( bv_8_184_n270 )  ;
assign n17362 = state_in[63:56] ;
assign n17363 =  ( n17362 ) == ( bv_8_183_n273 )  ;
assign n17364 = state_in[63:56] ;
assign n17365 =  ( n17364 ) == ( bv_8_182_n277 )  ;
assign n17366 = state_in[63:56] ;
assign n17367 =  ( n17366 ) == ( bv_8_181_n281 )  ;
assign n17368 = state_in[63:56] ;
assign n17369 =  ( n17368 ) == ( bv_8_180_n285 )  ;
assign n17370 = state_in[63:56] ;
assign n17371 =  ( n17370 ) == ( bv_8_179_n289 )  ;
assign n17372 = state_in[63:56] ;
assign n17373 =  ( n17372 ) == ( bv_8_178_n292 )  ;
assign n17374 = state_in[63:56] ;
assign n17375 =  ( n17374 ) == ( bv_8_177_n283 )  ;
assign n17376 = state_in[63:56] ;
assign n17377 =  ( n17376 ) == ( bv_8_176_n299 )  ;
assign n17378 = state_in[63:56] ;
assign n17379 =  ( n17378 ) == ( bv_8_175_n302 )  ;
assign n17380 = state_in[63:56] ;
assign n17381 =  ( n17380 ) == ( bv_8_174_n152 )  ;
assign n17382 = state_in[63:56] ;
assign n17383 =  ( n17382 ) == ( bv_8_173_n307 )  ;
assign n17384 = state_in[63:56] ;
assign n17385 =  ( n17384 ) == ( bv_8_172_n268 )  ;
assign n17386 = state_in[63:56] ;
assign n17387 =  ( n17386 ) == ( bv_8_171_n314 )  ;
assign n17388 = state_in[63:56] ;
assign n17389 =  ( n17388 ) == ( bv_8_170_n77 )  ;
assign n17390 = state_in[63:56] ;
assign n17391 =  ( n17390 ) == ( bv_8_169_n109 )  ;
assign n17392 = state_in[63:56] ;
assign n17393 =  ( n17392 ) == ( bv_8_168_n13 )  ;
assign n17394 = state_in[63:56] ;
assign n17395 =  ( n17394 ) == ( bv_8_167_n325 )  ;
assign n17396 = state_in[63:56] ;
assign n17397 =  ( n17396 ) == ( bv_8_166_n328 )  ;
assign n17398 = state_in[63:56] ;
assign n17399 =  ( n17398 ) == ( bv_8_165_n69 )  ;
assign n17400 = state_in[63:56] ;
assign n17401 =  ( n17400 ) == ( bv_8_164_n335 )  ;
assign n17402 = state_in[63:56] ;
assign n17403 =  ( n17402 ) == ( bv_8_163_n339 )  ;
assign n17404 = state_in[63:56] ;
assign n17405 =  ( n17404 ) == ( bv_8_162_n343 )  ;
assign n17406 = state_in[63:56] ;
assign n17407 =  ( n17406 ) == ( bv_8_161_n211 )  ;
assign n17408 = state_in[63:56] ;
assign n17409 =  ( n17408 ) == ( bv_8_160_n350 )  ;
assign n17410 = state_in[63:56] ;
assign n17411 =  ( n17410 ) == ( bv_8_159_n323 )  ;
assign n17412 = state_in[63:56] ;
assign n17413 =  ( n17412 ) == ( bv_8_158_n355 )  ;
assign n17414 = state_in[63:56] ;
assign n17415 =  ( n17414 ) == ( bv_8_157_n359 )  ;
assign n17416 = state_in[63:56] ;
assign n17417 =  ( n17416 ) == ( bv_8_156_n279 )  ;
assign n17418 = state_in[63:56] ;
assign n17419 =  ( n17418 ) == ( bv_8_155_n364 )  ;
assign n17420 = state_in[63:56] ;
assign n17421 =  ( n17420 ) == ( bv_8_154_n368 )  ;
assign n17422 = state_in[63:56] ;
assign n17423 =  ( n17422 ) == ( bv_8_153_n140 )  ;
assign n17424 = state_in[63:56] ;
assign n17425 =  ( n17424 ) == ( bv_8_152_n374 )  ;
assign n17426 = state_in[63:56] ;
assign n17427 =  ( n17426 ) == ( bv_8_151_n218 )  ;
assign n17428 = state_in[63:56] ;
assign n17429 =  ( n17428 ) == ( bv_8_150_n201 )  ;
assign n17430 = state_in[63:56] ;
assign n17431 =  ( n17430 ) == ( bv_8_149_n384 )  ;
assign n17432 = state_in[63:56] ;
assign n17433 =  ( n17432 ) == ( bv_8_148_n388 )  ;
assign n17434 = state_in[63:56] ;
assign n17435 =  ( n17434 ) == ( bv_8_147_n392 )  ;
assign n17436 = state_in[63:56] ;
assign n17437 =  ( n17436 ) == ( bv_8_146_n337 )  ;
assign n17438 = state_in[63:56] ;
assign n17439 =  ( n17438 ) == ( bv_8_145_n397 )  ;
assign n17440 = state_in[63:56] ;
assign n17441 =  ( n17440 ) == ( bv_8_144_n173 )  ;
assign n17442 = state_in[63:56] ;
assign n17443 =  ( n17442 ) == ( bv_8_143_n403 )  ;
assign n17444 = state_in[63:56] ;
assign n17445 =  ( n17444 ) == ( bv_8_142_n406 )  ;
assign n17446 = state_in[63:56] ;
assign n17447 =  ( n17446 ) == ( bv_8_141_n410 )  ;
assign n17448 = state_in[63:56] ;
assign n17449 =  ( n17448 ) == ( bv_8_140_n376 )  ;
assign n17450 = state_in[63:56] ;
assign n17451 =  ( n17450 ) == ( bv_8_139_n297 )  ;
assign n17452 = state_in[63:56] ;
assign n17453 =  ( n17452 ) == ( bv_8_138_n418 )  ;
assign n17454 = state_in[63:56] ;
assign n17455 =  ( n17454 ) == ( bv_8_137_n421 )  ;
assign n17456 = state_in[63:56] ;
assign n17457 =  ( n17456 ) == ( bv_8_136_n425 )  ;
assign n17458 = state_in[63:56] ;
assign n17459 =  ( n17458 ) == ( bv_8_135_n81 )  ;
assign n17460 = state_in[63:56] ;
assign n17461 =  ( n17460 ) == ( bv_8_134_n431 )  ;
assign n17462 = state_in[63:56] ;
assign n17463 =  ( n17462 ) == ( bv_8_133_n434 )  ;
assign n17464 = state_in[63:56] ;
assign n17465 =  ( n17464 ) == ( bv_8_132_n41 )  ;
assign n17466 = state_in[63:56] ;
assign n17467 =  ( n17466 ) == ( bv_8_131_n440 )  ;
assign n17468 = state_in[63:56] ;
assign n17469 =  ( n17468 ) == ( bv_8_130_n33 )  ;
assign n17470 = state_in[63:56] ;
assign n17471 =  ( n17470 ) == ( bv_8_129_n446 )  ;
assign n17472 = state_in[63:56] ;
assign n17473 =  ( n17472 ) == ( bv_8_128_n450 )  ;
assign n17474 = state_in[63:56] ;
assign n17475 =  ( n17474 ) == ( bv_8_127_n453 )  ;
assign n17476 = state_in[63:56] ;
assign n17477 =  ( n17476 ) == ( bv_8_126_n456 )  ;
assign n17478 = state_in[63:56] ;
assign n17479 =  ( n17478 ) == ( bv_8_125_n459 )  ;
assign n17480 = state_in[63:56] ;
assign n17481 =  ( n17480 ) == ( bv_8_124_n184 )  ;
assign n17482 = state_in[63:56] ;
assign n17483 =  ( n17482 ) == ( bv_8_123_n17 )  ;
assign n17484 = state_in[63:56] ;
assign n17485 =  ( n17484 ) == ( bv_8_122_n416 )  ;
assign n17486 = state_in[63:56] ;
assign n17487 =  ( n17486 ) == ( bv_8_121_n470 )  ;
assign n17488 = state_in[63:56] ;
assign n17489 =  ( n17488 ) == ( bv_8_120_n474 )  ;
assign n17490 = state_in[63:56] ;
assign n17491 =  ( n17490 ) == ( bv_8_119_n472 )  ;
assign n17492 = state_in[63:56] ;
assign n17493 =  ( n17492 ) == ( bv_8_118_n480 )  ;
assign n17494 = state_in[63:56] ;
assign n17495 =  ( n17494 ) == ( bv_8_117_n484 )  ;
assign n17496 = state_in[63:56] ;
assign n17497 =  ( n17496 ) == ( bv_8_116_n345 )  ;
assign n17498 = state_in[63:56] ;
assign n17499 =  ( n17498 ) == ( bv_8_115_n222 )  ;
assign n17500 = state_in[63:56] ;
assign n17501 =  ( n17500 ) == ( bv_8_114_n494 )  ;
assign n17502 = state_in[63:56] ;
assign n17503 =  ( n17502 ) == ( bv_8_113_n180 )  ;
assign n17504 = state_in[63:56] ;
assign n17505 =  ( n17504 ) == ( bv_8_112_n482 )  ;
assign n17506 = state_in[63:56] ;
assign n17507 =  ( n17506 ) == ( bv_8_111_n244 )  ;
assign n17508 = state_in[63:56] ;
assign n17509 =  ( n17508 ) == ( bv_8_110_n294 )  ;
assign n17510 = state_in[63:56] ;
assign n17511 =  ( n17510 ) == ( bv_8_109_n9 )  ;
assign n17512 = state_in[63:56] ;
assign n17513 =  ( n17512 ) == ( bv_8_108_n510 )  ;
assign n17514 = state_in[63:56] ;
assign n17515 =  ( n17514 ) == ( bv_8_107_n370 )  ;
assign n17516 = state_in[63:56] ;
assign n17517 =  ( n17516 ) == ( bv_8_106_n155 )  ;
assign n17518 = state_in[63:56] ;
assign n17519 =  ( n17518 ) == ( bv_8_105_n148 )  ;
assign n17520 = state_in[63:56] ;
assign n17521 =  ( n17520 ) == ( bv_8_104_n520 )  ;
assign n17522 = state_in[63:56] ;
assign n17523 =  ( n17522 ) == ( bv_8_103_n523 )  ;
assign n17524 = state_in[63:56] ;
assign n17525 =  ( n17524 ) == ( bv_8_102_n527 )  ;
assign n17526 = state_in[63:56] ;
assign n17527 =  ( n17526 ) == ( bv_8_101_n49 )  ;
assign n17528 = state_in[63:56] ;
assign n17529 =  ( n17528 ) == ( bv_8_100_n348 )  ;
assign n17530 = state_in[63:56] ;
assign n17531 =  ( n17530 ) == ( bv_8_99_n476 )  ;
assign n17532 = state_in[63:56] ;
assign n17533 =  ( n17532 ) == ( bv_8_98_n536 )  ;
assign n17534 = state_in[63:56] ;
assign n17535 =  ( n17534 ) == ( bv_8_97_n198 )  ;
assign n17536 = state_in[63:56] ;
assign n17537 =  ( n17536 ) == ( bv_8_96_n542 )  ;
assign n17538 = state_in[63:56] ;
assign n17539 =  ( n17538 ) == ( bv_8_95_n545 )  ;
assign n17540 = state_in[63:56] ;
assign n17541 =  ( n17540 ) == ( bv_8_94_n548 )  ;
assign n17542 = state_in[63:56] ;
assign n17543 =  ( n17542 ) == ( bv_8_93_n498 )  ;
assign n17544 = state_in[63:56] ;
assign n17545 =  ( n17544 ) == ( bv_8_92_n234 )  ;
assign n17546 = state_in[63:56] ;
assign n17547 =  ( n17546 ) == ( bv_8_91_n555 )  ;
assign n17548 = state_in[63:56] ;
assign n17549 =  ( n17548 ) == ( bv_8_90_n25 )  ;
assign n17550 = state_in[63:56] ;
assign n17551 =  ( n17550 ) == ( bv_8_89_n61 )  ;
assign n17552 = state_in[63:56] ;
assign n17553 =  ( n17552 ) == ( bv_8_88_n562 )  ;
assign n17554 = state_in[63:56] ;
assign n17555 =  ( n17554 ) == ( bv_8_87_n226 )  ;
assign n17556 = state_in[63:56] ;
assign n17557 =  ( n17556 ) == ( bv_8_86_n567 )  ;
assign n17558 = state_in[63:56] ;
assign n17559 =  ( n17558 ) == ( bv_8_85_n423 )  ;
assign n17560 = state_in[63:56] ;
assign n17561 =  ( n17560 ) == ( bv_8_84_n386 )  ;
assign n17562 = state_in[63:56] ;
assign n17563 =  ( n17562 ) == ( bv_8_83_n575 )  ;
assign n17564 = state_in[63:56] ;
assign n17565 =  ( n17564 ) == ( bv_8_82_n578 )  ;
assign n17566 = state_in[63:56] ;
assign n17567 =  ( n17566 ) == ( bv_8_81_n582 )  ;
assign n17568 = state_in[63:56] ;
assign n17569 =  ( n17568 ) == ( bv_8_80_n73 )  ;
assign n17570 = state_in[63:56] ;
assign n17571 =  ( n17570 ) == ( bv_8_79_n538 )  ;
assign n17572 = state_in[63:56] ;
assign n17573 =  ( n17572 ) == ( bv_8_78_n590 )  ;
assign n17574 = state_in[63:56] ;
assign n17575 =  ( n17574 ) == ( bv_8_77_n593 )  ;
assign n17576 = state_in[63:56] ;
assign n17577 =  ( n17576 ) == ( bv_8_76_n596 )  ;
assign n17578 = state_in[63:56] ;
assign n17579 =  ( n17578 ) == ( bv_8_75_n503 )  ;
assign n17580 = state_in[63:56] ;
assign n17581 =  ( n17580 ) == ( bv_8_74_n237 )  ;
assign n17582 = state_in[63:56] ;
assign n17583 =  ( n17582 ) == ( bv_8_73_n275 )  ;
assign n17584 = state_in[63:56] ;
assign n17585 =  ( n17584 ) == ( bv_8_72_n330 )  ;
assign n17586 = state_in[63:56] ;
assign n17587 =  ( n17586 ) == ( bv_8_71_n252 )  ;
assign n17588 = state_in[63:56] ;
assign n17589 =  ( n17588 ) == ( bv_8_70_n609 )  ;
assign n17590 = state_in[63:56] ;
assign n17591 =  ( n17590 ) == ( bv_8_69_n612 )  ;
assign n17592 = state_in[63:56] ;
assign n17593 =  ( n17592 ) == ( bv_8_68_n390 )  ;
assign n17594 = state_in[63:56] ;
assign n17595 =  ( n17594 ) == ( bv_8_67_n318 )  ;
assign n17596 = state_in[63:56] ;
assign n17597 =  ( n17596 ) == ( bv_8_66_n466 )  ;
assign n17598 = state_in[63:56] ;
assign n17599 =  ( n17598 ) == ( bv_8_65_n623 )  ;
assign n17600 = state_in[63:56] ;
assign n17601 =  ( n17600 ) == ( bv_8_64_n573 )  ;
assign n17602 = state_in[63:56] ;
assign n17603 =  ( n17602 ) == ( bv_8_63_n489 )  ;
assign n17604 = state_in[63:56] ;
assign n17605 =  ( n17604 ) == ( bv_8_62_n205 )  ;
assign n17606 = state_in[63:56] ;
assign n17607 =  ( n17606 ) == ( bv_8_61_n634 )  ;
assign n17608 = state_in[63:56] ;
assign n17609 =  ( n17608 ) == ( bv_8_60_n93 )  ;
assign n17610 = state_in[63:56] ;
assign n17611 =  ( n17610 ) == ( bv_8_59_n382 )  ;
assign n17612 = state_in[63:56] ;
assign n17613 =  ( n17612 ) == ( bv_8_58_n136 )  ;
assign n17614 = state_in[63:56] ;
assign n17615 =  ( n17614 ) == ( bv_8_57_n312 )  ;
assign n17616 = state_in[63:56] ;
assign n17617 =  ( n17616 ) == ( bv_8_56_n230 )  ;
assign n17618 = state_in[63:56] ;
assign n17619 =  ( n17618 ) == ( bv_8_55_n650 )  ;
assign n17620 = state_in[63:56] ;
assign n17621 =  ( n17620 ) == ( bv_8_54_n616 )  ;
assign n17622 = state_in[63:56] ;
assign n17623 =  ( n17622 ) == ( bv_8_53_n436 )  ;
assign n17624 = state_in[63:56] ;
assign n17625 =  ( n17624 ) == ( bv_8_52_n619 )  ;
assign n17626 = state_in[63:56] ;
assign n17627 =  ( n17626 ) == ( bv_8_51_n101 )  ;
assign n17628 = state_in[63:56] ;
assign n17629 =  ( n17628 ) == ( bv_8_50_n408 )  ;
assign n17630 = state_in[63:56] ;
assign n17631 =  ( n17630 ) == ( bv_8_49_n309 )  ;
assign n17632 = state_in[63:56] ;
assign n17633 =  ( n17632 ) == ( bv_8_48_n660 )  ;
assign n17634 = state_in[63:56] ;
assign n17635 =  ( n17634 ) == ( bv_8_47_n652 )  ;
assign n17636 = state_in[63:56] ;
assign n17637 =  ( n17636 ) == ( bv_8_46_n429 )  ;
assign n17638 = state_in[63:56] ;
assign n17639 =  ( n17638 ) == ( bv_8_45_n97 )  ;
assign n17640 = state_in[63:56] ;
assign n17641 =  ( n17640 ) == ( bv_8_44_n5 )  ;
assign n17642 = state_in[63:56] ;
assign n17643 =  ( n17642 ) == ( bv_8_43_n121 )  ;
assign n17644 = state_in[63:56] ;
assign n17645 =  ( n17644 ) == ( bv_8_42_n672 )  ;
assign n17646 = state_in[63:56] ;
assign n17647 =  ( n17646 ) == ( bv_8_41_n29 )  ;
assign n17648 = state_in[63:56] ;
assign n17649 =  ( n17648 ) == ( bv_8_40_n366 )  ;
assign n17650 = state_in[63:56] ;
assign n17651 =  ( n17650 ) == ( bv_8_39_n132 )  ;
assign n17652 = state_in[63:56] ;
assign n17653 =  ( n17652 ) == ( bv_8_38_n444 )  ;
assign n17654 = state_in[63:56] ;
assign n17655 =  ( n17654 ) == ( bv_8_37_n506 )  ;
assign n17656 = state_in[63:56] ;
assign n17657 =  ( n17656 ) == ( bv_8_36_n645 )  ;
assign n17658 = state_in[63:56] ;
assign n17659 =  ( n17658 ) == ( bv_8_35_n696 )  ;
assign n17660 = state_in[63:56] ;
assign n17661 =  ( n17660 ) == ( bv_8_34_n117 )  ;
assign n17662 = state_in[63:56] ;
assign n17663 =  ( n17662 ) == ( bv_8_33_n486 )  ;
assign n17664 = state_in[63:56] ;
assign n17665 =  ( n17664 ) == ( bv_8_32_n463 )  ;
assign n17666 = state_in[63:56] ;
assign n17667 =  ( n17666 ) == ( bv_8_31_n705 )  ;
assign n17668 = state_in[63:56] ;
assign n17669 =  ( n17668 ) == ( bv_8_30_n21 )  ;
assign n17670 = state_in[63:56] ;
assign n17671 =  ( n17670 ) == ( bv_8_29_n625 )  ;
assign n17672 = state_in[63:56] ;
assign n17673 =  ( n17672 ) == ( bv_8_28_n162 )  ;
assign n17674 = state_in[63:56] ;
assign n17675 =  ( n17674 ) == ( bv_8_27_n642 )  ;
assign n17676 = state_in[63:56] ;
assign n17677 =  ( n17676 ) == ( bv_8_26_n53 )  ;
assign n17678 = state_in[63:56] ;
assign n17679 =  ( n17678 ) == ( bv_8_25_n399 )  ;
assign n17680 = state_in[63:56] ;
assign n17681 =  ( n17680 ) == ( bv_8_24_n448 )  ;
assign n17682 = state_in[63:56] ;
assign n17683 =  ( n17682 ) == ( bv_8_23_n144 )  ;
assign n17684 = state_in[63:56] ;
assign n17685 =  ( n17684 ) == ( bv_8_22_n357 )  ;
assign n17686 = state_in[63:56] ;
assign n17687 =  ( n17686 ) == ( bv_8_21_n89 )  ;
assign n17688 = state_in[63:56] ;
assign n17689 =  ( n17688 ) == ( bv_8_20_n341 )  ;
assign n17690 = state_in[63:56] ;
assign n17691 =  ( n17690 ) == ( bv_8_19_n588 )  ;
assign n17692 = state_in[63:56] ;
assign n17693 =  ( n17692 ) == ( bv_8_18_n628 )  ;
assign n17694 = state_in[63:56] ;
assign n17695 =  ( n17694 ) == ( bv_8_17_n525 )  ;
assign n17696 = state_in[63:56] ;
assign n17697 =  ( n17696 ) == ( bv_8_16_n248 )  ;
assign n17698 = state_in[63:56] ;
assign n17699 =  ( n17698 ) == ( bv_8_15_n190 )  ;
assign n17700 = state_in[63:56] ;
assign n17701 =  ( n17700 ) == ( bv_8_14_n648 )  ;
assign n17702 = state_in[63:56] ;
assign n17703 =  ( n17702 ) == ( bv_8_13_n194 )  ;
assign n17704 = state_in[63:56] ;
assign n17705 =  ( n17704 ) == ( bv_8_12_n333 )  ;
assign n17706 = state_in[63:56] ;
assign n17707 =  ( n17706 ) == ( bv_8_11_n379 )  ;
assign n17708 = state_in[63:56] ;
assign n17709 =  ( n17708 ) == ( bv_8_10_n655 )  ;
assign n17710 = state_in[63:56] ;
assign n17711 =  ( n17710 ) == ( bv_8_9_n57 )  ;
assign n17712 = state_in[63:56] ;
assign n17713 =  ( n17712 ) == ( bv_8_8_n669 )  ;
assign n17714 = state_in[63:56] ;
assign n17715 =  ( n17714 ) == ( bv_8_7_n105 )  ;
assign n17716 = state_in[63:56] ;
assign n17717 =  ( n17716 ) == ( bv_8_6_n169 )  ;
assign n17718 = state_in[63:56] ;
assign n17719 =  ( n17718 ) == ( bv_8_5_n492 )  ;
assign n17720 = state_in[63:56] ;
assign n17721 =  ( n17720 ) == ( bv_8_4_n516 )  ;
assign n17722 = state_in[63:56] ;
assign n17723 =  ( n17722 ) == ( bv_8_3_n65 )  ;
assign n17724 = state_in[63:56] ;
assign n17725 =  ( n17724 ) == ( bv_8_2_n751 )  ;
assign n17726 = state_in[63:56] ;
assign n17727 =  ( n17726 ) == ( bv_8_1_n287 )  ;
assign n17728 = state_in[63:56] ;
assign n17729 =  ( n17728 ) == ( bv_8_0_n580 )  ;
assign n17730 =  ( n17729 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n17731 =  ( n17727 ) ? ( bv_8_124_n184 ) : ( n17730 ) ;
assign n17732 =  ( n17725 ) ? ( bv_8_119_n472 ) : ( n17731 ) ;
assign n17733 =  ( n17723 ) ? ( bv_8_123_n17 ) : ( n17732 ) ;
assign n17734 =  ( n17721 ) ? ( bv_8_242_n55 ) : ( n17733 ) ;
assign n17735 =  ( n17719 ) ? ( bv_8_107_n370 ) : ( n17734 ) ;
assign n17736 =  ( n17717 ) ? ( bv_8_111_n244 ) : ( n17735 ) ;
assign n17737 =  ( n17715 ) ? ( bv_8_197_n224 ) : ( n17736 ) ;
assign n17738 =  ( n17713 ) ? ( bv_8_48_n660 ) : ( n17737 ) ;
assign n17739 =  ( n17711 ) ? ( bv_8_1_n287 ) : ( n17738 ) ;
assign n17740 =  ( n17709 ) ? ( bv_8_103_n523 ) : ( n17739 ) ;
assign n17741 =  ( n17707 ) ? ( bv_8_43_n121 ) : ( n17740 ) ;
assign n17742 =  ( n17705 ) ? ( bv_8_254_n7 ) : ( n17741 ) ;
assign n17743 =  ( n17703 ) ? ( bv_8_215_n45 ) : ( n17742 ) ;
assign n17744 =  ( n17701 ) ? ( bv_8_171_n314 ) : ( n17743 ) ;
assign n17745 =  ( n17699 ) ? ( bv_8_118_n480 ) : ( n17744 ) ;
assign n17746 =  ( n17697 ) ? ( bv_8_202_n207 ) : ( n17745 ) ;
assign n17747 =  ( n17695 ) ? ( bv_8_130_n33 ) : ( n17746 ) ;
assign n17748 =  ( n17693 ) ? ( bv_8_201_n85 ) : ( n17747 ) ;
assign n17749 =  ( n17691 ) ? ( bv_8_125_n459 ) : ( n17748 ) ;
assign n17750 =  ( n17689 ) ? ( bv_8_250_n23 ) : ( n17749 ) ;
assign n17751 =  ( n17687 ) ? ( bv_8_89_n61 ) : ( n17750 ) ;
assign n17752 =  ( n17685 ) ? ( bv_8_71_n252 ) : ( n17751 ) ;
assign n17753 =  ( n17683 ) ? ( bv_8_240_n63 ) : ( n17752 ) ;
assign n17754 =  ( n17681 ) ? ( bv_8_173_n307 ) : ( n17753 ) ;
assign n17755 =  ( n17679 ) ? ( bv_8_212_n171 ) : ( n17754 ) ;
assign n17756 =  ( n17677 ) ? ( bv_8_162_n343 ) : ( n17755 ) ;
assign n17757 =  ( n17675 ) ? ( bv_8_175_n302 ) : ( n17756 ) ;
assign n17758 =  ( n17673 ) ? ( bv_8_156_n279 ) : ( n17757 ) ;
assign n17759 =  ( n17671 ) ? ( bv_8_164_n335 ) : ( n17758 ) ;
assign n17760 =  ( n17669 ) ? ( bv_8_114_n494 ) : ( n17759 ) ;
assign n17761 =  ( n17667 ) ? ( bv_8_192_n242 ) : ( n17760 ) ;
assign n17762 =  ( n17665 ) ? ( bv_8_183_n273 ) : ( n17761 ) ;
assign n17763 =  ( n17663 ) ? ( bv_8_253_n11 ) : ( n17762 ) ;
assign n17764 =  ( n17661 ) ? ( bv_8_147_n392 ) : ( n17763 ) ;
assign n17765 =  ( n17659 ) ? ( bv_8_38_n444 ) : ( n17764 ) ;
assign n17766 =  ( n17657 ) ? ( bv_8_54_n616 ) : ( n17765 ) ;
assign n17767 =  ( n17655 ) ? ( bv_8_63_n489 ) : ( n17766 ) ;
assign n17768 =  ( n17653 ) ? ( bv_8_247_n35 ) : ( n17767 ) ;
assign n17769 =  ( n17651 ) ? ( bv_8_204_n177 ) : ( n17768 ) ;
assign n17770 =  ( n17649 ) ? ( bv_8_52_n619 ) : ( n17769 ) ;
assign n17771 =  ( n17647 ) ? ( bv_8_165_n69 ) : ( n17770 ) ;
assign n17772 =  ( n17645 ) ? ( bv_8_229_n107 ) : ( n17771 ) ;
assign n17773 =  ( n17643 ) ? ( bv_8_241_n59 ) : ( n17772 ) ;
assign n17774 =  ( n17641 ) ? ( bv_8_113_n180 ) : ( n17773 ) ;
assign n17775 =  ( n17639 ) ? ( bv_8_216_n157 ) : ( n17774 ) ;
assign n17776 =  ( n17637 ) ? ( bv_8_49_n309 ) : ( n17775 ) ;
assign n17777 =  ( n17635 ) ? ( bv_8_21_n89 ) : ( n17776 ) ;
assign n17778 =  ( n17633 ) ? ( bv_8_4_n516 ) : ( n17777 ) ;
assign n17779 =  ( n17631 ) ? ( bv_8_199_n216 ) : ( n17778 ) ;
assign n17780 =  ( n17629 ) ? ( bv_8_35_n696 ) : ( n17779 ) ;
assign n17781 =  ( n17627 ) ? ( bv_8_195_n232 ) : ( n17780 ) ;
assign n17782 =  ( n17625 ) ? ( bv_8_24_n448 ) : ( n17781 ) ;
assign n17783 =  ( n17623 ) ? ( bv_8_150_n201 ) : ( n17782 ) ;
assign n17784 =  ( n17621 ) ? ( bv_8_5_n492 ) : ( n17783 ) ;
assign n17785 =  ( n17619 ) ? ( bv_8_154_n368 ) : ( n17784 ) ;
assign n17786 =  ( n17617 ) ? ( bv_8_7_n105 ) : ( n17785 ) ;
assign n17787 =  ( n17615 ) ? ( bv_8_18_n628 ) : ( n17786 ) ;
assign n17788 =  ( n17613 ) ? ( bv_8_128_n450 ) : ( n17787 ) ;
assign n17789 =  ( n17611 ) ? ( bv_8_226_n119 ) : ( n17788 ) ;
assign n17790 =  ( n17609 ) ? ( bv_8_235_n83 ) : ( n17789 ) ;
assign n17791 =  ( n17607 ) ? ( bv_8_39_n132 ) : ( n17790 ) ;
assign n17792 =  ( n17605 ) ? ( bv_8_178_n292 ) : ( n17791 ) ;
assign n17793 =  ( n17603 ) ? ( bv_8_117_n484 ) : ( n17792 ) ;
assign n17794 =  ( n17601 ) ? ( bv_8_9_n57 ) : ( n17793 ) ;
assign n17795 =  ( n17599 ) ? ( bv_8_131_n440 ) : ( n17794 ) ;
assign n17796 =  ( n17597 ) ? ( bv_8_44_n5 ) : ( n17795 ) ;
assign n17797 =  ( n17595 ) ? ( bv_8_26_n53 ) : ( n17796 ) ;
assign n17798 =  ( n17593 ) ? ( bv_8_27_n642 ) : ( n17797 ) ;
assign n17799 =  ( n17591 ) ? ( bv_8_110_n294 ) : ( n17798 ) ;
assign n17800 =  ( n17589 ) ? ( bv_8_90_n25 ) : ( n17799 ) ;
assign n17801 =  ( n17587 ) ? ( bv_8_160_n350 ) : ( n17800 ) ;
assign n17802 =  ( n17585 ) ? ( bv_8_82_n578 ) : ( n17801 ) ;
assign n17803 =  ( n17583 ) ? ( bv_8_59_n382 ) : ( n17802 ) ;
assign n17804 =  ( n17581 ) ? ( bv_8_214_n164 ) : ( n17803 ) ;
assign n17805 =  ( n17579 ) ? ( bv_8_179_n289 ) : ( n17804 ) ;
assign n17806 =  ( n17577 ) ? ( bv_8_41_n29 ) : ( n17805 ) ;
assign n17807 =  ( n17575 ) ? ( bv_8_227_n115 ) : ( n17806 ) ;
assign n17808 =  ( n17573 ) ? ( bv_8_47_n652 ) : ( n17807 ) ;
assign n17809 =  ( n17571 ) ? ( bv_8_132_n41 ) : ( n17808 ) ;
assign n17810 =  ( n17569 ) ? ( bv_8_83_n575 ) : ( n17809 ) ;
assign n17811 =  ( n17567 ) ? ( bv_8_209_n182 ) : ( n17810 ) ;
assign n17812 =  ( n17565 ) ? ( bv_8_0_n580 ) : ( n17811 ) ;
assign n17813 =  ( n17563 ) ? ( bv_8_237_n75 ) : ( n17812 ) ;
assign n17814 =  ( n17561 ) ? ( bv_8_32_n463 ) : ( n17813 ) ;
assign n17815 =  ( n17559 ) ? ( bv_8_252_n15 ) : ( n17814 ) ;
assign n17816 =  ( n17557 ) ? ( bv_8_177_n283 ) : ( n17815 ) ;
assign n17817 =  ( n17555 ) ? ( bv_8_91_n555 ) : ( n17816 ) ;
assign n17818 =  ( n17553 ) ? ( bv_8_106_n155 ) : ( n17817 ) ;
assign n17819 =  ( n17551 ) ? ( bv_8_203_n203 ) : ( n17818 ) ;
assign n17820 =  ( n17549 ) ? ( bv_8_190_n250 ) : ( n17819 ) ;
assign n17821 =  ( n17547 ) ? ( bv_8_57_n312 ) : ( n17820 ) ;
assign n17822 =  ( n17545 ) ? ( bv_8_74_n237 ) : ( n17821 ) ;
assign n17823 =  ( n17543 ) ? ( bv_8_76_n596 ) : ( n17822 ) ;
assign n17824 =  ( n17541 ) ? ( bv_8_88_n562 ) : ( n17823 ) ;
assign n17825 =  ( n17539 ) ? ( bv_8_207_n188 ) : ( n17824 ) ;
assign n17826 =  ( n17537 ) ? ( bv_8_208_n37 ) : ( n17825 ) ;
assign n17827 =  ( n17535 ) ? ( bv_8_239_n67 ) : ( n17826 ) ;
assign n17828 =  ( n17533 ) ? ( bv_8_170_n77 ) : ( n17827 ) ;
assign n17829 =  ( n17531 ) ? ( bv_8_251_n19 ) : ( n17828 ) ;
assign n17830 =  ( n17529 ) ? ( bv_8_67_n318 ) : ( n17829 ) ;
assign n17831 =  ( n17527 ) ? ( bv_8_77_n593 ) : ( n17830 ) ;
assign n17832 =  ( n17525 ) ? ( bv_8_51_n101 ) : ( n17831 ) ;
assign n17833 =  ( n17523 ) ? ( bv_8_133_n434 ) : ( n17832 ) ;
assign n17834 =  ( n17521 ) ? ( bv_8_69_n612 ) : ( n17833 ) ;
assign n17835 =  ( n17519 ) ? ( bv_8_249_n27 ) : ( n17834 ) ;
assign n17836 =  ( n17517 ) ? ( bv_8_2_n751 ) : ( n17835 ) ;
assign n17837 =  ( n17515 ) ? ( bv_8_127_n453 ) : ( n17836 ) ;
assign n17838 =  ( n17513 ) ? ( bv_8_80_n73 ) : ( n17837 ) ;
assign n17839 =  ( n17511 ) ? ( bv_8_60_n93 ) : ( n17838 ) ;
assign n17840 =  ( n17509 ) ? ( bv_8_159_n323 ) : ( n17839 ) ;
assign n17841 =  ( n17507 ) ? ( bv_8_168_n13 ) : ( n17840 ) ;
assign n17842 =  ( n17505 ) ? ( bv_8_81_n582 ) : ( n17841 ) ;
assign n17843 =  ( n17503 ) ? ( bv_8_163_n339 ) : ( n17842 ) ;
assign n17844 =  ( n17501 ) ? ( bv_8_64_n573 ) : ( n17843 ) ;
assign n17845 =  ( n17499 ) ? ( bv_8_143_n403 ) : ( n17844 ) ;
assign n17846 =  ( n17497 ) ? ( bv_8_146_n337 ) : ( n17845 ) ;
assign n17847 =  ( n17495 ) ? ( bv_8_157_n359 ) : ( n17846 ) ;
assign n17848 =  ( n17493 ) ? ( bv_8_56_n230 ) : ( n17847 ) ;
assign n17849 =  ( n17491 ) ? ( bv_8_245_n43 ) : ( n17848 ) ;
assign n17850 =  ( n17489 ) ? ( bv_8_188_n257 ) : ( n17849 ) ;
assign n17851 =  ( n17487 ) ? ( bv_8_182_n277 ) : ( n17850 ) ;
assign n17852 =  ( n17485 ) ? ( bv_8_218_n150 ) : ( n17851 ) ;
assign n17853 =  ( n17483 ) ? ( bv_8_33_n486 ) : ( n17852 ) ;
assign n17854 =  ( n17481 ) ? ( bv_8_16_n248 ) : ( n17853 ) ;
assign n17855 =  ( n17479 ) ? ( bv_8_255_n3 ) : ( n17854 ) ;
assign n17856 =  ( n17477 ) ? ( bv_8_243_n51 ) : ( n17855 ) ;
assign n17857 =  ( n17475 ) ? ( bv_8_210_n113 ) : ( n17856 ) ;
assign n17858 =  ( n17473 ) ? ( bv_8_205_n196 ) : ( n17857 ) ;
assign n17859 =  ( n17471 ) ? ( bv_8_12_n333 ) : ( n17858 ) ;
assign n17860 =  ( n17469 ) ? ( bv_8_19_n588 ) : ( n17859 ) ;
assign n17861 =  ( n17467 ) ? ( bv_8_236_n79 ) : ( n17860 ) ;
assign n17862 =  ( n17465 ) ? ( bv_8_95_n545 ) : ( n17861 ) ;
assign n17863 =  ( n17463 ) ? ( bv_8_151_n218 ) : ( n17862 ) ;
assign n17864 =  ( n17461 ) ? ( bv_8_68_n390 ) : ( n17863 ) ;
assign n17865 =  ( n17459 ) ? ( bv_8_23_n144 ) : ( n17864 ) ;
assign n17866 =  ( n17457 ) ? ( bv_8_196_n228 ) : ( n17865 ) ;
assign n17867 =  ( n17455 ) ? ( bv_8_167_n325 ) : ( n17866 ) ;
assign n17868 =  ( n17453 ) ? ( bv_8_126_n456 ) : ( n17867 ) ;
assign n17869 =  ( n17451 ) ? ( bv_8_61_n634 ) : ( n17868 ) ;
assign n17870 =  ( n17449 ) ? ( bv_8_100_n348 ) : ( n17869 ) ;
assign n17871 =  ( n17447 ) ? ( bv_8_93_n498 ) : ( n17870 ) ;
assign n17872 =  ( n17445 ) ? ( bv_8_25_n399 ) : ( n17871 ) ;
assign n17873 =  ( n17443 ) ? ( bv_8_115_n222 ) : ( n17872 ) ;
assign n17874 =  ( n17441 ) ? ( bv_8_96_n542 ) : ( n17873 ) ;
assign n17875 =  ( n17439 ) ? ( bv_8_129_n446 ) : ( n17874 ) ;
assign n17876 =  ( n17437 ) ? ( bv_8_79_n538 ) : ( n17875 ) ;
assign n17877 =  ( n17435 ) ? ( bv_8_220_n142 ) : ( n17876 ) ;
assign n17878 =  ( n17433 ) ? ( bv_8_34_n117 ) : ( n17877 ) ;
assign n17879 =  ( n17431 ) ? ( bv_8_42_n672 ) : ( n17878 ) ;
assign n17880 =  ( n17429 ) ? ( bv_8_144_n173 ) : ( n17879 ) ;
assign n17881 =  ( n17427 ) ? ( bv_8_136_n425 ) : ( n17880 ) ;
assign n17882 =  ( n17425 ) ? ( bv_8_70_n609 ) : ( n17881 ) ;
assign n17883 =  ( n17423 ) ? ( bv_8_238_n71 ) : ( n17882 ) ;
assign n17884 =  ( n17421 ) ? ( bv_8_184_n270 ) : ( n17883 ) ;
assign n17885 =  ( n17419 ) ? ( bv_8_20_n341 ) : ( n17884 ) ;
assign n17886 =  ( n17417 ) ? ( bv_8_222_n134 ) : ( n17885 ) ;
assign n17887 =  ( n17415 ) ? ( bv_8_94_n548 ) : ( n17886 ) ;
assign n17888 =  ( n17413 ) ? ( bv_8_11_n379 ) : ( n17887 ) ;
assign n17889 =  ( n17411 ) ? ( bv_8_219_n146 ) : ( n17888 ) ;
assign n17890 =  ( n17409 ) ? ( bv_8_224_n126 ) : ( n17889 ) ;
assign n17891 =  ( n17407 ) ? ( bv_8_50_n408 ) : ( n17890 ) ;
assign n17892 =  ( n17405 ) ? ( bv_8_58_n136 ) : ( n17891 ) ;
assign n17893 =  ( n17403 ) ? ( bv_8_10_n655 ) : ( n17892 ) ;
assign n17894 =  ( n17401 ) ? ( bv_8_73_n275 ) : ( n17893 ) ;
assign n17895 =  ( n17399 ) ? ( bv_8_6_n169 ) : ( n17894 ) ;
assign n17896 =  ( n17397 ) ? ( bv_8_36_n645 ) : ( n17895 ) ;
assign n17897 =  ( n17395 ) ? ( bv_8_92_n234 ) : ( n17896 ) ;
assign n17898 =  ( n17393 ) ? ( bv_8_194_n159 ) : ( n17897 ) ;
assign n17899 =  ( n17391 ) ? ( bv_8_211_n175 ) : ( n17898 ) ;
assign n17900 =  ( n17389 ) ? ( bv_8_172_n268 ) : ( n17899 ) ;
assign n17901 =  ( n17387 ) ? ( bv_8_98_n536 ) : ( n17900 ) ;
assign n17902 =  ( n17385 ) ? ( bv_8_145_n397 ) : ( n17901 ) ;
assign n17903 =  ( n17383 ) ? ( bv_8_149_n384 ) : ( n17902 ) ;
assign n17904 =  ( n17381 ) ? ( bv_8_228_n111 ) : ( n17903 ) ;
assign n17905 =  ( n17379 ) ? ( bv_8_121_n470 ) : ( n17904 ) ;
assign n17906 =  ( n17377 ) ? ( bv_8_231_n99 ) : ( n17905 ) ;
assign n17907 =  ( n17375 ) ? ( bv_8_200_n213 ) : ( n17906 ) ;
assign n17908 =  ( n17373 ) ? ( bv_8_55_n650 ) : ( n17907 ) ;
assign n17909 =  ( n17371 ) ? ( bv_8_109_n9 ) : ( n17908 ) ;
assign n17910 =  ( n17369 ) ? ( bv_8_141_n410 ) : ( n17909 ) ;
assign n17911 =  ( n17367 ) ? ( bv_8_213_n167 ) : ( n17910 ) ;
assign n17912 =  ( n17365 ) ? ( bv_8_78_n590 ) : ( n17911 ) ;
assign n17913 =  ( n17363 ) ? ( bv_8_169_n109 ) : ( n17912 ) ;
assign n17914 =  ( n17361 ) ? ( bv_8_108_n510 ) : ( n17913 ) ;
assign n17915 =  ( n17359 ) ? ( bv_8_86_n567 ) : ( n17914 ) ;
assign n17916 =  ( n17357 ) ? ( bv_8_244_n47 ) : ( n17915 ) ;
assign n17917 =  ( n17355 ) ? ( bv_8_234_n87 ) : ( n17916 ) ;
assign n17918 =  ( n17353 ) ? ( bv_8_101_n49 ) : ( n17917 ) ;
assign n17919 =  ( n17351 ) ? ( bv_8_122_n416 ) : ( n17918 ) ;
assign n17920 =  ( n17349 ) ? ( bv_8_174_n152 ) : ( n17919 ) ;
assign n17921 =  ( n17347 ) ? ( bv_8_8_n669 ) : ( n17920 ) ;
assign n17922 =  ( n17345 ) ? ( bv_8_186_n263 ) : ( n17921 ) ;
assign n17923 =  ( n17343 ) ? ( bv_8_120_n474 ) : ( n17922 ) ;
assign n17924 =  ( n17341 ) ? ( bv_8_37_n506 ) : ( n17923 ) ;
assign n17925 =  ( n17339 ) ? ( bv_8_46_n429 ) : ( n17924 ) ;
assign n17926 =  ( n17337 ) ? ( bv_8_28_n162 ) : ( n17925 ) ;
assign n17927 =  ( n17335 ) ? ( bv_8_166_n328 ) : ( n17926 ) ;
assign n17928 =  ( n17333 ) ? ( bv_8_180_n285 ) : ( n17927 ) ;
assign n17929 =  ( n17331 ) ? ( bv_8_198_n220 ) : ( n17928 ) ;
assign n17930 =  ( n17329 ) ? ( bv_8_232_n95 ) : ( n17929 ) ;
assign n17931 =  ( n17327 ) ? ( bv_8_221_n138 ) : ( n17930 ) ;
assign n17932 =  ( n17325 ) ? ( bv_8_116_n345 ) : ( n17931 ) ;
assign n17933 =  ( n17323 ) ? ( bv_8_31_n705 ) : ( n17932 ) ;
assign n17934 =  ( n17321 ) ? ( bv_8_75_n503 ) : ( n17933 ) ;
assign n17935 =  ( n17319 ) ? ( bv_8_189_n254 ) : ( n17934 ) ;
assign n17936 =  ( n17317 ) ? ( bv_8_139_n297 ) : ( n17935 ) ;
assign n17937 =  ( n17315 ) ? ( bv_8_138_n418 ) : ( n17936 ) ;
assign n17938 =  ( n17313 ) ? ( bv_8_112_n482 ) : ( n17937 ) ;
assign n17939 =  ( n17311 ) ? ( bv_8_62_n205 ) : ( n17938 ) ;
assign n17940 =  ( n17309 ) ? ( bv_8_181_n281 ) : ( n17939 ) ;
assign n17941 =  ( n17307 ) ? ( bv_8_102_n527 ) : ( n17940 ) ;
assign n17942 =  ( n17305 ) ? ( bv_8_72_n330 ) : ( n17941 ) ;
assign n17943 =  ( n17303 ) ? ( bv_8_3_n65 ) : ( n17942 ) ;
assign n17944 =  ( n17301 ) ? ( bv_8_246_n39 ) : ( n17943 ) ;
assign n17945 =  ( n17299 ) ? ( bv_8_14_n648 ) : ( n17944 ) ;
assign n17946 =  ( n17297 ) ? ( bv_8_97_n198 ) : ( n17945 ) ;
assign n17947 =  ( n17295 ) ? ( bv_8_53_n436 ) : ( n17946 ) ;
assign n17948 =  ( n17293 ) ? ( bv_8_87_n226 ) : ( n17947 ) ;
assign n17949 =  ( n17291 ) ? ( bv_8_185_n266 ) : ( n17948 ) ;
assign n17950 =  ( n17289 ) ? ( bv_8_134_n431 ) : ( n17949 ) ;
assign n17951 =  ( n17287 ) ? ( bv_8_193_n239 ) : ( n17950 ) ;
assign n17952 =  ( n17285 ) ? ( bv_8_29_n625 ) : ( n17951 ) ;
assign n17953 =  ( n17283 ) ? ( bv_8_158_n355 ) : ( n17952 ) ;
assign n17954 =  ( n17281 ) ? ( bv_8_225_n123 ) : ( n17953 ) ;
assign n17955 =  ( n17279 ) ? ( bv_8_248_n31 ) : ( n17954 ) ;
assign n17956 =  ( n17277 ) ? ( bv_8_152_n374 ) : ( n17955 ) ;
assign n17957 =  ( n17275 ) ? ( bv_8_17_n525 ) : ( n17956 ) ;
assign n17958 =  ( n17273 ) ? ( bv_8_105_n148 ) : ( n17957 ) ;
assign n17959 =  ( n17271 ) ? ( bv_8_217_n128 ) : ( n17958 ) ;
assign n17960 =  ( n17269 ) ? ( bv_8_142_n406 ) : ( n17959 ) ;
assign n17961 =  ( n17267 ) ? ( bv_8_148_n388 ) : ( n17960 ) ;
assign n17962 =  ( n17265 ) ? ( bv_8_155_n364 ) : ( n17961 ) ;
assign n17963 =  ( n17263 ) ? ( bv_8_30_n21 ) : ( n17962 ) ;
assign n17964 =  ( n17261 ) ? ( bv_8_135_n81 ) : ( n17963 ) ;
assign n17965 =  ( n17259 ) ? ( bv_8_233_n91 ) : ( n17964 ) ;
assign n17966 =  ( n17257 ) ? ( bv_8_206_n192 ) : ( n17965 ) ;
assign n17967 =  ( n17255 ) ? ( bv_8_85_n423 ) : ( n17966 ) ;
assign n17968 =  ( n17253 ) ? ( bv_8_40_n366 ) : ( n17967 ) ;
assign n17969 =  ( n17251 ) ? ( bv_8_223_n130 ) : ( n17968 ) ;
assign n17970 =  ( n17249 ) ? ( bv_8_140_n376 ) : ( n17969 ) ;
assign n17971 =  ( n17247 ) ? ( bv_8_161_n211 ) : ( n17970 ) ;
assign n17972 =  ( n17245 ) ? ( bv_8_137_n421 ) : ( n17971 ) ;
assign n17973 =  ( n17243 ) ? ( bv_8_13_n194 ) : ( n17972 ) ;
assign n17974 =  ( n17241 ) ? ( bv_8_191_n246 ) : ( n17973 ) ;
assign n17975 =  ( n17239 ) ? ( bv_8_230_n103 ) : ( n17974 ) ;
assign n17976 =  ( n17237 ) ? ( bv_8_66_n466 ) : ( n17975 ) ;
assign n17977 =  ( n17235 ) ? ( bv_8_104_n520 ) : ( n17976 ) ;
assign n17978 =  ( n17233 ) ? ( bv_8_65_n623 ) : ( n17977 ) ;
assign n17979 =  ( n17231 ) ? ( bv_8_153_n140 ) : ( n17978 ) ;
assign n17980 =  ( n17229 ) ? ( bv_8_45_n97 ) : ( n17979 ) ;
assign n17981 =  ( n17227 ) ? ( bv_8_15_n190 ) : ( n17980 ) ;
assign n17982 =  ( n17225 ) ? ( bv_8_176_n299 ) : ( n17981 ) ;
assign n17983 =  ( n17223 ) ? ( bv_8_84_n386 ) : ( n17982 ) ;
assign n17984 =  ( n17221 ) ? ( bv_8_187_n260 ) : ( n17983 ) ;
assign n17985 =  ( n17219 ) ? ( bv_8_22_n357 ) : ( n17984 ) ;
assign n17986 =  ( n17217 ) ^ ( n17985 )  ;
assign n17987 =  ( n17986 ) ^ ( n16443 )  ;
assign n17988 = key[55:48] ;
assign n17989 =  ( n17987 ) ^ ( n17988 )  ;
assign n17990 =  { ( n16447 ) , ( n17989 ) }  ;
assign n17991 =  ( n17215 ) ^ ( n14136 )  ;
assign n17992 = state_in[71:64] ;
assign n17993 =  ( n17992 ) == ( bv_8_255_n3 )  ;
assign n17994 = state_in[71:64] ;
assign n17995 =  ( n17994 ) == ( bv_8_254_n7 )  ;
assign n17996 = state_in[71:64] ;
assign n17997 =  ( n17996 ) == ( bv_8_253_n11 )  ;
assign n17998 = state_in[71:64] ;
assign n17999 =  ( n17998 ) == ( bv_8_252_n15 )  ;
assign n18000 = state_in[71:64] ;
assign n18001 =  ( n18000 ) == ( bv_8_251_n19 )  ;
assign n18002 = state_in[71:64] ;
assign n18003 =  ( n18002 ) == ( bv_8_250_n23 )  ;
assign n18004 = state_in[71:64] ;
assign n18005 =  ( n18004 ) == ( bv_8_249_n27 )  ;
assign n18006 = state_in[71:64] ;
assign n18007 =  ( n18006 ) == ( bv_8_248_n31 )  ;
assign n18008 = state_in[71:64] ;
assign n18009 =  ( n18008 ) == ( bv_8_247_n35 )  ;
assign n18010 = state_in[71:64] ;
assign n18011 =  ( n18010 ) == ( bv_8_246_n39 )  ;
assign n18012 = state_in[71:64] ;
assign n18013 =  ( n18012 ) == ( bv_8_245_n43 )  ;
assign n18014 = state_in[71:64] ;
assign n18015 =  ( n18014 ) == ( bv_8_244_n47 )  ;
assign n18016 = state_in[71:64] ;
assign n18017 =  ( n18016 ) == ( bv_8_243_n51 )  ;
assign n18018 = state_in[71:64] ;
assign n18019 =  ( n18018 ) == ( bv_8_242_n55 )  ;
assign n18020 = state_in[71:64] ;
assign n18021 =  ( n18020 ) == ( bv_8_241_n59 )  ;
assign n18022 = state_in[71:64] ;
assign n18023 =  ( n18022 ) == ( bv_8_240_n63 )  ;
assign n18024 = state_in[71:64] ;
assign n18025 =  ( n18024 ) == ( bv_8_239_n67 )  ;
assign n18026 = state_in[71:64] ;
assign n18027 =  ( n18026 ) == ( bv_8_238_n71 )  ;
assign n18028 = state_in[71:64] ;
assign n18029 =  ( n18028 ) == ( bv_8_237_n75 )  ;
assign n18030 = state_in[71:64] ;
assign n18031 =  ( n18030 ) == ( bv_8_236_n79 )  ;
assign n18032 = state_in[71:64] ;
assign n18033 =  ( n18032 ) == ( bv_8_235_n83 )  ;
assign n18034 = state_in[71:64] ;
assign n18035 =  ( n18034 ) == ( bv_8_234_n87 )  ;
assign n18036 = state_in[71:64] ;
assign n18037 =  ( n18036 ) == ( bv_8_233_n91 )  ;
assign n18038 = state_in[71:64] ;
assign n18039 =  ( n18038 ) == ( bv_8_232_n95 )  ;
assign n18040 = state_in[71:64] ;
assign n18041 =  ( n18040 ) == ( bv_8_231_n99 )  ;
assign n18042 = state_in[71:64] ;
assign n18043 =  ( n18042 ) == ( bv_8_230_n103 )  ;
assign n18044 = state_in[71:64] ;
assign n18045 =  ( n18044 ) == ( bv_8_229_n107 )  ;
assign n18046 = state_in[71:64] ;
assign n18047 =  ( n18046 ) == ( bv_8_228_n111 )  ;
assign n18048 = state_in[71:64] ;
assign n18049 =  ( n18048 ) == ( bv_8_227_n115 )  ;
assign n18050 = state_in[71:64] ;
assign n18051 =  ( n18050 ) == ( bv_8_226_n119 )  ;
assign n18052 = state_in[71:64] ;
assign n18053 =  ( n18052 ) == ( bv_8_225_n123 )  ;
assign n18054 = state_in[71:64] ;
assign n18055 =  ( n18054 ) == ( bv_8_224_n126 )  ;
assign n18056 = state_in[71:64] ;
assign n18057 =  ( n18056 ) == ( bv_8_223_n130 )  ;
assign n18058 = state_in[71:64] ;
assign n18059 =  ( n18058 ) == ( bv_8_222_n134 )  ;
assign n18060 = state_in[71:64] ;
assign n18061 =  ( n18060 ) == ( bv_8_221_n138 )  ;
assign n18062 = state_in[71:64] ;
assign n18063 =  ( n18062 ) == ( bv_8_220_n142 )  ;
assign n18064 = state_in[71:64] ;
assign n18065 =  ( n18064 ) == ( bv_8_219_n146 )  ;
assign n18066 = state_in[71:64] ;
assign n18067 =  ( n18066 ) == ( bv_8_218_n150 )  ;
assign n18068 = state_in[71:64] ;
assign n18069 =  ( n18068 ) == ( bv_8_217_n128 )  ;
assign n18070 = state_in[71:64] ;
assign n18071 =  ( n18070 ) == ( bv_8_216_n157 )  ;
assign n18072 = state_in[71:64] ;
assign n18073 =  ( n18072 ) == ( bv_8_215_n45 )  ;
assign n18074 = state_in[71:64] ;
assign n18075 =  ( n18074 ) == ( bv_8_214_n164 )  ;
assign n18076 = state_in[71:64] ;
assign n18077 =  ( n18076 ) == ( bv_8_213_n167 )  ;
assign n18078 = state_in[71:64] ;
assign n18079 =  ( n18078 ) == ( bv_8_212_n171 )  ;
assign n18080 = state_in[71:64] ;
assign n18081 =  ( n18080 ) == ( bv_8_211_n175 )  ;
assign n18082 = state_in[71:64] ;
assign n18083 =  ( n18082 ) == ( bv_8_210_n113 )  ;
assign n18084 = state_in[71:64] ;
assign n18085 =  ( n18084 ) == ( bv_8_209_n182 )  ;
assign n18086 = state_in[71:64] ;
assign n18087 =  ( n18086 ) == ( bv_8_208_n37 )  ;
assign n18088 = state_in[71:64] ;
assign n18089 =  ( n18088 ) == ( bv_8_207_n188 )  ;
assign n18090 = state_in[71:64] ;
assign n18091 =  ( n18090 ) == ( bv_8_206_n192 )  ;
assign n18092 = state_in[71:64] ;
assign n18093 =  ( n18092 ) == ( bv_8_205_n196 )  ;
assign n18094 = state_in[71:64] ;
assign n18095 =  ( n18094 ) == ( bv_8_204_n177 )  ;
assign n18096 = state_in[71:64] ;
assign n18097 =  ( n18096 ) == ( bv_8_203_n203 )  ;
assign n18098 = state_in[71:64] ;
assign n18099 =  ( n18098 ) == ( bv_8_202_n207 )  ;
assign n18100 = state_in[71:64] ;
assign n18101 =  ( n18100 ) == ( bv_8_201_n85 )  ;
assign n18102 = state_in[71:64] ;
assign n18103 =  ( n18102 ) == ( bv_8_200_n213 )  ;
assign n18104 = state_in[71:64] ;
assign n18105 =  ( n18104 ) == ( bv_8_199_n216 )  ;
assign n18106 = state_in[71:64] ;
assign n18107 =  ( n18106 ) == ( bv_8_198_n220 )  ;
assign n18108 = state_in[71:64] ;
assign n18109 =  ( n18108 ) == ( bv_8_197_n224 )  ;
assign n18110 = state_in[71:64] ;
assign n18111 =  ( n18110 ) == ( bv_8_196_n228 )  ;
assign n18112 = state_in[71:64] ;
assign n18113 =  ( n18112 ) == ( bv_8_195_n232 )  ;
assign n18114 = state_in[71:64] ;
assign n18115 =  ( n18114 ) == ( bv_8_194_n159 )  ;
assign n18116 = state_in[71:64] ;
assign n18117 =  ( n18116 ) == ( bv_8_193_n239 )  ;
assign n18118 = state_in[71:64] ;
assign n18119 =  ( n18118 ) == ( bv_8_192_n242 )  ;
assign n18120 = state_in[71:64] ;
assign n18121 =  ( n18120 ) == ( bv_8_191_n246 )  ;
assign n18122 = state_in[71:64] ;
assign n18123 =  ( n18122 ) == ( bv_8_190_n250 )  ;
assign n18124 = state_in[71:64] ;
assign n18125 =  ( n18124 ) == ( bv_8_189_n254 )  ;
assign n18126 = state_in[71:64] ;
assign n18127 =  ( n18126 ) == ( bv_8_188_n257 )  ;
assign n18128 = state_in[71:64] ;
assign n18129 =  ( n18128 ) == ( bv_8_187_n260 )  ;
assign n18130 = state_in[71:64] ;
assign n18131 =  ( n18130 ) == ( bv_8_186_n263 )  ;
assign n18132 = state_in[71:64] ;
assign n18133 =  ( n18132 ) == ( bv_8_185_n266 )  ;
assign n18134 = state_in[71:64] ;
assign n18135 =  ( n18134 ) == ( bv_8_184_n270 )  ;
assign n18136 = state_in[71:64] ;
assign n18137 =  ( n18136 ) == ( bv_8_183_n273 )  ;
assign n18138 = state_in[71:64] ;
assign n18139 =  ( n18138 ) == ( bv_8_182_n277 )  ;
assign n18140 = state_in[71:64] ;
assign n18141 =  ( n18140 ) == ( bv_8_181_n281 )  ;
assign n18142 = state_in[71:64] ;
assign n18143 =  ( n18142 ) == ( bv_8_180_n285 )  ;
assign n18144 = state_in[71:64] ;
assign n18145 =  ( n18144 ) == ( bv_8_179_n289 )  ;
assign n18146 = state_in[71:64] ;
assign n18147 =  ( n18146 ) == ( bv_8_178_n292 )  ;
assign n18148 = state_in[71:64] ;
assign n18149 =  ( n18148 ) == ( bv_8_177_n283 )  ;
assign n18150 = state_in[71:64] ;
assign n18151 =  ( n18150 ) == ( bv_8_176_n299 )  ;
assign n18152 = state_in[71:64] ;
assign n18153 =  ( n18152 ) == ( bv_8_175_n302 )  ;
assign n18154 = state_in[71:64] ;
assign n18155 =  ( n18154 ) == ( bv_8_174_n152 )  ;
assign n18156 = state_in[71:64] ;
assign n18157 =  ( n18156 ) == ( bv_8_173_n307 )  ;
assign n18158 = state_in[71:64] ;
assign n18159 =  ( n18158 ) == ( bv_8_172_n268 )  ;
assign n18160 = state_in[71:64] ;
assign n18161 =  ( n18160 ) == ( bv_8_171_n314 )  ;
assign n18162 = state_in[71:64] ;
assign n18163 =  ( n18162 ) == ( bv_8_170_n77 )  ;
assign n18164 = state_in[71:64] ;
assign n18165 =  ( n18164 ) == ( bv_8_169_n109 )  ;
assign n18166 = state_in[71:64] ;
assign n18167 =  ( n18166 ) == ( bv_8_168_n13 )  ;
assign n18168 = state_in[71:64] ;
assign n18169 =  ( n18168 ) == ( bv_8_167_n325 )  ;
assign n18170 = state_in[71:64] ;
assign n18171 =  ( n18170 ) == ( bv_8_166_n328 )  ;
assign n18172 = state_in[71:64] ;
assign n18173 =  ( n18172 ) == ( bv_8_165_n69 )  ;
assign n18174 = state_in[71:64] ;
assign n18175 =  ( n18174 ) == ( bv_8_164_n335 )  ;
assign n18176 = state_in[71:64] ;
assign n18177 =  ( n18176 ) == ( bv_8_163_n339 )  ;
assign n18178 = state_in[71:64] ;
assign n18179 =  ( n18178 ) == ( bv_8_162_n343 )  ;
assign n18180 = state_in[71:64] ;
assign n18181 =  ( n18180 ) == ( bv_8_161_n211 )  ;
assign n18182 = state_in[71:64] ;
assign n18183 =  ( n18182 ) == ( bv_8_160_n350 )  ;
assign n18184 = state_in[71:64] ;
assign n18185 =  ( n18184 ) == ( bv_8_159_n323 )  ;
assign n18186 = state_in[71:64] ;
assign n18187 =  ( n18186 ) == ( bv_8_158_n355 )  ;
assign n18188 = state_in[71:64] ;
assign n18189 =  ( n18188 ) == ( bv_8_157_n359 )  ;
assign n18190 = state_in[71:64] ;
assign n18191 =  ( n18190 ) == ( bv_8_156_n279 )  ;
assign n18192 = state_in[71:64] ;
assign n18193 =  ( n18192 ) == ( bv_8_155_n364 )  ;
assign n18194 = state_in[71:64] ;
assign n18195 =  ( n18194 ) == ( bv_8_154_n368 )  ;
assign n18196 = state_in[71:64] ;
assign n18197 =  ( n18196 ) == ( bv_8_153_n140 )  ;
assign n18198 = state_in[71:64] ;
assign n18199 =  ( n18198 ) == ( bv_8_152_n374 )  ;
assign n18200 = state_in[71:64] ;
assign n18201 =  ( n18200 ) == ( bv_8_151_n218 )  ;
assign n18202 = state_in[71:64] ;
assign n18203 =  ( n18202 ) == ( bv_8_150_n201 )  ;
assign n18204 = state_in[71:64] ;
assign n18205 =  ( n18204 ) == ( bv_8_149_n384 )  ;
assign n18206 = state_in[71:64] ;
assign n18207 =  ( n18206 ) == ( bv_8_148_n388 )  ;
assign n18208 = state_in[71:64] ;
assign n18209 =  ( n18208 ) == ( bv_8_147_n392 )  ;
assign n18210 = state_in[71:64] ;
assign n18211 =  ( n18210 ) == ( bv_8_146_n337 )  ;
assign n18212 = state_in[71:64] ;
assign n18213 =  ( n18212 ) == ( bv_8_145_n397 )  ;
assign n18214 = state_in[71:64] ;
assign n18215 =  ( n18214 ) == ( bv_8_144_n173 )  ;
assign n18216 = state_in[71:64] ;
assign n18217 =  ( n18216 ) == ( bv_8_143_n403 )  ;
assign n18218 = state_in[71:64] ;
assign n18219 =  ( n18218 ) == ( bv_8_142_n406 )  ;
assign n18220 = state_in[71:64] ;
assign n18221 =  ( n18220 ) == ( bv_8_141_n410 )  ;
assign n18222 = state_in[71:64] ;
assign n18223 =  ( n18222 ) == ( bv_8_140_n376 )  ;
assign n18224 = state_in[71:64] ;
assign n18225 =  ( n18224 ) == ( bv_8_139_n297 )  ;
assign n18226 = state_in[71:64] ;
assign n18227 =  ( n18226 ) == ( bv_8_138_n418 )  ;
assign n18228 = state_in[71:64] ;
assign n18229 =  ( n18228 ) == ( bv_8_137_n421 )  ;
assign n18230 = state_in[71:64] ;
assign n18231 =  ( n18230 ) == ( bv_8_136_n425 )  ;
assign n18232 = state_in[71:64] ;
assign n18233 =  ( n18232 ) == ( bv_8_135_n81 )  ;
assign n18234 = state_in[71:64] ;
assign n18235 =  ( n18234 ) == ( bv_8_134_n431 )  ;
assign n18236 = state_in[71:64] ;
assign n18237 =  ( n18236 ) == ( bv_8_133_n434 )  ;
assign n18238 = state_in[71:64] ;
assign n18239 =  ( n18238 ) == ( bv_8_132_n41 )  ;
assign n18240 = state_in[71:64] ;
assign n18241 =  ( n18240 ) == ( bv_8_131_n440 )  ;
assign n18242 = state_in[71:64] ;
assign n18243 =  ( n18242 ) == ( bv_8_130_n33 )  ;
assign n18244 = state_in[71:64] ;
assign n18245 =  ( n18244 ) == ( bv_8_129_n446 )  ;
assign n18246 = state_in[71:64] ;
assign n18247 =  ( n18246 ) == ( bv_8_128_n450 )  ;
assign n18248 = state_in[71:64] ;
assign n18249 =  ( n18248 ) == ( bv_8_127_n453 )  ;
assign n18250 = state_in[71:64] ;
assign n18251 =  ( n18250 ) == ( bv_8_126_n456 )  ;
assign n18252 = state_in[71:64] ;
assign n18253 =  ( n18252 ) == ( bv_8_125_n459 )  ;
assign n18254 = state_in[71:64] ;
assign n18255 =  ( n18254 ) == ( bv_8_124_n184 )  ;
assign n18256 = state_in[71:64] ;
assign n18257 =  ( n18256 ) == ( bv_8_123_n17 )  ;
assign n18258 = state_in[71:64] ;
assign n18259 =  ( n18258 ) == ( bv_8_122_n416 )  ;
assign n18260 = state_in[71:64] ;
assign n18261 =  ( n18260 ) == ( bv_8_121_n470 )  ;
assign n18262 = state_in[71:64] ;
assign n18263 =  ( n18262 ) == ( bv_8_120_n474 )  ;
assign n18264 = state_in[71:64] ;
assign n18265 =  ( n18264 ) == ( bv_8_119_n472 )  ;
assign n18266 = state_in[71:64] ;
assign n18267 =  ( n18266 ) == ( bv_8_118_n480 )  ;
assign n18268 = state_in[71:64] ;
assign n18269 =  ( n18268 ) == ( bv_8_117_n484 )  ;
assign n18270 = state_in[71:64] ;
assign n18271 =  ( n18270 ) == ( bv_8_116_n345 )  ;
assign n18272 = state_in[71:64] ;
assign n18273 =  ( n18272 ) == ( bv_8_115_n222 )  ;
assign n18274 = state_in[71:64] ;
assign n18275 =  ( n18274 ) == ( bv_8_114_n494 )  ;
assign n18276 = state_in[71:64] ;
assign n18277 =  ( n18276 ) == ( bv_8_113_n180 )  ;
assign n18278 = state_in[71:64] ;
assign n18279 =  ( n18278 ) == ( bv_8_112_n482 )  ;
assign n18280 = state_in[71:64] ;
assign n18281 =  ( n18280 ) == ( bv_8_111_n244 )  ;
assign n18282 = state_in[71:64] ;
assign n18283 =  ( n18282 ) == ( bv_8_110_n294 )  ;
assign n18284 = state_in[71:64] ;
assign n18285 =  ( n18284 ) == ( bv_8_109_n9 )  ;
assign n18286 = state_in[71:64] ;
assign n18287 =  ( n18286 ) == ( bv_8_108_n510 )  ;
assign n18288 = state_in[71:64] ;
assign n18289 =  ( n18288 ) == ( bv_8_107_n370 )  ;
assign n18290 = state_in[71:64] ;
assign n18291 =  ( n18290 ) == ( bv_8_106_n155 )  ;
assign n18292 = state_in[71:64] ;
assign n18293 =  ( n18292 ) == ( bv_8_105_n148 )  ;
assign n18294 = state_in[71:64] ;
assign n18295 =  ( n18294 ) == ( bv_8_104_n520 )  ;
assign n18296 = state_in[71:64] ;
assign n18297 =  ( n18296 ) == ( bv_8_103_n523 )  ;
assign n18298 = state_in[71:64] ;
assign n18299 =  ( n18298 ) == ( bv_8_102_n527 )  ;
assign n18300 = state_in[71:64] ;
assign n18301 =  ( n18300 ) == ( bv_8_101_n49 )  ;
assign n18302 = state_in[71:64] ;
assign n18303 =  ( n18302 ) == ( bv_8_100_n348 )  ;
assign n18304 = state_in[71:64] ;
assign n18305 =  ( n18304 ) == ( bv_8_99_n476 )  ;
assign n18306 = state_in[71:64] ;
assign n18307 =  ( n18306 ) == ( bv_8_98_n536 )  ;
assign n18308 = state_in[71:64] ;
assign n18309 =  ( n18308 ) == ( bv_8_97_n198 )  ;
assign n18310 = state_in[71:64] ;
assign n18311 =  ( n18310 ) == ( bv_8_96_n542 )  ;
assign n18312 = state_in[71:64] ;
assign n18313 =  ( n18312 ) == ( bv_8_95_n545 )  ;
assign n18314 = state_in[71:64] ;
assign n18315 =  ( n18314 ) == ( bv_8_94_n548 )  ;
assign n18316 = state_in[71:64] ;
assign n18317 =  ( n18316 ) == ( bv_8_93_n498 )  ;
assign n18318 = state_in[71:64] ;
assign n18319 =  ( n18318 ) == ( bv_8_92_n234 )  ;
assign n18320 = state_in[71:64] ;
assign n18321 =  ( n18320 ) == ( bv_8_91_n555 )  ;
assign n18322 = state_in[71:64] ;
assign n18323 =  ( n18322 ) == ( bv_8_90_n25 )  ;
assign n18324 = state_in[71:64] ;
assign n18325 =  ( n18324 ) == ( bv_8_89_n61 )  ;
assign n18326 = state_in[71:64] ;
assign n18327 =  ( n18326 ) == ( bv_8_88_n562 )  ;
assign n18328 = state_in[71:64] ;
assign n18329 =  ( n18328 ) == ( bv_8_87_n226 )  ;
assign n18330 = state_in[71:64] ;
assign n18331 =  ( n18330 ) == ( bv_8_86_n567 )  ;
assign n18332 = state_in[71:64] ;
assign n18333 =  ( n18332 ) == ( bv_8_85_n423 )  ;
assign n18334 = state_in[71:64] ;
assign n18335 =  ( n18334 ) == ( bv_8_84_n386 )  ;
assign n18336 = state_in[71:64] ;
assign n18337 =  ( n18336 ) == ( bv_8_83_n575 )  ;
assign n18338 = state_in[71:64] ;
assign n18339 =  ( n18338 ) == ( bv_8_82_n578 )  ;
assign n18340 = state_in[71:64] ;
assign n18341 =  ( n18340 ) == ( bv_8_81_n582 )  ;
assign n18342 = state_in[71:64] ;
assign n18343 =  ( n18342 ) == ( bv_8_80_n73 )  ;
assign n18344 = state_in[71:64] ;
assign n18345 =  ( n18344 ) == ( bv_8_79_n538 )  ;
assign n18346 = state_in[71:64] ;
assign n18347 =  ( n18346 ) == ( bv_8_78_n590 )  ;
assign n18348 = state_in[71:64] ;
assign n18349 =  ( n18348 ) == ( bv_8_77_n593 )  ;
assign n18350 = state_in[71:64] ;
assign n18351 =  ( n18350 ) == ( bv_8_76_n596 )  ;
assign n18352 = state_in[71:64] ;
assign n18353 =  ( n18352 ) == ( bv_8_75_n503 )  ;
assign n18354 = state_in[71:64] ;
assign n18355 =  ( n18354 ) == ( bv_8_74_n237 )  ;
assign n18356 = state_in[71:64] ;
assign n18357 =  ( n18356 ) == ( bv_8_73_n275 )  ;
assign n18358 = state_in[71:64] ;
assign n18359 =  ( n18358 ) == ( bv_8_72_n330 )  ;
assign n18360 = state_in[71:64] ;
assign n18361 =  ( n18360 ) == ( bv_8_71_n252 )  ;
assign n18362 = state_in[71:64] ;
assign n18363 =  ( n18362 ) == ( bv_8_70_n609 )  ;
assign n18364 = state_in[71:64] ;
assign n18365 =  ( n18364 ) == ( bv_8_69_n612 )  ;
assign n18366 = state_in[71:64] ;
assign n18367 =  ( n18366 ) == ( bv_8_68_n390 )  ;
assign n18368 = state_in[71:64] ;
assign n18369 =  ( n18368 ) == ( bv_8_67_n318 )  ;
assign n18370 = state_in[71:64] ;
assign n18371 =  ( n18370 ) == ( bv_8_66_n466 )  ;
assign n18372 = state_in[71:64] ;
assign n18373 =  ( n18372 ) == ( bv_8_65_n623 )  ;
assign n18374 = state_in[71:64] ;
assign n18375 =  ( n18374 ) == ( bv_8_64_n573 )  ;
assign n18376 = state_in[71:64] ;
assign n18377 =  ( n18376 ) == ( bv_8_63_n489 )  ;
assign n18378 = state_in[71:64] ;
assign n18379 =  ( n18378 ) == ( bv_8_62_n205 )  ;
assign n18380 = state_in[71:64] ;
assign n18381 =  ( n18380 ) == ( bv_8_61_n634 )  ;
assign n18382 = state_in[71:64] ;
assign n18383 =  ( n18382 ) == ( bv_8_60_n93 )  ;
assign n18384 = state_in[71:64] ;
assign n18385 =  ( n18384 ) == ( bv_8_59_n382 )  ;
assign n18386 = state_in[71:64] ;
assign n18387 =  ( n18386 ) == ( bv_8_58_n136 )  ;
assign n18388 = state_in[71:64] ;
assign n18389 =  ( n18388 ) == ( bv_8_57_n312 )  ;
assign n18390 = state_in[71:64] ;
assign n18391 =  ( n18390 ) == ( bv_8_56_n230 )  ;
assign n18392 = state_in[71:64] ;
assign n18393 =  ( n18392 ) == ( bv_8_55_n650 )  ;
assign n18394 = state_in[71:64] ;
assign n18395 =  ( n18394 ) == ( bv_8_54_n616 )  ;
assign n18396 = state_in[71:64] ;
assign n18397 =  ( n18396 ) == ( bv_8_53_n436 )  ;
assign n18398 = state_in[71:64] ;
assign n18399 =  ( n18398 ) == ( bv_8_52_n619 )  ;
assign n18400 = state_in[71:64] ;
assign n18401 =  ( n18400 ) == ( bv_8_51_n101 )  ;
assign n18402 = state_in[71:64] ;
assign n18403 =  ( n18402 ) == ( bv_8_50_n408 )  ;
assign n18404 = state_in[71:64] ;
assign n18405 =  ( n18404 ) == ( bv_8_49_n309 )  ;
assign n18406 = state_in[71:64] ;
assign n18407 =  ( n18406 ) == ( bv_8_48_n660 )  ;
assign n18408 = state_in[71:64] ;
assign n18409 =  ( n18408 ) == ( bv_8_47_n652 )  ;
assign n18410 = state_in[71:64] ;
assign n18411 =  ( n18410 ) == ( bv_8_46_n429 )  ;
assign n18412 = state_in[71:64] ;
assign n18413 =  ( n18412 ) == ( bv_8_45_n97 )  ;
assign n18414 = state_in[71:64] ;
assign n18415 =  ( n18414 ) == ( bv_8_44_n5 )  ;
assign n18416 = state_in[71:64] ;
assign n18417 =  ( n18416 ) == ( bv_8_43_n121 )  ;
assign n18418 = state_in[71:64] ;
assign n18419 =  ( n18418 ) == ( bv_8_42_n672 )  ;
assign n18420 = state_in[71:64] ;
assign n18421 =  ( n18420 ) == ( bv_8_41_n29 )  ;
assign n18422 = state_in[71:64] ;
assign n18423 =  ( n18422 ) == ( bv_8_40_n366 )  ;
assign n18424 = state_in[71:64] ;
assign n18425 =  ( n18424 ) == ( bv_8_39_n132 )  ;
assign n18426 = state_in[71:64] ;
assign n18427 =  ( n18426 ) == ( bv_8_38_n444 )  ;
assign n18428 = state_in[71:64] ;
assign n18429 =  ( n18428 ) == ( bv_8_37_n506 )  ;
assign n18430 = state_in[71:64] ;
assign n18431 =  ( n18430 ) == ( bv_8_36_n645 )  ;
assign n18432 = state_in[71:64] ;
assign n18433 =  ( n18432 ) == ( bv_8_35_n696 )  ;
assign n18434 = state_in[71:64] ;
assign n18435 =  ( n18434 ) == ( bv_8_34_n117 )  ;
assign n18436 = state_in[71:64] ;
assign n18437 =  ( n18436 ) == ( bv_8_33_n486 )  ;
assign n18438 = state_in[71:64] ;
assign n18439 =  ( n18438 ) == ( bv_8_32_n463 )  ;
assign n18440 = state_in[71:64] ;
assign n18441 =  ( n18440 ) == ( bv_8_31_n705 )  ;
assign n18442 = state_in[71:64] ;
assign n18443 =  ( n18442 ) == ( bv_8_30_n21 )  ;
assign n18444 = state_in[71:64] ;
assign n18445 =  ( n18444 ) == ( bv_8_29_n625 )  ;
assign n18446 = state_in[71:64] ;
assign n18447 =  ( n18446 ) == ( bv_8_28_n162 )  ;
assign n18448 = state_in[71:64] ;
assign n18449 =  ( n18448 ) == ( bv_8_27_n642 )  ;
assign n18450 = state_in[71:64] ;
assign n18451 =  ( n18450 ) == ( bv_8_26_n53 )  ;
assign n18452 = state_in[71:64] ;
assign n18453 =  ( n18452 ) == ( bv_8_25_n399 )  ;
assign n18454 = state_in[71:64] ;
assign n18455 =  ( n18454 ) == ( bv_8_24_n448 )  ;
assign n18456 = state_in[71:64] ;
assign n18457 =  ( n18456 ) == ( bv_8_23_n144 )  ;
assign n18458 = state_in[71:64] ;
assign n18459 =  ( n18458 ) == ( bv_8_22_n357 )  ;
assign n18460 = state_in[71:64] ;
assign n18461 =  ( n18460 ) == ( bv_8_21_n89 )  ;
assign n18462 = state_in[71:64] ;
assign n18463 =  ( n18462 ) == ( bv_8_20_n341 )  ;
assign n18464 = state_in[71:64] ;
assign n18465 =  ( n18464 ) == ( bv_8_19_n588 )  ;
assign n18466 = state_in[71:64] ;
assign n18467 =  ( n18466 ) == ( bv_8_18_n628 )  ;
assign n18468 = state_in[71:64] ;
assign n18469 =  ( n18468 ) == ( bv_8_17_n525 )  ;
assign n18470 = state_in[71:64] ;
assign n18471 =  ( n18470 ) == ( bv_8_16_n248 )  ;
assign n18472 = state_in[71:64] ;
assign n18473 =  ( n18472 ) == ( bv_8_15_n190 )  ;
assign n18474 = state_in[71:64] ;
assign n18475 =  ( n18474 ) == ( bv_8_14_n648 )  ;
assign n18476 = state_in[71:64] ;
assign n18477 =  ( n18476 ) == ( bv_8_13_n194 )  ;
assign n18478 = state_in[71:64] ;
assign n18479 =  ( n18478 ) == ( bv_8_12_n333 )  ;
assign n18480 = state_in[71:64] ;
assign n18481 =  ( n18480 ) == ( bv_8_11_n379 )  ;
assign n18482 = state_in[71:64] ;
assign n18483 =  ( n18482 ) == ( bv_8_10_n655 )  ;
assign n18484 = state_in[71:64] ;
assign n18485 =  ( n18484 ) == ( bv_8_9_n57 )  ;
assign n18486 = state_in[71:64] ;
assign n18487 =  ( n18486 ) == ( bv_8_8_n669 )  ;
assign n18488 = state_in[71:64] ;
assign n18489 =  ( n18488 ) == ( bv_8_7_n105 )  ;
assign n18490 = state_in[71:64] ;
assign n18491 =  ( n18490 ) == ( bv_8_6_n169 )  ;
assign n18492 = state_in[71:64] ;
assign n18493 =  ( n18492 ) == ( bv_8_5_n492 )  ;
assign n18494 = state_in[71:64] ;
assign n18495 =  ( n18494 ) == ( bv_8_4_n516 )  ;
assign n18496 = state_in[71:64] ;
assign n18497 =  ( n18496 ) == ( bv_8_3_n65 )  ;
assign n18498 = state_in[71:64] ;
assign n18499 =  ( n18498 ) == ( bv_8_2_n751 )  ;
assign n18500 = state_in[71:64] ;
assign n18501 =  ( n18500 ) == ( bv_8_1_n287 )  ;
assign n18502 = state_in[71:64] ;
assign n18503 =  ( n18502 ) == ( bv_8_0_n580 )  ;
assign n18504 =  ( n18503 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n18505 =  ( n18501 ) ? ( bv_8_248_n31 ) : ( n18504 ) ;
assign n18506 =  ( n18499 ) ? ( bv_8_238_n71 ) : ( n18505 ) ;
assign n18507 =  ( n18497 ) ? ( bv_8_246_n39 ) : ( n18506 ) ;
assign n18508 =  ( n18495 ) ? ( bv_8_255_n3 ) : ( n18507 ) ;
assign n18509 =  ( n18493 ) ? ( bv_8_214_n164 ) : ( n18508 ) ;
assign n18510 =  ( n18491 ) ? ( bv_8_222_n134 ) : ( n18509 ) ;
assign n18511 =  ( n18489 ) ? ( bv_8_145_n397 ) : ( n18510 ) ;
assign n18512 =  ( n18487 ) ? ( bv_8_96_n542 ) : ( n18511 ) ;
assign n18513 =  ( n18485 ) ? ( bv_8_2_n751 ) : ( n18512 ) ;
assign n18514 =  ( n18483 ) ? ( bv_8_206_n192 ) : ( n18513 ) ;
assign n18515 =  ( n18481 ) ? ( bv_8_86_n567 ) : ( n18514 ) ;
assign n18516 =  ( n18479 ) ? ( bv_8_231_n99 ) : ( n18515 ) ;
assign n18517 =  ( n18477 ) ? ( bv_8_181_n281 ) : ( n18516 ) ;
assign n18518 =  ( n18475 ) ? ( bv_8_77_n593 ) : ( n18517 ) ;
assign n18519 =  ( n18473 ) ? ( bv_8_236_n79 ) : ( n18518 ) ;
assign n18520 =  ( n18471 ) ? ( bv_8_143_n403 ) : ( n18519 ) ;
assign n18521 =  ( n18469 ) ? ( bv_8_31_n705 ) : ( n18520 ) ;
assign n18522 =  ( n18467 ) ? ( bv_8_137_n421 ) : ( n18521 ) ;
assign n18523 =  ( n18465 ) ? ( bv_8_250_n23 ) : ( n18522 ) ;
assign n18524 =  ( n18463 ) ? ( bv_8_239_n67 ) : ( n18523 ) ;
assign n18525 =  ( n18461 ) ? ( bv_8_178_n292 ) : ( n18524 ) ;
assign n18526 =  ( n18459 ) ? ( bv_8_142_n406 ) : ( n18525 ) ;
assign n18527 =  ( n18457 ) ? ( bv_8_251_n19 ) : ( n18526 ) ;
assign n18528 =  ( n18455 ) ? ( bv_8_65_n623 ) : ( n18527 ) ;
assign n18529 =  ( n18453 ) ? ( bv_8_179_n289 ) : ( n18528 ) ;
assign n18530 =  ( n18451 ) ? ( bv_8_95_n545 ) : ( n18529 ) ;
assign n18531 =  ( n18449 ) ? ( bv_8_69_n612 ) : ( n18530 ) ;
assign n18532 =  ( n18447 ) ? ( bv_8_35_n696 ) : ( n18531 ) ;
assign n18533 =  ( n18445 ) ? ( bv_8_83_n575 ) : ( n18532 ) ;
assign n18534 =  ( n18443 ) ? ( bv_8_228_n111 ) : ( n18533 ) ;
assign n18535 =  ( n18441 ) ? ( bv_8_155_n364 ) : ( n18534 ) ;
assign n18536 =  ( n18439 ) ? ( bv_8_117_n484 ) : ( n18535 ) ;
assign n18537 =  ( n18437 ) ? ( bv_8_225_n123 ) : ( n18536 ) ;
assign n18538 =  ( n18435 ) ? ( bv_8_61_n634 ) : ( n18537 ) ;
assign n18539 =  ( n18433 ) ? ( bv_8_76_n596 ) : ( n18538 ) ;
assign n18540 =  ( n18431 ) ? ( bv_8_108_n510 ) : ( n18539 ) ;
assign n18541 =  ( n18429 ) ? ( bv_8_126_n456 ) : ( n18540 ) ;
assign n18542 =  ( n18427 ) ? ( bv_8_245_n43 ) : ( n18541 ) ;
assign n18543 =  ( n18425 ) ? ( bv_8_131_n440 ) : ( n18542 ) ;
assign n18544 =  ( n18423 ) ? ( bv_8_104_n520 ) : ( n18543 ) ;
assign n18545 =  ( n18421 ) ? ( bv_8_81_n582 ) : ( n18544 ) ;
assign n18546 =  ( n18419 ) ? ( bv_8_209_n182 ) : ( n18545 ) ;
assign n18547 =  ( n18417 ) ? ( bv_8_249_n27 ) : ( n18546 ) ;
assign n18548 =  ( n18415 ) ? ( bv_8_226_n119 ) : ( n18547 ) ;
assign n18549 =  ( n18413 ) ? ( bv_8_171_n314 ) : ( n18548 ) ;
assign n18550 =  ( n18411 ) ? ( bv_8_98_n536 ) : ( n18549 ) ;
assign n18551 =  ( n18409 ) ? ( bv_8_42_n672 ) : ( n18550 ) ;
assign n18552 =  ( n18407 ) ? ( bv_8_8_n669 ) : ( n18551 ) ;
assign n18553 =  ( n18405 ) ? ( bv_8_149_n384 ) : ( n18552 ) ;
assign n18554 =  ( n18403 ) ? ( bv_8_70_n609 ) : ( n18553 ) ;
assign n18555 =  ( n18401 ) ? ( bv_8_157_n359 ) : ( n18554 ) ;
assign n18556 =  ( n18399 ) ? ( bv_8_48_n660 ) : ( n18555 ) ;
assign n18557 =  ( n18397 ) ? ( bv_8_55_n650 ) : ( n18556 ) ;
assign n18558 =  ( n18395 ) ? ( bv_8_10_n655 ) : ( n18557 ) ;
assign n18559 =  ( n18393 ) ? ( bv_8_47_n652 ) : ( n18558 ) ;
assign n18560 =  ( n18391 ) ? ( bv_8_14_n648 ) : ( n18559 ) ;
assign n18561 =  ( n18389 ) ? ( bv_8_36_n645 ) : ( n18560 ) ;
assign n18562 =  ( n18387 ) ? ( bv_8_27_n642 ) : ( n18561 ) ;
assign n18563 =  ( n18385 ) ? ( bv_8_223_n130 ) : ( n18562 ) ;
assign n18564 =  ( n18383 ) ? ( bv_8_205_n196 ) : ( n18563 ) ;
assign n18565 =  ( n18381 ) ? ( bv_8_78_n590 ) : ( n18564 ) ;
assign n18566 =  ( n18379 ) ? ( bv_8_127_n453 ) : ( n18565 ) ;
assign n18567 =  ( n18377 ) ? ( bv_8_234_n87 ) : ( n18566 ) ;
assign n18568 =  ( n18375 ) ? ( bv_8_18_n628 ) : ( n18567 ) ;
assign n18569 =  ( n18373 ) ? ( bv_8_29_n625 ) : ( n18568 ) ;
assign n18570 =  ( n18371 ) ? ( bv_8_88_n562 ) : ( n18569 ) ;
assign n18571 =  ( n18369 ) ? ( bv_8_52_n619 ) : ( n18570 ) ;
assign n18572 =  ( n18367 ) ? ( bv_8_54_n616 ) : ( n18571 ) ;
assign n18573 =  ( n18365 ) ? ( bv_8_220_n142 ) : ( n18572 ) ;
assign n18574 =  ( n18363 ) ? ( bv_8_180_n285 ) : ( n18573 ) ;
assign n18575 =  ( n18361 ) ? ( bv_8_91_n555 ) : ( n18574 ) ;
assign n18576 =  ( n18359 ) ? ( bv_8_164_n335 ) : ( n18575 ) ;
assign n18577 =  ( n18357 ) ? ( bv_8_118_n480 ) : ( n18576 ) ;
assign n18578 =  ( n18355 ) ? ( bv_8_183_n273 ) : ( n18577 ) ;
assign n18579 =  ( n18353 ) ? ( bv_8_125_n459 ) : ( n18578 ) ;
assign n18580 =  ( n18351 ) ? ( bv_8_82_n578 ) : ( n18579 ) ;
assign n18581 =  ( n18349 ) ? ( bv_8_221_n138 ) : ( n18580 ) ;
assign n18582 =  ( n18347 ) ? ( bv_8_94_n548 ) : ( n18581 ) ;
assign n18583 =  ( n18345 ) ? ( bv_8_19_n588 ) : ( n18582 ) ;
assign n18584 =  ( n18343 ) ? ( bv_8_166_n328 ) : ( n18583 ) ;
assign n18585 =  ( n18341 ) ? ( bv_8_185_n266 ) : ( n18584 ) ;
assign n18586 =  ( n18339 ) ? ( bv_8_0_n580 ) : ( n18585 ) ;
assign n18587 =  ( n18337 ) ? ( bv_8_193_n239 ) : ( n18586 ) ;
assign n18588 =  ( n18335 ) ? ( bv_8_64_n573 ) : ( n18587 ) ;
assign n18589 =  ( n18333 ) ? ( bv_8_227_n115 ) : ( n18588 ) ;
assign n18590 =  ( n18331 ) ? ( bv_8_121_n470 ) : ( n18589 ) ;
assign n18591 =  ( n18329 ) ? ( bv_8_182_n277 ) : ( n18590 ) ;
assign n18592 =  ( n18327 ) ? ( bv_8_212_n171 ) : ( n18591 ) ;
assign n18593 =  ( n18325 ) ? ( bv_8_141_n410 ) : ( n18592 ) ;
assign n18594 =  ( n18323 ) ? ( bv_8_103_n523 ) : ( n18593 ) ;
assign n18595 =  ( n18321 ) ? ( bv_8_114_n494 ) : ( n18594 ) ;
assign n18596 =  ( n18319 ) ? ( bv_8_148_n388 ) : ( n18595 ) ;
assign n18597 =  ( n18317 ) ? ( bv_8_152_n374 ) : ( n18596 ) ;
assign n18598 =  ( n18315 ) ? ( bv_8_176_n299 ) : ( n18597 ) ;
assign n18599 =  ( n18313 ) ? ( bv_8_133_n434 ) : ( n18598 ) ;
assign n18600 =  ( n18311 ) ? ( bv_8_187_n260 ) : ( n18599 ) ;
assign n18601 =  ( n18309 ) ? ( bv_8_197_n224 ) : ( n18600 ) ;
assign n18602 =  ( n18307 ) ? ( bv_8_79_n538 ) : ( n18601 ) ;
assign n18603 =  ( n18305 ) ? ( bv_8_237_n75 ) : ( n18602 ) ;
assign n18604 =  ( n18303 ) ? ( bv_8_134_n431 ) : ( n18603 ) ;
assign n18605 =  ( n18301 ) ? ( bv_8_154_n368 ) : ( n18604 ) ;
assign n18606 =  ( n18299 ) ? ( bv_8_102_n527 ) : ( n18605 ) ;
assign n18607 =  ( n18297 ) ? ( bv_8_17_n525 ) : ( n18606 ) ;
assign n18608 =  ( n18295 ) ? ( bv_8_138_n418 ) : ( n18607 ) ;
assign n18609 =  ( n18293 ) ? ( bv_8_233_n91 ) : ( n18608 ) ;
assign n18610 =  ( n18291 ) ? ( bv_8_4_n516 ) : ( n18609 ) ;
assign n18611 =  ( n18289 ) ? ( bv_8_254_n7 ) : ( n18610 ) ;
assign n18612 =  ( n18287 ) ? ( bv_8_160_n350 ) : ( n18611 ) ;
assign n18613 =  ( n18285 ) ? ( bv_8_120_n474 ) : ( n18612 ) ;
assign n18614 =  ( n18283 ) ? ( bv_8_37_n506 ) : ( n18613 ) ;
assign n18615 =  ( n18281 ) ? ( bv_8_75_n503 ) : ( n18614 ) ;
assign n18616 =  ( n18279 ) ? ( bv_8_162_n343 ) : ( n18615 ) ;
assign n18617 =  ( n18277 ) ? ( bv_8_93_n498 ) : ( n18616 ) ;
assign n18618 =  ( n18275 ) ? ( bv_8_128_n450 ) : ( n18617 ) ;
assign n18619 =  ( n18273 ) ? ( bv_8_5_n492 ) : ( n18618 ) ;
assign n18620 =  ( n18271 ) ? ( bv_8_63_n489 ) : ( n18619 ) ;
assign n18621 =  ( n18269 ) ? ( bv_8_33_n486 ) : ( n18620 ) ;
assign n18622 =  ( n18267 ) ? ( bv_8_112_n482 ) : ( n18621 ) ;
assign n18623 =  ( n18265 ) ? ( bv_8_241_n59 ) : ( n18622 ) ;
assign n18624 =  ( n18263 ) ? ( bv_8_99_n476 ) : ( n18623 ) ;
assign n18625 =  ( n18261 ) ? ( bv_8_119_n472 ) : ( n18624 ) ;
assign n18626 =  ( n18259 ) ? ( bv_8_175_n302 ) : ( n18625 ) ;
assign n18627 =  ( n18257 ) ? ( bv_8_66_n466 ) : ( n18626 ) ;
assign n18628 =  ( n18255 ) ? ( bv_8_32_n463 ) : ( n18627 ) ;
assign n18629 =  ( n18253 ) ? ( bv_8_229_n107 ) : ( n18628 ) ;
assign n18630 =  ( n18251 ) ? ( bv_8_253_n11 ) : ( n18629 ) ;
assign n18631 =  ( n18249 ) ? ( bv_8_191_n246 ) : ( n18630 ) ;
assign n18632 =  ( n18247 ) ? ( bv_8_129_n446 ) : ( n18631 ) ;
assign n18633 =  ( n18245 ) ? ( bv_8_24_n448 ) : ( n18632 ) ;
assign n18634 =  ( n18243 ) ? ( bv_8_38_n444 ) : ( n18633 ) ;
assign n18635 =  ( n18241 ) ? ( bv_8_195_n232 ) : ( n18634 ) ;
assign n18636 =  ( n18239 ) ? ( bv_8_190_n250 ) : ( n18635 ) ;
assign n18637 =  ( n18237 ) ? ( bv_8_53_n436 ) : ( n18636 ) ;
assign n18638 =  ( n18235 ) ? ( bv_8_136_n425 ) : ( n18637 ) ;
assign n18639 =  ( n18233 ) ? ( bv_8_46_n429 ) : ( n18638 ) ;
assign n18640 =  ( n18231 ) ? ( bv_8_147_n392 ) : ( n18639 ) ;
assign n18641 =  ( n18229 ) ? ( bv_8_85_n423 ) : ( n18640 ) ;
assign n18642 =  ( n18227 ) ? ( bv_8_252_n15 ) : ( n18641 ) ;
assign n18643 =  ( n18225 ) ? ( bv_8_122_n416 ) : ( n18642 ) ;
assign n18644 =  ( n18223 ) ? ( bv_8_200_n213 ) : ( n18643 ) ;
assign n18645 =  ( n18221 ) ? ( bv_8_186_n263 ) : ( n18644 ) ;
assign n18646 =  ( n18219 ) ? ( bv_8_50_n408 ) : ( n18645 ) ;
assign n18647 =  ( n18217 ) ? ( bv_8_230_n103 ) : ( n18646 ) ;
assign n18648 =  ( n18215 ) ? ( bv_8_192_n242 ) : ( n18647 ) ;
assign n18649 =  ( n18213 ) ? ( bv_8_25_n399 ) : ( n18648 ) ;
assign n18650 =  ( n18211 ) ? ( bv_8_158_n355 ) : ( n18649 ) ;
assign n18651 =  ( n18209 ) ? ( bv_8_163_n339 ) : ( n18650 ) ;
assign n18652 =  ( n18207 ) ? ( bv_8_68_n390 ) : ( n18651 ) ;
assign n18653 =  ( n18205 ) ? ( bv_8_84_n386 ) : ( n18652 ) ;
assign n18654 =  ( n18203 ) ? ( bv_8_59_n382 ) : ( n18653 ) ;
assign n18655 =  ( n18201 ) ? ( bv_8_11_n379 ) : ( n18654 ) ;
assign n18656 =  ( n18199 ) ? ( bv_8_140_n376 ) : ( n18655 ) ;
assign n18657 =  ( n18197 ) ? ( bv_8_199_n216 ) : ( n18656 ) ;
assign n18658 =  ( n18195 ) ? ( bv_8_107_n370 ) : ( n18657 ) ;
assign n18659 =  ( n18193 ) ? ( bv_8_40_n366 ) : ( n18658 ) ;
assign n18660 =  ( n18191 ) ? ( bv_8_167_n325 ) : ( n18659 ) ;
assign n18661 =  ( n18189 ) ? ( bv_8_188_n257 ) : ( n18660 ) ;
assign n18662 =  ( n18187 ) ? ( bv_8_22_n357 ) : ( n18661 ) ;
assign n18663 =  ( n18185 ) ? ( bv_8_173_n307 ) : ( n18662 ) ;
assign n18664 =  ( n18183 ) ? ( bv_8_219_n146 ) : ( n18663 ) ;
assign n18665 =  ( n18181 ) ? ( bv_8_100_n348 ) : ( n18664 ) ;
assign n18666 =  ( n18179 ) ? ( bv_8_116_n345 ) : ( n18665 ) ;
assign n18667 =  ( n18177 ) ? ( bv_8_20_n341 ) : ( n18666 ) ;
assign n18668 =  ( n18175 ) ? ( bv_8_146_n337 ) : ( n18667 ) ;
assign n18669 =  ( n18173 ) ? ( bv_8_12_n333 ) : ( n18668 ) ;
assign n18670 =  ( n18171 ) ? ( bv_8_72_n330 ) : ( n18669 ) ;
assign n18671 =  ( n18169 ) ? ( bv_8_184_n270 ) : ( n18670 ) ;
assign n18672 =  ( n18167 ) ? ( bv_8_159_n323 ) : ( n18671 ) ;
assign n18673 =  ( n18165 ) ? ( bv_8_189_n254 ) : ( n18672 ) ;
assign n18674 =  ( n18163 ) ? ( bv_8_67_n318 ) : ( n18673 ) ;
assign n18675 =  ( n18161 ) ? ( bv_8_196_n228 ) : ( n18674 ) ;
assign n18676 =  ( n18159 ) ? ( bv_8_57_n312 ) : ( n18675 ) ;
assign n18677 =  ( n18157 ) ? ( bv_8_49_n309 ) : ( n18676 ) ;
assign n18678 =  ( n18155 ) ? ( bv_8_211_n175 ) : ( n18677 ) ;
assign n18679 =  ( n18153 ) ? ( bv_8_242_n55 ) : ( n18678 ) ;
assign n18680 =  ( n18151 ) ? ( bv_8_213_n167 ) : ( n18679 ) ;
assign n18681 =  ( n18149 ) ? ( bv_8_139_n297 ) : ( n18680 ) ;
assign n18682 =  ( n18147 ) ? ( bv_8_110_n294 ) : ( n18681 ) ;
assign n18683 =  ( n18145 ) ? ( bv_8_218_n150 ) : ( n18682 ) ;
assign n18684 =  ( n18143 ) ? ( bv_8_1_n287 ) : ( n18683 ) ;
assign n18685 =  ( n18141 ) ? ( bv_8_177_n283 ) : ( n18684 ) ;
assign n18686 =  ( n18139 ) ? ( bv_8_156_n279 ) : ( n18685 ) ;
assign n18687 =  ( n18137 ) ? ( bv_8_73_n275 ) : ( n18686 ) ;
assign n18688 =  ( n18135 ) ? ( bv_8_216_n157 ) : ( n18687 ) ;
assign n18689 =  ( n18133 ) ? ( bv_8_172_n268 ) : ( n18688 ) ;
assign n18690 =  ( n18131 ) ? ( bv_8_243_n51 ) : ( n18689 ) ;
assign n18691 =  ( n18129 ) ? ( bv_8_207_n188 ) : ( n18690 ) ;
assign n18692 =  ( n18127 ) ? ( bv_8_202_n207 ) : ( n18691 ) ;
assign n18693 =  ( n18125 ) ? ( bv_8_244_n47 ) : ( n18692 ) ;
assign n18694 =  ( n18123 ) ? ( bv_8_71_n252 ) : ( n18693 ) ;
assign n18695 =  ( n18121 ) ? ( bv_8_16_n248 ) : ( n18694 ) ;
assign n18696 =  ( n18119 ) ? ( bv_8_111_n244 ) : ( n18695 ) ;
assign n18697 =  ( n18117 ) ? ( bv_8_240_n63 ) : ( n18696 ) ;
assign n18698 =  ( n18115 ) ? ( bv_8_74_n237 ) : ( n18697 ) ;
assign n18699 =  ( n18113 ) ? ( bv_8_92_n234 ) : ( n18698 ) ;
assign n18700 =  ( n18111 ) ? ( bv_8_56_n230 ) : ( n18699 ) ;
assign n18701 =  ( n18109 ) ? ( bv_8_87_n226 ) : ( n18700 ) ;
assign n18702 =  ( n18107 ) ? ( bv_8_115_n222 ) : ( n18701 ) ;
assign n18703 =  ( n18105 ) ? ( bv_8_151_n218 ) : ( n18702 ) ;
assign n18704 =  ( n18103 ) ? ( bv_8_203_n203 ) : ( n18703 ) ;
assign n18705 =  ( n18101 ) ? ( bv_8_161_n211 ) : ( n18704 ) ;
assign n18706 =  ( n18099 ) ? ( bv_8_232_n95 ) : ( n18705 ) ;
assign n18707 =  ( n18097 ) ? ( bv_8_62_n205 ) : ( n18706 ) ;
assign n18708 =  ( n18095 ) ? ( bv_8_150_n201 ) : ( n18707 ) ;
assign n18709 =  ( n18093 ) ? ( bv_8_97_n198 ) : ( n18708 ) ;
assign n18710 =  ( n18091 ) ? ( bv_8_13_n194 ) : ( n18709 ) ;
assign n18711 =  ( n18089 ) ? ( bv_8_15_n190 ) : ( n18710 ) ;
assign n18712 =  ( n18087 ) ? ( bv_8_224_n126 ) : ( n18711 ) ;
assign n18713 =  ( n18085 ) ? ( bv_8_124_n184 ) : ( n18712 ) ;
assign n18714 =  ( n18083 ) ? ( bv_8_113_n180 ) : ( n18713 ) ;
assign n18715 =  ( n18081 ) ? ( bv_8_204_n177 ) : ( n18714 ) ;
assign n18716 =  ( n18079 ) ? ( bv_8_144_n173 ) : ( n18715 ) ;
assign n18717 =  ( n18077 ) ? ( bv_8_6_n169 ) : ( n18716 ) ;
assign n18718 =  ( n18075 ) ? ( bv_8_247_n35 ) : ( n18717 ) ;
assign n18719 =  ( n18073 ) ? ( bv_8_28_n162 ) : ( n18718 ) ;
assign n18720 =  ( n18071 ) ? ( bv_8_194_n159 ) : ( n18719 ) ;
assign n18721 =  ( n18069 ) ? ( bv_8_106_n155 ) : ( n18720 ) ;
assign n18722 =  ( n18067 ) ? ( bv_8_174_n152 ) : ( n18721 ) ;
assign n18723 =  ( n18065 ) ? ( bv_8_105_n148 ) : ( n18722 ) ;
assign n18724 =  ( n18063 ) ? ( bv_8_23_n144 ) : ( n18723 ) ;
assign n18725 =  ( n18061 ) ? ( bv_8_153_n140 ) : ( n18724 ) ;
assign n18726 =  ( n18059 ) ? ( bv_8_58_n136 ) : ( n18725 ) ;
assign n18727 =  ( n18057 ) ? ( bv_8_39_n132 ) : ( n18726 ) ;
assign n18728 =  ( n18055 ) ? ( bv_8_217_n128 ) : ( n18727 ) ;
assign n18729 =  ( n18053 ) ? ( bv_8_235_n83 ) : ( n18728 ) ;
assign n18730 =  ( n18051 ) ? ( bv_8_43_n121 ) : ( n18729 ) ;
assign n18731 =  ( n18049 ) ? ( bv_8_34_n117 ) : ( n18730 ) ;
assign n18732 =  ( n18047 ) ? ( bv_8_210_n113 ) : ( n18731 ) ;
assign n18733 =  ( n18045 ) ? ( bv_8_169_n109 ) : ( n18732 ) ;
assign n18734 =  ( n18043 ) ? ( bv_8_7_n105 ) : ( n18733 ) ;
assign n18735 =  ( n18041 ) ? ( bv_8_51_n101 ) : ( n18734 ) ;
assign n18736 =  ( n18039 ) ? ( bv_8_45_n97 ) : ( n18735 ) ;
assign n18737 =  ( n18037 ) ? ( bv_8_60_n93 ) : ( n18736 ) ;
assign n18738 =  ( n18035 ) ? ( bv_8_21_n89 ) : ( n18737 ) ;
assign n18739 =  ( n18033 ) ? ( bv_8_201_n85 ) : ( n18738 ) ;
assign n18740 =  ( n18031 ) ? ( bv_8_135_n81 ) : ( n18739 ) ;
assign n18741 =  ( n18029 ) ? ( bv_8_170_n77 ) : ( n18740 ) ;
assign n18742 =  ( n18027 ) ? ( bv_8_80_n73 ) : ( n18741 ) ;
assign n18743 =  ( n18025 ) ? ( bv_8_165_n69 ) : ( n18742 ) ;
assign n18744 =  ( n18023 ) ? ( bv_8_3_n65 ) : ( n18743 ) ;
assign n18745 =  ( n18021 ) ? ( bv_8_89_n61 ) : ( n18744 ) ;
assign n18746 =  ( n18019 ) ? ( bv_8_9_n57 ) : ( n18745 ) ;
assign n18747 =  ( n18017 ) ? ( bv_8_26_n53 ) : ( n18746 ) ;
assign n18748 =  ( n18015 ) ? ( bv_8_101_n49 ) : ( n18747 ) ;
assign n18749 =  ( n18013 ) ? ( bv_8_215_n45 ) : ( n18748 ) ;
assign n18750 =  ( n18011 ) ? ( bv_8_132_n41 ) : ( n18749 ) ;
assign n18751 =  ( n18009 ) ? ( bv_8_208_n37 ) : ( n18750 ) ;
assign n18752 =  ( n18007 ) ? ( bv_8_130_n33 ) : ( n18751 ) ;
assign n18753 =  ( n18005 ) ? ( bv_8_41_n29 ) : ( n18752 ) ;
assign n18754 =  ( n18003 ) ? ( bv_8_90_n25 ) : ( n18753 ) ;
assign n18755 =  ( n18001 ) ? ( bv_8_30_n21 ) : ( n18754 ) ;
assign n18756 =  ( n17999 ) ? ( bv_8_123_n17 ) : ( n18755 ) ;
assign n18757 =  ( n17997 ) ? ( bv_8_168_n13 ) : ( n18756 ) ;
assign n18758 =  ( n17995 ) ? ( bv_8_109_n9 ) : ( n18757 ) ;
assign n18759 =  ( n17993 ) ? ( bv_8_44_n5 ) : ( n18758 ) ;
assign n18760 =  ( n17991 ) ^ ( n18759 )  ;
assign n18761 =  ( n18760 ) ^ ( n17985 )  ;
assign n18762 =  ( n18761 ) ^ ( n15674 )  ;
assign n18763 = key[47:40] ;
assign n18764 =  ( n18762 ) ^ ( n18763 )  ;
assign n18765 =  { ( n17990 ) , ( n18764 ) }  ;
assign n18766 =  ( n13368 ) ^ ( n18759 )  ;
assign n18767 =  ( n18766 ) ^ ( n17985 )  ;
assign n18768 =  ( n18767 ) ^ ( n14905 )  ;
assign n18769 =  ( n18768 ) ^ ( n15674 )  ;
assign n18770 = key[39:32] ;
assign n18771 =  ( n18769 ) ^ ( n18770 )  ;
assign n18772 =  { ( n18765 ) , ( n18771 ) }  ;
assign n18773 = state_in[119:112] ;
assign n18774 =  ( n18773 ) == ( bv_8_255_n3 )  ;
assign n18775 = state_in[119:112] ;
assign n18776 =  ( n18775 ) == ( bv_8_254_n7 )  ;
assign n18777 = state_in[119:112] ;
assign n18778 =  ( n18777 ) == ( bv_8_253_n11 )  ;
assign n18779 = state_in[119:112] ;
assign n18780 =  ( n18779 ) == ( bv_8_252_n15 )  ;
assign n18781 = state_in[119:112] ;
assign n18782 =  ( n18781 ) == ( bv_8_251_n19 )  ;
assign n18783 = state_in[119:112] ;
assign n18784 =  ( n18783 ) == ( bv_8_250_n23 )  ;
assign n18785 = state_in[119:112] ;
assign n18786 =  ( n18785 ) == ( bv_8_249_n27 )  ;
assign n18787 = state_in[119:112] ;
assign n18788 =  ( n18787 ) == ( bv_8_248_n31 )  ;
assign n18789 = state_in[119:112] ;
assign n18790 =  ( n18789 ) == ( bv_8_247_n35 )  ;
assign n18791 = state_in[119:112] ;
assign n18792 =  ( n18791 ) == ( bv_8_246_n39 )  ;
assign n18793 = state_in[119:112] ;
assign n18794 =  ( n18793 ) == ( bv_8_245_n43 )  ;
assign n18795 = state_in[119:112] ;
assign n18796 =  ( n18795 ) == ( bv_8_244_n47 )  ;
assign n18797 = state_in[119:112] ;
assign n18798 =  ( n18797 ) == ( bv_8_243_n51 )  ;
assign n18799 = state_in[119:112] ;
assign n18800 =  ( n18799 ) == ( bv_8_242_n55 )  ;
assign n18801 = state_in[119:112] ;
assign n18802 =  ( n18801 ) == ( bv_8_241_n59 )  ;
assign n18803 = state_in[119:112] ;
assign n18804 =  ( n18803 ) == ( bv_8_240_n63 )  ;
assign n18805 = state_in[119:112] ;
assign n18806 =  ( n18805 ) == ( bv_8_239_n67 )  ;
assign n18807 = state_in[119:112] ;
assign n18808 =  ( n18807 ) == ( bv_8_238_n71 )  ;
assign n18809 = state_in[119:112] ;
assign n18810 =  ( n18809 ) == ( bv_8_237_n75 )  ;
assign n18811 = state_in[119:112] ;
assign n18812 =  ( n18811 ) == ( bv_8_236_n79 )  ;
assign n18813 = state_in[119:112] ;
assign n18814 =  ( n18813 ) == ( bv_8_235_n83 )  ;
assign n18815 = state_in[119:112] ;
assign n18816 =  ( n18815 ) == ( bv_8_234_n87 )  ;
assign n18817 = state_in[119:112] ;
assign n18818 =  ( n18817 ) == ( bv_8_233_n91 )  ;
assign n18819 = state_in[119:112] ;
assign n18820 =  ( n18819 ) == ( bv_8_232_n95 )  ;
assign n18821 = state_in[119:112] ;
assign n18822 =  ( n18821 ) == ( bv_8_231_n99 )  ;
assign n18823 = state_in[119:112] ;
assign n18824 =  ( n18823 ) == ( bv_8_230_n103 )  ;
assign n18825 = state_in[119:112] ;
assign n18826 =  ( n18825 ) == ( bv_8_229_n107 )  ;
assign n18827 = state_in[119:112] ;
assign n18828 =  ( n18827 ) == ( bv_8_228_n111 )  ;
assign n18829 = state_in[119:112] ;
assign n18830 =  ( n18829 ) == ( bv_8_227_n115 )  ;
assign n18831 = state_in[119:112] ;
assign n18832 =  ( n18831 ) == ( bv_8_226_n119 )  ;
assign n18833 = state_in[119:112] ;
assign n18834 =  ( n18833 ) == ( bv_8_225_n123 )  ;
assign n18835 = state_in[119:112] ;
assign n18836 =  ( n18835 ) == ( bv_8_224_n126 )  ;
assign n18837 = state_in[119:112] ;
assign n18838 =  ( n18837 ) == ( bv_8_223_n130 )  ;
assign n18839 = state_in[119:112] ;
assign n18840 =  ( n18839 ) == ( bv_8_222_n134 )  ;
assign n18841 = state_in[119:112] ;
assign n18842 =  ( n18841 ) == ( bv_8_221_n138 )  ;
assign n18843 = state_in[119:112] ;
assign n18844 =  ( n18843 ) == ( bv_8_220_n142 )  ;
assign n18845 = state_in[119:112] ;
assign n18846 =  ( n18845 ) == ( bv_8_219_n146 )  ;
assign n18847 = state_in[119:112] ;
assign n18848 =  ( n18847 ) == ( bv_8_218_n150 )  ;
assign n18849 = state_in[119:112] ;
assign n18850 =  ( n18849 ) == ( bv_8_217_n128 )  ;
assign n18851 = state_in[119:112] ;
assign n18852 =  ( n18851 ) == ( bv_8_216_n157 )  ;
assign n18853 = state_in[119:112] ;
assign n18854 =  ( n18853 ) == ( bv_8_215_n45 )  ;
assign n18855 = state_in[119:112] ;
assign n18856 =  ( n18855 ) == ( bv_8_214_n164 )  ;
assign n18857 = state_in[119:112] ;
assign n18858 =  ( n18857 ) == ( bv_8_213_n167 )  ;
assign n18859 = state_in[119:112] ;
assign n18860 =  ( n18859 ) == ( bv_8_212_n171 )  ;
assign n18861 = state_in[119:112] ;
assign n18862 =  ( n18861 ) == ( bv_8_211_n175 )  ;
assign n18863 = state_in[119:112] ;
assign n18864 =  ( n18863 ) == ( bv_8_210_n113 )  ;
assign n18865 = state_in[119:112] ;
assign n18866 =  ( n18865 ) == ( bv_8_209_n182 )  ;
assign n18867 = state_in[119:112] ;
assign n18868 =  ( n18867 ) == ( bv_8_208_n37 )  ;
assign n18869 = state_in[119:112] ;
assign n18870 =  ( n18869 ) == ( bv_8_207_n188 )  ;
assign n18871 = state_in[119:112] ;
assign n18872 =  ( n18871 ) == ( bv_8_206_n192 )  ;
assign n18873 = state_in[119:112] ;
assign n18874 =  ( n18873 ) == ( bv_8_205_n196 )  ;
assign n18875 = state_in[119:112] ;
assign n18876 =  ( n18875 ) == ( bv_8_204_n177 )  ;
assign n18877 = state_in[119:112] ;
assign n18878 =  ( n18877 ) == ( bv_8_203_n203 )  ;
assign n18879 = state_in[119:112] ;
assign n18880 =  ( n18879 ) == ( bv_8_202_n207 )  ;
assign n18881 = state_in[119:112] ;
assign n18882 =  ( n18881 ) == ( bv_8_201_n85 )  ;
assign n18883 = state_in[119:112] ;
assign n18884 =  ( n18883 ) == ( bv_8_200_n213 )  ;
assign n18885 = state_in[119:112] ;
assign n18886 =  ( n18885 ) == ( bv_8_199_n216 )  ;
assign n18887 = state_in[119:112] ;
assign n18888 =  ( n18887 ) == ( bv_8_198_n220 )  ;
assign n18889 = state_in[119:112] ;
assign n18890 =  ( n18889 ) == ( bv_8_197_n224 )  ;
assign n18891 = state_in[119:112] ;
assign n18892 =  ( n18891 ) == ( bv_8_196_n228 )  ;
assign n18893 = state_in[119:112] ;
assign n18894 =  ( n18893 ) == ( bv_8_195_n232 )  ;
assign n18895 = state_in[119:112] ;
assign n18896 =  ( n18895 ) == ( bv_8_194_n159 )  ;
assign n18897 = state_in[119:112] ;
assign n18898 =  ( n18897 ) == ( bv_8_193_n239 )  ;
assign n18899 = state_in[119:112] ;
assign n18900 =  ( n18899 ) == ( bv_8_192_n242 )  ;
assign n18901 = state_in[119:112] ;
assign n18902 =  ( n18901 ) == ( bv_8_191_n246 )  ;
assign n18903 = state_in[119:112] ;
assign n18904 =  ( n18903 ) == ( bv_8_190_n250 )  ;
assign n18905 = state_in[119:112] ;
assign n18906 =  ( n18905 ) == ( bv_8_189_n254 )  ;
assign n18907 = state_in[119:112] ;
assign n18908 =  ( n18907 ) == ( bv_8_188_n257 )  ;
assign n18909 = state_in[119:112] ;
assign n18910 =  ( n18909 ) == ( bv_8_187_n260 )  ;
assign n18911 = state_in[119:112] ;
assign n18912 =  ( n18911 ) == ( bv_8_186_n263 )  ;
assign n18913 = state_in[119:112] ;
assign n18914 =  ( n18913 ) == ( bv_8_185_n266 )  ;
assign n18915 = state_in[119:112] ;
assign n18916 =  ( n18915 ) == ( bv_8_184_n270 )  ;
assign n18917 = state_in[119:112] ;
assign n18918 =  ( n18917 ) == ( bv_8_183_n273 )  ;
assign n18919 = state_in[119:112] ;
assign n18920 =  ( n18919 ) == ( bv_8_182_n277 )  ;
assign n18921 = state_in[119:112] ;
assign n18922 =  ( n18921 ) == ( bv_8_181_n281 )  ;
assign n18923 = state_in[119:112] ;
assign n18924 =  ( n18923 ) == ( bv_8_180_n285 )  ;
assign n18925 = state_in[119:112] ;
assign n18926 =  ( n18925 ) == ( bv_8_179_n289 )  ;
assign n18927 = state_in[119:112] ;
assign n18928 =  ( n18927 ) == ( bv_8_178_n292 )  ;
assign n18929 = state_in[119:112] ;
assign n18930 =  ( n18929 ) == ( bv_8_177_n283 )  ;
assign n18931 = state_in[119:112] ;
assign n18932 =  ( n18931 ) == ( bv_8_176_n299 )  ;
assign n18933 = state_in[119:112] ;
assign n18934 =  ( n18933 ) == ( bv_8_175_n302 )  ;
assign n18935 = state_in[119:112] ;
assign n18936 =  ( n18935 ) == ( bv_8_174_n152 )  ;
assign n18937 = state_in[119:112] ;
assign n18938 =  ( n18937 ) == ( bv_8_173_n307 )  ;
assign n18939 = state_in[119:112] ;
assign n18940 =  ( n18939 ) == ( bv_8_172_n268 )  ;
assign n18941 = state_in[119:112] ;
assign n18942 =  ( n18941 ) == ( bv_8_171_n314 )  ;
assign n18943 = state_in[119:112] ;
assign n18944 =  ( n18943 ) == ( bv_8_170_n77 )  ;
assign n18945 = state_in[119:112] ;
assign n18946 =  ( n18945 ) == ( bv_8_169_n109 )  ;
assign n18947 = state_in[119:112] ;
assign n18948 =  ( n18947 ) == ( bv_8_168_n13 )  ;
assign n18949 = state_in[119:112] ;
assign n18950 =  ( n18949 ) == ( bv_8_167_n325 )  ;
assign n18951 = state_in[119:112] ;
assign n18952 =  ( n18951 ) == ( bv_8_166_n328 )  ;
assign n18953 = state_in[119:112] ;
assign n18954 =  ( n18953 ) == ( bv_8_165_n69 )  ;
assign n18955 = state_in[119:112] ;
assign n18956 =  ( n18955 ) == ( bv_8_164_n335 )  ;
assign n18957 = state_in[119:112] ;
assign n18958 =  ( n18957 ) == ( bv_8_163_n339 )  ;
assign n18959 = state_in[119:112] ;
assign n18960 =  ( n18959 ) == ( bv_8_162_n343 )  ;
assign n18961 = state_in[119:112] ;
assign n18962 =  ( n18961 ) == ( bv_8_161_n211 )  ;
assign n18963 = state_in[119:112] ;
assign n18964 =  ( n18963 ) == ( bv_8_160_n350 )  ;
assign n18965 = state_in[119:112] ;
assign n18966 =  ( n18965 ) == ( bv_8_159_n323 )  ;
assign n18967 = state_in[119:112] ;
assign n18968 =  ( n18967 ) == ( bv_8_158_n355 )  ;
assign n18969 = state_in[119:112] ;
assign n18970 =  ( n18969 ) == ( bv_8_157_n359 )  ;
assign n18971 = state_in[119:112] ;
assign n18972 =  ( n18971 ) == ( bv_8_156_n279 )  ;
assign n18973 = state_in[119:112] ;
assign n18974 =  ( n18973 ) == ( bv_8_155_n364 )  ;
assign n18975 = state_in[119:112] ;
assign n18976 =  ( n18975 ) == ( bv_8_154_n368 )  ;
assign n18977 = state_in[119:112] ;
assign n18978 =  ( n18977 ) == ( bv_8_153_n140 )  ;
assign n18979 = state_in[119:112] ;
assign n18980 =  ( n18979 ) == ( bv_8_152_n374 )  ;
assign n18981 = state_in[119:112] ;
assign n18982 =  ( n18981 ) == ( bv_8_151_n218 )  ;
assign n18983 = state_in[119:112] ;
assign n18984 =  ( n18983 ) == ( bv_8_150_n201 )  ;
assign n18985 = state_in[119:112] ;
assign n18986 =  ( n18985 ) == ( bv_8_149_n384 )  ;
assign n18987 = state_in[119:112] ;
assign n18988 =  ( n18987 ) == ( bv_8_148_n388 )  ;
assign n18989 = state_in[119:112] ;
assign n18990 =  ( n18989 ) == ( bv_8_147_n392 )  ;
assign n18991 = state_in[119:112] ;
assign n18992 =  ( n18991 ) == ( bv_8_146_n337 )  ;
assign n18993 = state_in[119:112] ;
assign n18994 =  ( n18993 ) == ( bv_8_145_n397 )  ;
assign n18995 = state_in[119:112] ;
assign n18996 =  ( n18995 ) == ( bv_8_144_n173 )  ;
assign n18997 = state_in[119:112] ;
assign n18998 =  ( n18997 ) == ( bv_8_143_n403 )  ;
assign n18999 = state_in[119:112] ;
assign n19000 =  ( n18999 ) == ( bv_8_142_n406 )  ;
assign n19001 = state_in[119:112] ;
assign n19002 =  ( n19001 ) == ( bv_8_141_n410 )  ;
assign n19003 = state_in[119:112] ;
assign n19004 =  ( n19003 ) == ( bv_8_140_n376 )  ;
assign n19005 = state_in[119:112] ;
assign n19006 =  ( n19005 ) == ( bv_8_139_n297 )  ;
assign n19007 = state_in[119:112] ;
assign n19008 =  ( n19007 ) == ( bv_8_138_n418 )  ;
assign n19009 = state_in[119:112] ;
assign n19010 =  ( n19009 ) == ( bv_8_137_n421 )  ;
assign n19011 = state_in[119:112] ;
assign n19012 =  ( n19011 ) == ( bv_8_136_n425 )  ;
assign n19013 = state_in[119:112] ;
assign n19014 =  ( n19013 ) == ( bv_8_135_n81 )  ;
assign n19015 = state_in[119:112] ;
assign n19016 =  ( n19015 ) == ( bv_8_134_n431 )  ;
assign n19017 = state_in[119:112] ;
assign n19018 =  ( n19017 ) == ( bv_8_133_n434 )  ;
assign n19019 = state_in[119:112] ;
assign n19020 =  ( n19019 ) == ( bv_8_132_n41 )  ;
assign n19021 = state_in[119:112] ;
assign n19022 =  ( n19021 ) == ( bv_8_131_n440 )  ;
assign n19023 = state_in[119:112] ;
assign n19024 =  ( n19023 ) == ( bv_8_130_n33 )  ;
assign n19025 = state_in[119:112] ;
assign n19026 =  ( n19025 ) == ( bv_8_129_n446 )  ;
assign n19027 = state_in[119:112] ;
assign n19028 =  ( n19027 ) == ( bv_8_128_n450 )  ;
assign n19029 = state_in[119:112] ;
assign n19030 =  ( n19029 ) == ( bv_8_127_n453 )  ;
assign n19031 = state_in[119:112] ;
assign n19032 =  ( n19031 ) == ( bv_8_126_n456 )  ;
assign n19033 = state_in[119:112] ;
assign n19034 =  ( n19033 ) == ( bv_8_125_n459 )  ;
assign n19035 = state_in[119:112] ;
assign n19036 =  ( n19035 ) == ( bv_8_124_n184 )  ;
assign n19037 = state_in[119:112] ;
assign n19038 =  ( n19037 ) == ( bv_8_123_n17 )  ;
assign n19039 = state_in[119:112] ;
assign n19040 =  ( n19039 ) == ( bv_8_122_n416 )  ;
assign n19041 = state_in[119:112] ;
assign n19042 =  ( n19041 ) == ( bv_8_121_n470 )  ;
assign n19043 = state_in[119:112] ;
assign n19044 =  ( n19043 ) == ( bv_8_120_n474 )  ;
assign n19045 = state_in[119:112] ;
assign n19046 =  ( n19045 ) == ( bv_8_119_n472 )  ;
assign n19047 = state_in[119:112] ;
assign n19048 =  ( n19047 ) == ( bv_8_118_n480 )  ;
assign n19049 = state_in[119:112] ;
assign n19050 =  ( n19049 ) == ( bv_8_117_n484 )  ;
assign n19051 = state_in[119:112] ;
assign n19052 =  ( n19051 ) == ( bv_8_116_n345 )  ;
assign n19053 = state_in[119:112] ;
assign n19054 =  ( n19053 ) == ( bv_8_115_n222 )  ;
assign n19055 = state_in[119:112] ;
assign n19056 =  ( n19055 ) == ( bv_8_114_n494 )  ;
assign n19057 = state_in[119:112] ;
assign n19058 =  ( n19057 ) == ( bv_8_113_n180 )  ;
assign n19059 = state_in[119:112] ;
assign n19060 =  ( n19059 ) == ( bv_8_112_n482 )  ;
assign n19061 = state_in[119:112] ;
assign n19062 =  ( n19061 ) == ( bv_8_111_n244 )  ;
assign n19063 = state_in[119:112] ;
assign n19064 =  ( n19063 ) == ( bv_8_110_n294 )  ;
assign n19065 = state_in[119:112] ;
assign n19066 =  ( n19065 ) == ( bv_8_109_n9 )  ;
assign n19067 = state_in[119:112] ;
assign n19068 =  ( n19067 ) == ( bv_8_108_n510 )  ;
assign n19069 = state_in[119:112] ;
assign n19070 =  ( n19069 ) == ( bv_8_107_n370 )  ;
assign n19071 = state_in[119:112] ;
assign n19072 =  ( n19071 ) == ( bv_8_106_n155 )  ;
assign n19073 = state_in[119:112] ;
assign n19074 =  ( n19073 ) == ( bv_8_105_n148 )  ;
assign n19075 = state_in[119:112] ;
assign n19076 =  ( n19075 ) == ( bv_8_104_n520 )  ;
assign n19077 = state_in[119:112] ;
assign n19078 =  ( n19077 ) == ( bv_8_103_n523 )  ;
assign n19079 = state_in[119:112] ;
assign n19080 =  ( n19079 ) == ( bv_8_102_n527 )  ;
assign n19081 = state_in[119:112] ;
assign n19082 =  ( n19081 ) == ( bv_8_101_n49 )  ;
assign n19083 = state_in[119:112] ;
assign n19084 =  ( n19083 ) == ( bv_8_100_n348 )  ;
assign n19085 = state_in[119:112] ;
assign n19086 =  ( n19085 ) == ( bv_8_99_n476 )  ;
assign n19087 = state_in[119:112] ;
assign n19088 =  ( n19087 ) == ( bv_8_98_n536 )  ;
assign n19089 = state_in[119:112] ;
assign n19090 =  ( n19089 ) == ( bv_8_97_n198 )  ;
assign n19091 = state_in[119:112] ;
assign n19092 =  ( n19091 ) == ( bv_8_96_n542 )  ;
assign n19093 = state_in[119:112] ;
assign n19094 =  ( n19093 ) == ( bv_8_95_n545 )  ;
assign n19095 = state_in[119:112] ;
assign n19096 =  ( n19095 ) == ( bv_8_94_n548 )  ;
assign n19097 = state_in[119:112] ;
assign n19098 =  ( n19097 ) == ( bv_8_93_n498 )  ;
assign n19099 = state_in[119:112] ;
assign n19100 =  ( n19099 ) == ( bv_8_92_n234 )  ;
assign n19101 = state_in[119:112] ;
assign n19102 =  ( n19101 ) == ( bv_8_91_n555 )  ;
assign n19103 = state_in[119:112] ;
assign n19104 =  ( n19103 ) == ( bv_8_90_n25 )  ;
assign n19105 = state_in[119:112] ;
assign n19106 =  ( n19105 ) == ( bv_8_89_n61 )  ;
assign n19107 = state_in[119:112] ;
assign n19108 =  ( n19107 ) == ( bv_8_88_n562 )  ;
assign n19109 = state_in[119:112] ;
assign n19110 =  ( n19109 ) == ( bv_8_87_n226 )  ;
assign n19111 = state_in[119:112] ;
assign n19112 =  ( n19111 ) == ( bv_8_86_n567 )  ;
assign n19113 = state_in[119:112] ;
assign n19114 =  ( n19113 ) == ( bv_8_85_n423 )  ;
assign n19115 = state_in[119:112] ;
assign n19116 =  ( n19115 ) == ( bv_8_84_n386 )  ;
assign n19117 = state_in[119:112] ;
assign n19118 =  ( n19117 ) == ( bv_8_83_n575 )  ;
assign n19119 = state_in[119:112] ;
assign n19120 =  ( n19119 ) == ( bv_8_82_n578 )  ;
assign n19121 = state_in[119:112] ;
assign n19122 =  ( n19121 ) == ( bv_8_81_n582 )  ;
assign n19123 = state_in[119:112] ;
assign n19124 =  ( n19123 ) == ( bv_8_80_n73 )  ;
assign n19125 = state_in[119:112] ;
assign n19126 =  ( n19125 ) == ( bv_8_79_n538 )  ;
assign n19127 = state_in[119:112] ;
assign n19128 =  ( n19127 ) == ( bv_8_78_n590 )  ;
assign n19129 = state_in[119:112] ;
assign n19130 =  ( n19129 ) == ( bv_8_77_n593 )  ;
assign n19131 = state_in[119:112] ;
assign n19132 =  ( n19131 ) == ( bv_8_76_n596 )  ;
assign n19133 = state_in[119:112] ;
assign n19134 =  ( n19133 ) == ( bv_8_75_n503 )  ;
assign n19135 = state_in[119:112] ;
assign n19136 =  ( n19135 ) == ( bv_8_74_n237 )  ;
assign n19137 = state_in[119:112] ;
assign n19138 =  ( n19137 ) == ( bv_8_73_n275 )  ;
assign n19139 = state_in[119:112] ;
assign n19140 =  ( n19139 ) == ( bv_8_72_n330 )  ;
assign n19141 = state_in[119:112] ;
assign n19142 =  ( n19141 ) == ( bv_8_71_n252 )  ;
assign n19143 = state_in[119:112] ;
assign n19144 =  ( n19143 ) == ( bv_8_70_n609 )  ;
assign n19145 = state_in[119:112] ;
assign n19146 =  ( n19145 ) == ( bv_8_69_n612 )  ;
assign n19147 = state_in[119:112] ;
assign n19148 =  ( n19147 ) == ( bv_8_68_n390 )  ;
assign n19149 = state_in[119:112] ;
assign n19150 =  ( n19149 ) == ( bv_8_67_n318 )  ;
assign n19151 = state_in[119:112] ;
assign n19152 =  ( n19151 ) == ( bv_8_66_n466 )  ;
assign n19153 = state_in[119:112] ;
assign n19154 =  ( n19153 ) == ( bv_8_65_n623 )  ;
assign n19155 = state_in[119:112] ;
assign n19156 =  ( n19155 ) == ( bv_8_64_n573 )  ;
assign n19157 = state_in[119:112] ;
assign n19158 =  ( n19157 ) == ( bv_8_63_n489 )  ;
assign n19159 = state_in[119:112] ;
assign n19160 =  ( n19159 ) == ( bv_8_62_n205 )  ;
assign n19161 = state_in[119:112] ;
assign n19162 =  ( n19161 ) == ( bv_8_61_n634 )  ;
assign n19163 = state_in[119:112] ;
assign n19164 =  ( n19163 ) == ( bv_8_60_n93 )  ;
assign n19165 = state_in[119:112] ;
assign n19166 =  ( n19165 ) == ( bv_8_59_n382 )  ;
assign n19167 = state_in[119:112] ;
assign n19168 =  ( n19167 ) == ( bv_8_58_n136 )  ;
assign n19169 = state_in[119:112] ;
assign n19170 =  ( n19169 ) == ( bv_8_57_n312 )  ;
assign n19171 = state_in[119:112] ;
assign n19172 =  ( n19171 ) == ( bv_8_56_n230 )  ;
assign n19173 = state_in[119:112] ;
assign n19174 =  ( n19173 ) == ( bv_8_55_n650 )  ;
assign n19175 = state_in[119:112] ;
assign n19176 =  ( n19175 ) == ( bv_8_54_n616 )  ;
assign n19177 = state_in[119:112] ;
assign n19178 =  ( n19177 ) == ( bv_8_53_n436 )  ;
assign n19179 = state_in[119:112] ;
assign n19180 =  ( n19179 ) == ( bv_8_52_n619 )  ;
assign n19181 = state_in[119:112] ;
assign n19182 =  ( n19181 ) == ( bv_8_51_n101 )  ;
assign n19183 = state_in[119:112] ;
assign n19184 =  ( n19183 ) == ( bv_8_50_n408 )  ;
assign n19185 = state_in[119:112] ;
assign n19186 =  ( n19185 ) == ( bv_8_49_n309 )  ;
assign n19187 = state_in[119:112] ;
assign n19188 =  ( n19187 ) == ( bv_8_48_n660 )  ;
assign n19189 = state_in[119:112] ;
assign n19190 =  ( n19189 ) == ( bv_8_47_n652 )  ;
assign n19191 = state_in[119:112] ;
assign n19192 =  ( n19191 ) == ( bv_8_46_n429 )  ;
assign n19193 = state_in[119:112] ;
assign n19194 =  ( n19193 ) == ( bv_8_45_n97 )  ;
assign n19195 = state_in[119:112] ;
assign n19196 =  ( n19195 ) == ( bv_8_44_n5 )  ;
assign n19197 = state_in[119:112] ;
assign n19198 =  ( n19197 ) == ( bv_8_43_n121 )  ;
assign n19199 = state_in[119:112] ;
assign n19200 =  ( n19199 ) == ( bv_8_42_n672 )  ;
assign n19201 = state_in[119:112] ;
assign n19202 =  ( n19201 ) == ( bv_8_41_n29 )  ;
assign n19203 = state_in[119:112] ;
assign n19204 =  ( n19203 ) == ( bv_8_40_n366 )  ;
assign n19205 = state_in[119:112] ;
assign n19206 =  ( n19205 ) == ( bv_8_39_n132 )  ;
assign n19207 = state_in[119:112] ;
assign n19208 =  ( n19207 ) == ( bv_8_38_n444 )  ;
assign n19209 = state_in[119:112] ;
assign n19210 =  ( n19209 ) == ( bv_8_37_n506 )  ;
assign n19211 = state_in[119:112] ;
assign n19212 =  ( n19211 ) == ( bv_8_36_n645 )  ;
assign n19213 = state_in[119:112] ;
assign n19214 =  ( n19213 ) == ( bv_8_35_n696 )  ;
assign n19215 = state_in[119:112] ;
assign n19216 =  ( n19215 ) == ( bv_8_34_n117 )  ;
assign n19217 = state_in[119:112] ;
assign n19218 =  ( n19217 ) == ( bv_8_33_n486 )  ;
assign n19219 = state_in[119:112] ;
assign n19220 =  ( n19219 ) == ( bv_8_32_n463 )  ;
assign n19221 = state_in[119:112] ;
assign n19222 =  ( n19221 ) == ( bv_8_31_n705 )  ;
assign n19223 = state_in[119:112] ;
assign n19224 =  ( n19223 ) == ( bv_8_30_n21 )  ;
assign n19225 = state_in[119:112] ;
assign n19226 =  ( n19225 ) == ( bv_8_29_n625 )  ;
assign n19227 = state_in[119:112] ;
assign n19228 =  ( n19227 ) == ( bv_8_28_n162 )  ;
assign n19229 = state_in[119:112] ;
assign n19230 =  ( n19229 ) == ( bv_8_27_n642 )  ;
assign n19231 = state_in[119:112] ;
assign n19232 =  ( n19231 ) == ( bv_8_26_n53 )  ;
assign n19233 = state_in[119:112] ;
assign n19234 =  ( n19233 ) == ( bv_8_25_n399 )  ;
assign n19235 = state_in[119:112] ;
assign n19236 =  ( n19235 ) == ( bv_8_24_n448 )  ;
assign n19237 = state_in[119:112] ;
assign n19238 =  ( n19237 ) == ( bv_8_23_n144 )  ;
assign n19239 = state_in[119:112] ;
assign n19240 =  ( n19239 ) == ( bv_8_22_n357 )  ;
assign n19241 = state_in[119:112] ;
assign n19242 =  ( n19241 ) == ( bv_8_21_n89 )  ;
assign n19243 = state_in[119:112] ;
assign n19244 =  ( n19243 ) == ( bv_8_20_n341 )  ;
assign n19245 = state_in[119:112] ;
assign n19246 =  ( n19245 ) == ( bv_8_19_n588 )  ;
assign n19247 = state_in[119:112] ;
assign n19248 =  ( n19247 ) == ( bv_8_18_n628 )  ;
assign n19249 = state_in[119:112] ;
assign n19250 =  ( n19249 ) == ( bv_8_17_n525 )  ;
assign n19251 = state_in[119:112] ;
assign n19252 =  ( n19251 ) == ( bv_8_16_n248 )  ;
assign n19253 = state_in[119:112] ;
assign n19254 =  ( n19253 ) == ( bv_8_15_n190 )  ;
assign n19255 = state_in[119:112] ;
assign n19256 =  ( n19255 ) == ( bv_8_14_n648 )  ;
assign n19257 = state_in[119:112] ;
assign n19258 =  ( n19257 ) == ( bv_8_13_n194 )  ;
assign n19259 = state_in[119:112] ;
assign n19260 =  ( n19259 ) == ( bv_8_12_n333 )  ;
assign n19261 = state_in[119:112] ;
assign n19262 =  ( n19261 ) == ( bv_8_11_n379 )  ;
assign n19263 = state_in[119:112] ;
assign n19264 =  ( n19263 ) == ( bv_8_10_n655 )  ;
assign n19265 = state_in[119:112] ;
assign n19266 =  ( n19265 ) == ( bv_8_9_n57 )  ;
assign n19267 = state_in[119:112] ;
assign n19268 =  ( n19267 ) == ( bv_8_8_n669 )  ;
assign n19269 = state_in[119:112] ;
assign n19270 =  ( n19269 ) == ( bv_8_7_n105 )  ;
assign n19271 = state_in[119:112] ;
assign n19272 =  ( n19271 ) == ( bv_8_6_n169 )  ;
assign n19273 = state_in[119:112] ;
assign n19274 =  ( n19273 ) == ( bv_8_5_n492 )  ;
assign n19275 = state_in[119:112] ;
assign n19276 =  ( n19275 ) == ( bv_8_4_n516 )  ;
assign n19277 = state_in[119:112] ;
assign n19278 =  ( n19277 ) == ( bv_8_3_n65 )  ;
assign n19279 = state_in[119:112] ;
assign n19280 =  ( n19279 ) == ( bv_8_2_n751 )  ;
assign n19281 = state_in[119:112] ;
assign n19282 =  ( n19281 ) == ( bv_8_1_n287 )  ;
assign n19283 = state_in[119:112] ;
assign n19284 =  ( n19283 ) == ( bv_8_0_n580 )  ;
assign n19285 =  ( n19284 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n19286 =  ( n19282 ) ? ( bv_8_124_n184 ) : ( n19285 ) ;
assign n19287 =  ( n19280 ) ? ( bv_8_119_n472 ) : ( n19286 ) ;
assign n19288 =  ( n19278 ) ? ( bv_8_123_n17 ) : ( n19287 ) ;
assign n19289 =  ( n19276 ) ? ( bv_8_242_n55 ) : ( n19288 ) ;
assign n19290 =  ( n19274 ) ? ( bv_8_107_n370 ) : ( n19289 ) ;
assign n19291 =  ( n19272 ) ? ( bv_8_111_n244 ) : ( n19290 ) ;
assign n19292 =  ( n19270 ) ? ( bv_8_197_n224 ) : ( n19291 ) ;
assign n19293 =  ( n19268 ) ? ( bv_8_48_n660 ) : ( n19292 ) ;
assign n19294 =  ( n19266 ) ? ( bv_8_1_n287 ) : ( n19293 ) ;
assign n19295 =  ( n19264 ) ? ( bv_8_103_n523 ) : ( n19294 ) ;
assign n19296 =  ( n19262 ) ? ( bv_8_43_n121 ) : ( n19295 ) ;
assign n19297 =  ( n19260 ) ? ( bv_8_254_n7 ) : ( n19296 ) ;
assign n19298 =  ( n19258 ) ? ( bv_8_215_n45 ) : ( n19297 ) ;
assign n19299 =  ( n19256 ) ? ( bv_8_171_n314 ) : ( n19298 ) ;
assign n19300 =  ( n19254 ) ? ( bv_8_118_n480 ) : ( n19299 ) ;
assign n19301 =  ( n19252 ) ? ( bv_8_202_n207 ) : ( n19300 ) ;
assign n19302 =  ( n19250 ) ? ( bv_8_130_n33 ) : ( n19301 ) ;
assign n19303 =  ( n19248 ) ? ( bv_8_201_n85 ) : ( n19302 ) ;
assign n19304 =  ( n19246 ) ? ( bv_8_125_n459 ) : ( n19303 ) ;
assign n19305 =  ( n19244 ) ? ( bv_8_250_n23 ) : ( n19304 ) ;
assign n19306 =  ( n19242 ) ? ( bv_8_89_n61 ) : ( n19305 ) ;
assign n19307 =  ( n19240 ) ? ( bv_8_71_n252 ) : ( n19306 ) ;
assign n19308 =  ( n19238 ) ? ( bv_8_240_n63 ) : ( n19307 ) ;
assign n19309 =  ( n19236 ) ? ( bv_8_173_n307 ) : ( n19308 ) ;
assign n19310 =  ( n19234 ) ? ( bv_8_212_n171 ) : ( n19309 ) ;
assign n19311 =  ( n19232 ) ? ( bv_8_162_n343 ) : ( n19310 ) ;
assign n19312 =  ( n19230 ) ? ( bv_8_175_n302 ) : ( n19311 ) ;
assign n19313 =  ( n19228 ) ? ( bv_8_156_n279 ) : ( n19312 ) ;
assign n19314 =  ( n19226 ) ? ( bv_8_164_n335 ) : ( n19313 ) ;
assign n19315 =  ( n19224 ) ? ( bv_8_114_n494 ) : ( n19314 ) ;
assign n19316 =  ( n19222 ) ? ( bv_8_192_n242 ) : ( n19315 ) ;
assign n19317 =  ( n19220 ) ? ( bv_8_183_n273 ) : ( n19316 ) ;
assign n19318 =  ( n19218 ) ? ( bv_8_253_n11 ) : ( n19317 ) ;
assign n19319 =  ( n19216 ) ? ( bv_8_147_n392 ) : ( n19318 ) ;
assign n19320 =  ( n19214 ) ? ( bv_8_38_n444 ) : ( n19319 ) ;
assign n19321 =  ( n19212 ) ? ( bv_8_54_n616 ) : ( n19320 ) ;
assign n19322 =  ( n19210 ) ? ( bv_8_63_n489 ) : ( n19321 ) ;
assign n19323 =  ( n19208 ) ? ( bv_8_247_n35 ) : ( n19322 ) ;
assign n19324 =  ( n19206 ) ? ( bv_8_204_n177 ) : ( n19323 ) ;
assign n19325 =  ( n19204 ) ? ( bv_8_52_n619 ) : ( n19324 ) ;
assign n19326 =  ( n19202 ) ? ( bv_8_165_n69 ) : ( n19325 ) ;
assign n19327 =  ( n19200 ) ? ( bv_8_229_n107 ) : ( n19326 ) ;
assign n19328 =  ( n19198 ) ? ( bv_8_241_n59 ) : ( n19327 ) ;
assign n19329 =  ( n19196 ) ? ( bv_8_113_n180 ) : ( n19328 ) ;
assign n19330 =  ( n19194 ) ? ( bv_8_216_n157 ) : ( n19329 ) ;
assign n19331 =  ( n19192 ) ? ( bv_8_49_n309 ) : ( n19330 ) ;
assign n19332 =  ( n19190 ) ? ( bv_8_21_n89 ) : ( n19331 ) ;
assign n19333 =  ( n19188 ) ? ( bv_8_4_n516 ) : ( n19332 ) ;
assign n19334 =  ( n19186 ) ? ( bv_8_199_n216 ) : ( n19333 ) ;
assign n19335 =  ( n19184 ) ? ( bv_8_35_n696 ) : ( n19334 ) ;
assign n19336 =  ( n19182 ) ? ( bv_8_195_n232 ) : ( n19335 ) ;
assign n19337 =  ( n19180 ) ? ( bv_8_24_n448 ) : ( n19336 ) ;
assign n19338 =  ( n19178 ) ? ( bv_8_150_n201 ) : ( n19337 ) ;
assign n19339 =  ( n19176 ) ? ( bv_8_5_n492 ) : ( n19338 ) ;
assign n19340 =  ( n19174 ) ? ( bv_8_154_n368 ) : ( n19339 ) ;
assign n19341 =  ( n19172 ) ? ( bv_8_7_n105 ) : ( n19340 ) ;
assign n19342 =  ( n19170 ) ? ( bv_8_18_n628 ) : ( n19341 ) ;
assign n19343 =  ( n19168 ) ? ( bv_8_128_n450 ) : ( n19342 ) ;
assign n19344 =  ( n19166 ) ? ( bv_8_226_n119 ) : ( n19343 ) ;
assign n19345 =  ( n19164 ) ? ( bv_8_235_n83 ) : ( n19344 ) ;
assign n19346 =  ( n19162 ) ? ( bv_8_39_n132 ) : ( n19345 ) ;
assign n19347 =  ( n19160 ) ? ( bv_8_178_n292 ) : ( n19346 ) ;
assign n19348 =  ( n19158 ) ? ( bv_8_117_n484 ) : ( n19347 ) ;
assign n19349 =  ( n19156 ) ? ( bv_8_9_n57 ) : ( n19348 ) ;
assign n19350 =  ( n19154 ) ? ( bv_8_131_n440 ) : ( n19349 ) ;
assign n19351 =  ( n19152 ) ? ( bv_8_44_n5 ) : ( n19350 ) ;
assign n19352 =  ( n19150 ) ? ( bv_8_26_n53 ) : ( n19351 ) ;
assign n19353 =  ( n19148 ) ? ( bv_8_27_n642 ) : ( n19352 ) ;
assign n19354 =  ( n19146 ) ? ( bv_8_110_n294 ) : ( n19353 ) ;
assign n19355 =  ( n19144 ) ? ( bv_8_90_n25 ) : ( n19354 ) ;
assign n19356 =  ( n19142 ) ? ( bv_8_160_n350 ) : ( n19355 ) ;
assign n19357 =  ( n19140 ) ? ( bv_8_82_n578 ) : ( n19356 ) ;
assign n19358 =  ( n19138 ) ? ( bv_8_59_n382 ) : ( n19357 ) ;
assign n19359 =  ( n19136 ) ? ( bv_8_214_n164 ) : ( n19358 ) ;
assign n19360 =  ( n19134 ) ? ( bv_8_179_n289 ) : ( n19359 ) ;
assign n19361 =  ( n19132 ) ? ( bv_8_41_n29 ) : ( n19360 ) ;
assign n19362 =  ( n19130 ) ? ( bv_8_227_n115 ) : ( n19361 ) ;
assign n19363 =  ( n19128 ) ? ( bv_8_47_n652 ) : ( n19362 ) ;
assign n19364 =  ( n19126 ) ? ( bv_8_132_n41 ) : ( n19363 ) ;
assign n19365 =  ( n19124 ) ? ( bv_8_83_n575 ) : ( n19364 ) ;
assign n19366 =  ( n19122 ) ? ( bv_8_209_n182 ) : ( n19365 ) ;
assign n19367 =  ( n19120 ) ? ( bv_8_0_n580 ) : ( n19366 ) ;
assign n19368 =  ( n19118 ) ? ( bv_8_237_n75 ) : ( n19367 ) ;
assign n19369 =  ( n19116 ) ? ( bv_8_32_n463 ) : ( n19368 ) ;
assign n19370 =  ( n19114 ) ? ( bv_8_252_n15 ) : ( n19369 ) ;
assign n19371 =  ( n19112 ) ? ( bv_8_177_n283 ) : ( n19370 ) ;
assign n19372 =  ( n19110 ) ? ( bv_8_91_n555 ) : ( n19371 ) ;
assign n19373 =  ( n19108 ) ? ( bv_8_106_n155 ) : ( n19372 ) ;
assign n19374 =  ( n19106 ) ? ( bv_8_203_n203 ) : ( n19373 ) ;
assign n19375 =  ( n19104 ) ? ( bv_8_190_n250 ) : ( n19374 ) ;
assign n19376 =  ( n19102 ) ? ( bv_8_57_n312 ) : ( n19375 ) ;
assign n19377 =  ( n19100 ) ? ( bv_8_74_n237 ) : ( n19376 ) ;
assign n19378 =  ( n19098 ) ? ( bv_8_76_n596 ) : ( n19377 ) ;
assign n19379 =  ( n19096 ) ? ( bv_8_88_n562 ) : ( n19378 ) ;
assign n19380 =  ( n19094 ) ? ( bv_8_207_n188 ) : ( n19379 ) ;
assign n19381 =  ( n19092 ) ? ( bv_8_208_n37 ) : ( n19380 ) ;
assign n19382 =  ( n19090 ) ? ( bv_8_239_n67 ) : ( n19381 ) ;
assign n19383 =  ( n19088 ) ? ( bv_8_170_n77 ) : ( n19382 ) ;
assign n19384 =  ( n19086 ) ? ( bv_8_251_n19 ) : ( n19383 ) ;
assign n19385 =  ( n19084 ) ? ( bv_8_67_n318 ) : ( n19384 ) ;
assign n19386 =  ( n19082 ) ? ( bv_8_77_n593 ) : ( n19385 ) ;
assign n19387 =  ( n19080 ) ? ( bv_8_51_n101 ) : ( n19386 ) ;
assign n19388 =  ( n19078 ) ? ( bv_8_133_n434 ) : ( n19387 ) ;
assign n19389 =  ( n19076 ) ? ( bv_8_69_n612 ) : ( n19388 ) ;
assign n19390 =  ( n19074 ) ? ( bv_8_249_n27 ) : ( n19389 ) ;
assign n19391 =  ( n19072 ) ? ( bv_8_2_n751 ) : ( n19390 ) ;
assign n19392 =  ( n19070 ) ? ( bv_8_127_n453 ) : ( n19391 ) ;
assign n19393 =  ( n19068 ) ? ( bv_8_80_n73 ) : ( n19392 ) ;
assign n19394 =  ( n19066 ) ? ( bv_8_60_n93 ) : ( n19393 ) ;
assign n19395 =  ( n19064 ) ? ( bv_8_159_n323 ) : ( n19394 ) ;
assign n19396 =  ( n19062 ) ? ( bv_8_168_n13 ) : ( n19395 ) ;
assign n19397 =  ( n19060 ) ? ( bv_8_81_n582 ) : ( n19396 ) ;
assign n19398 =  ( n19058 ) ? ( bv_8_163_n339 ) : ( n19397 ) ;
assign n19399 =  ( n19056 ) ? ( bv_8_64_n573 ) : ( n19398 ) ;
assign n19400 =  ( n19054 ) ? ( bv_8_143_n403 ) : ( n19399 ) ;
assign n19401 =  ( n19052 ) ? ( bv_8_146_n337 ) : ( n19400 ) ;
assign n19402 =  ( n19050 ) ? ( bv_8_157_n359 ) : ( n19401 ) ;
assign n19403 =  ( n19048 ) ? ( bv_8_56_n230 ) : ( n19402 ) ;
assign n19404 =  ( n19046 ) ? ( bv_8_245_n43 ) : ( n19403 ) ;
assign n19405 =  ( n19044 ) ? ( bv_8_188_n257 ) : ( n19404 ) ;
assign n19406 =  ( n19042 ) ? ( bv_8_182_n277 ) : ( n19405 ) ;
assign n19407 =  ( n19040 ) ? ( bv_8_218_n150 ) : ( n19406 ) ;
assign n19408 =  ( n19038 ) ? ( bv_8_33_n486 ) : ( n19407 ) ;
assign n19409 =  ( n19036 ) ? ( bv_8_16_n248 ) : ( n19408 ) ;
assign n19410 =  ( n19034 ) ? ( bv_8_255_n3 ) : ( n19409 ) ;
assign n19411 =  ( n19032 ) ? ( bv_8_243_n51 ) : ( n19410 ) ;
assign n19412 =  ( n19030 ) ? ( bv_8_210_n113 ) : ( n19411 ) ;
assign n19413 =  ( n19028 ) ? ( bv_8_205_n196 ) : ( n19412 ) ;
assign n19414 =  ( n19026 ) ? ( bv_8_12_n333 ) : ( n19413 ) ;
assign n19415 =  ( n19024 ) ? ( bv_8_19_n588 ) : ( n19414 ) ;
assign n19416 =  ( n19022 ) ? ( bv_8_236_n79 ) : ( n19415 ) ;
assign n19417 =  ( n19020 ) ? ( bv_8_95_n545 ) : ( n19416 ) ;
assign n19418 =  ( n19018 ) ? ( bv_8_151_n218 ) : ( n19417 ) ;
assign n19419 =  ( n19016 ) ? ( bv_8_68_n390 ) : ( n19418 ) ;
assign n19420 =  ( n19014 ) ? ( bv_8_23_n144 ) : ( n19419 ) ;
assign n19421 =  ( n19012 ) ? ( bv_8_196_n228 ) : ( n19420 ) ;
assign n19422 =  ( n19010 ) ? ( bv_8_167_n325 ) : ( n19421 ) ;
assign n19423 =  ( n19008 ) ? ( bv_8_126_n456 ) : ( n19422 ) ;
assign n19424 =  ( n19006 ) ? ( bv_8_61_n634 ) : ( n19423 ) ;
assign n19425 =  ( n19004 ) ? ( bv_8_100_n348 ) : ( n19424 ) ;
assign n19426 =  ( n19002 ) ? ( bv_8_93_n498 ) : ( n19425 ) ;
assign n19427 =  ( n19000 ) ? ( bv_8_25_n399 ) : ( n19426 ) ;
assign n19428 =  ( n18998 ) ? ( bv_8_115_n222 ) : ( n19427 ) ;
assign n19429 =  ( n18996 ) ? ( bv_8_96_n542 ) : ( n19428 ) ;
assign n19430 =  ( n18994 ) ? ( bv_8_129_n446 ) : ( n19429 ) ;
assign n19431 =  ( n18992 ) ? ( bv_8_79_n538 ) : ( n19430 ) ;
assign n19432 =  ( n18990 ) ? ( bv_8_220_n142 ) : ( n19431 ) ;
assign n19433 =  ( n18988 ) ? ( bv_8_34_n117 ) : ( n19432 ) ;
assign n19434 =  ( n18986 ) ? ( bv_8_42_n672 ) : ( n19433 ) ;
assign n19435 =  ( n18984 ) ? ( bv_8_144_n173 ) : ( n19434 ) ;
assign n19436 =  ( n18982 ) ? ( bv_8_136_n425 ) : ( n19435 ) ;
assign n19437 =  ( n18980 ) ? ( bv_8_70_n609 ) : ( n19436 ) ;
assign n19438 =  ( n18978 ) ? ( bv_8_238_n71 ) : ( n19437 ) ;
assign n19439 =  ( n18976 ) ? ( bv_8_184_n270 ) : ( n19438 ) ;
assign n19440 =  ( n18974 ) ? ( bv_8_20_n341 ) : ( n19439 ) ;
assign n19441 =  ( n18972 ) ? ( bv_8_222_n134 ) : ( n19440 ) ;
assign n19442 =  ( n18970 ) ? ( bv_8_94_n548 ) : ( n19441 ) ;
assign n19443 =  ( n18968 ) ? ( bv_8_11_n379 ) : ( n19442 ) ;
assign n19444 =  ( n18966 ) ? ( bv_8_219_n146 ) : ( n19443 ) ;
assign n19445 =  ( n18964 ) ? ( bv_8_224_n126 ) : ( n19444 ) ;
assign n19446 =  ( n18962 ) ? ( bv_8_50_n408 ) : ( n19445 ) ;
assign n19447 =  ( n18960 ) ? ( bv_8_58_n136 ) : ( n19446 ) ;
assign n19448 =  ( n18958 ) ? ( bv_8_10_n655 ) : ( n19447 ) ;
assign n19449 =  ( n18956 ) ? ( bv_8_73_n275 ) : ( n19448 ) ;
assign n19450 =  ( n18954 ) ? ( bv_8_6_n169 ) : ( n19449 ) ;
assign n19451 =  ( n18952 ) ? ( bv_8_36_n645 ) : ( n19450 ) ;
assign n19452 =  ( n18950 ) ? ( bv_8_92_n234 ) : ( n19451 ) ;
assign n19453 =  ( n18948 ) ? ( bv_8_194_n159 ) : ( n19452 ) ;
assign n19454 =  ( n18946 ) ? ( bv_8_211_n175 ) : ( n19453 ) ;
assign n19455 =  ( n18944 ) ? ( bv_8_172_n268 ) : ( n19454 ) ;
assign n19456 =  ( n18942 ) ? ( bv_8_98_n536 ) : ( n19455 ) ;
assign n19457 =  ( n18940 ) ? ( bv_8_145_n397 ) : ( n19456 ) ;
assign n19458 =  ( n18938 ) ? ( bv_8_149_n384 ) : ( n19457 ) ;
assign n19459 =  ( n18936 ) ? ( bv_8_228_n111 ) : ( n19458 ) ;
assign n19460 =  ( n18934 ) ? ( bv_8_121_n470 ) : ( n19459 ) ;
assign n19461 =  ( n18932 ) ? ( bv_8_231_n99 ) : ( n19460 ) ;
assign n19462 =  ( n18930 ) ? ( bv_8_200_n213 ) : ( n19461 ) ;
assign n19463 =  ( n18928 ) ? ( bv_8_55_n650 ) : ( n19462 ) ;
assign n19464 =  ( n18926 ) ? ( bv_8_109_n9 ) : ( n19463 ) ;
assign n19465 =  ( n18924 ) ? ( bv_8_141_n410 ) : ( n19464 ) ;
assign n19466 =  ( n18922 ) ? ( bv_8_213_n167 ) : ( n19465 ) ;
assign n19467 =  ( n18920 ) ? ( bv_8_78_n590 ) : ( n19466 ) ;
assign n19468 =  ( n18918 ) ? ( bv_8_169_n109 ) : ( n19467 ) ;
assign n19469 =  ( n18916 ) ? ( bv_8_108_n510 ) : ( n19468 ) ;
assign n19470 =  ( n18914 ) ? ( bv_8_86_n567 ) : ( n19469 ) ;
assign n19471 =  ( n18912 ) ? ( bv_8_244_n47 ) : ( n19470 ) ;
assign n19472 =  ( n18910 ) ? ( bv_8_234_n87 ) : ( n19471 ) ;
assign n19473 =  ( n18908 ) ? ( bv_8_101_n49 ) : ( n19472 ) ;
assign n19474 =  ( n18906 ) ? ( bv_8_122_n416 ) : ( n19473 ) ;
assign n19475 =  ( n18904 ) ? ( bv_8_174_n152 ) : ( n19474 ) ;
assign n19476 =  ( n18902 ) ? ( bv_8_8_n669 ) : ( n19475 ) ;
assign n19477 =  ( n18900 ) ? ( bv_8_186_n263 ) : ( n19476 ) ;
assign n19478 =  ( n18898 ) ? ( bv_8_120_n474 ) : ( n19477 ) ;
assign n19479 =  ( n18896 ) ? ( bv_8_37_n506 ) : ( n19478 ) ;
assign n19480 =  ( n18894 ) ? ( bv_8_46_n429 ) : ( n19479 ) ;
assign n19481 =  ( n18892 ) ? ( bv_8_28_n162 ) : ( n19480 ) ;
assign n19482 =  ( n18890 ) ? ( bv_8_166_n328 ) : ( n19481 ) ;
assign n19483 =  ( n18888 ) ? ( bv_8_180_n285 ) : ( n19482 ) ;
assign n19484 =  ( n18886 ) ? ( bv_8_198_n220 ) : ( n19483 ) ;
assign n19485 =  ( n18884 ) ? ( bv_8_232_n95 ) : ( n19484 ) ;
assign n19486 =  ( n18882 ) ? ( bv_8_221_n138 ) : ( n19485 ) ;
assign n19487 =  ( n18880 ) ? ( bv_8_116_n345 ) : ( n19486 ) ;
assign n19488 =  ( n18878 ) ? ( bv_8_31_n705 ) : ( n19487 ) ;
assign n19489 =  ( n18876 ) ? ( bv_8_75_n503 ) : ( n19488 ) ;
assign n19490 =  ( n18874 ) ? ( bv_8_189_n254 ) : ( n19489 ) ;
assign n19491 =  ( n18872 ) ? ( bv_8_139_n297 ) : ( n19490 ) ;
assign n19492 =  ( n18870 ) ? ( bv_8_138_n418 ) : ( n19491 ) ;
assign n19493 =  ( n18868 ) ? ( bv_8_112_n482 ) : ( n19492 ) ;
assign n19494 =  ( n18866 ) ? ( bv_8_62_n205 ) : ( n19493 ) ;
assign n19495 =  ( n18864 ) ? ( bv_8_181_n281 ) : ( n19494 ) ;
assign n19496 =  ( n18862 ) ? ( bv_8_102_n527 ) : ( n19495 ) ;
assign n19497 =  ( n18860 ) ? ( bv_8_72_n330 ) : ( n19496 ) ;
assign n19498 =  ( n18858 ) ? ( bv_8_3_n65 ) : ( n19497 ) ;
assign n19499 =  ( n18856 ) ? ( bv_8_246_n39 ) : ( n19498 ) ;
assign n19500 =  ( n18854 ) ? ( bv_8_14_n648 ) : ( n19499 ) ;
assign n19501 =  ( n18852 ) ? ( bv_8_97_n198 ) : ( n19500 ) ;
assign n19502 =  ( n18850 ) ? ( bv_8_53_n436 ) : ( n19501 ) ;
assign n19503 =  ( n18848 ) ? ( bv_8_87_n226 ) : ( n19502 ) ;
assign n19504 =  ( n18846 ) ? ( bv_8_185_n266 ) : ( n19503 ) ;
assign n19505 =  ( n18844 ) ? ( bv_8_134_n431 ) : ( n19504 ) ;
assign n19506 =  ( n18842 ) ? ( bv_8_193_n239 ) : ( n19505 ) ;
assign n19507 =  ( n18840 ) ? ( bv_8_29_n625 ) : ( n19506 ) ;
assign n19508 =  ( n18838 ) ? ( bv_8_158_n355 ) : ( n19507 ) ;
assign n19509 =  ( n18836 ) ? ( bv_8_225_n123 ) : ( n19508 ) ;
assign n19510 =  ( n18834 ) ? ( bv_8_248_n31 ) : ( n19509 ) ;
assign n19511 =  ( n18832 ) ? ( bv_8_152_n374 ) : ( n19510 ) ;
assign n19512 =  ( n18830 ) ? ( bv_8_17_n525 ) : ( n19511 ) ;
assign n19513 =  ( n18828 ) ? ( bv_8_105_n148 ) : ( n19512 ) ;
assign n19514 =  ( n18826 ) ? ( bv_8_217_n128 ) : ( n19513 ) ;
assign n19515 =  ( n18824 ) ? ( bv_8_142_n406 ) : ( n19514 ) ;
assign n19516 =  ( n18822 ) ? ( bv_8_148_n388 ) : ( n19515 ) ;
assign n19517 =  ( n18820 ) ? ( bv_8_155_n364 ) : ( n19516 ) ;
assign n19518 =  ( n18818 ) ? ( bv_8_30_n21 ) : ( n19517 ) ;
assign n19519 =  ( n18816 ) ? ( bv_8_135_n81 ) : ( n19518 ) ;
assign n19520 =  ( n18814 ) ? ( bv_8_233_n91 ) : ( n19519 ) ;
assign n19521 =  ( n18812 ) ? ( bv_8_206_n192 ) : ( n19520 ) ;
assign n19522 =  ( n18810 ) ? ( bv_8_85_n423 ) : ( n19521 ) ;
assign n19523 =  ( n18808 ) ? ( bv_8_40_n366 ) : ( n19522 ) ;
assign n19524 =  ( n18806 ) ? ( bv_8_223_n130 ) : ( n19523 ) ;
assign n19525 =  ( n18804 ) ? ( bv_8_140_n376 ) : ( n19524 ) ;
assign n19526 =  ( n18802 ) ? ( bv_8_161_n211 ) : ( n19525 ) ;
assign n19527 =  ( n18800 ) ? ( bv_8_137_n421 ) : ( n19526 ) ;
assign n19528 =  ( n18798 ) ? ( bv_8_13_n194 ) : ( n19527 ) ;
assign n19529 =  ( n18796 ) ? ( bv_8_191_n246 ) : ( n19528 ) ;
assign n19530 =  ( n18794 ) ? ( bv_8_230_n103 ) : ( n19529 ) ;
assign n19531 =  ( n18792 ) ? ( bv_8_66_n466 ) : ( n19530 ) ;
assign n19532 =  ( n18790 ) ? ( bv_8_104_n520 ) : ( n19531 ) ;
assign n19533 =  ( n18788 ) ? ( bv_8_65_n623 ) : ( n19532 ) ;
assign n19534 =  ( n18786 ) ? ( bv_8_153_n140 ) : ( n19533 ) ;
assign n19535 =  ( n18784 ) ? ( bv_8_45_n97 ) : ( n19534 ) ;
assign n19536 =  ( n18782 ) ? ( bv_8_15_n190 ) : ( n19535 ) ;
assign n19537 =  ( n18780 ) ? ( bv_8_176_n299 ) : ( n19536 ) ;
assign n19538 =  ( n18778 ) ? ( bv_8_84_n386 ) : ( n19537 ) ;
assign n19539 =  ( n18776 ) ? ( bv_8_187_n260 ) : ( n19538 ) ;
assign n19540 =  ( n18774 ) ? ( bv_8_22_n357 ) : ( n19539 ) ;
assign n19541 = state_in[119:112] ;
assign n19542 =  ( n19541 ) == ( bv_8_255_n3 )  ;
assign n19543 = state_in[119:112] ;
assign n19544 =  ( n19543 ) == ( bv_8_254_n7 )  ;
assign n19545 = state_in[119:112] ;
assign n19546 =  ( n19545 ) == ( bv_8_253_n11 )  ;
assign n19547 = state_in[119:112] ;
assign n19548 =  ( n19547 ) == ( bv_8_252_n15 )  ;
assign n19549 = state_in[119:112] ;
assign n19550 =  ( n19549 ) == ( bv_8_251_n19 )  ;
assign n19551 = state_in[119:112] ;
assign n19552 =  ( n19551 ) == ( bv_8_250_n23 )  ;
assign n19553 = state_in[119:112] ;
assign n19554 =  ( n19553 ) == ( bv_8_249_n27 )  ;
assign n19555 = state_in[119:112] ;
assign n19556 =  ( n19555 ) == ( bv_8_248_n31 )  ;
assign n19557 = state_in[119:112] ;
assign n19558 =  ( n19557 ) == ( bv_8_247_n35 )  ;
assign n19559 = state_in[119:112] ;
assign n19560 =  ( n19559 ) == ( bv_8_246_n39 )  ;
assign n19561 = state_in[119:112] ;
assign n19562 =  ( n19561 ) == ( bv_8_245_n43 )  ;
assign n19563 = state_in[119:112] ;
assign n19564 =  ( n19563 ) == ( bv_8_244_n47 )  ;
assign n19565 = state_in[119:112] ;
assign n19566 =  ( n19565 ) == ( bv_8_243_n51 )  ;
assign n19567 = state_in[119:112] ;
assign n19568 =  ( n19567 ) == ( bv_8_242_n55 )  ;
assign n19569 = state_in[119:112] ;
assign n19570 =  ( n19569 ) == ( bv_8_241_n59 )  ;
assign n19571 = state_in[119:112] ;
assign n19572 =  ( n19571 ) == ( bv_8_240_n63 )  ;
assign n19573 = state_in[119:112] ;
assign n19574 =  ( n19573 ) == ( bv_8_239_n67 )  ;
assign n19575 = state_in[119:112] ;
assign n19576 =  ( n19575 ) == ( bv_8_238_n71 )  ;
assign n19577 = state_in[119:112] ;
assign n19578 =  ( n19577 ) == ( bv_8_237_n75 )  ;
assign n19579 = state_in[119:112] ;
assign n19580 =  ( n19579 ) == ( bv_8_236_n79 )  ;
assign n19581 = state_in[119:112] ;
assign n19582 =  ( n19581 ) == ( bv_8_235_n83 )  ;
assign n19583 = state_in[119:112] ;
assign n19584 =  ( n19583 ) == ( bv_8_234_n87 )  ;
assign n19585 = state_in[119:112] ;
assign n19586 =  ( n19585 ) == ( bv_8_233_n91 )  ;
assign n19587 = state_in[119:112] ;
assign n19588 =  ( n19587 ) == ( bv_8_232_n95 )  ;
assign n19589 = state_in[119:112] ;
assign n19590 =  ( n19589 ) == ( bv_8_231_n99 )  ;
assign n19591 = state_in[119:112] ;
assign n19592 =  ( n19591 ) == ( bv_8_230_n103 )  ;
assign n19593 = state_in[119:112] ;
assign n19594 =  ( n19593 ) == ( bv_8_229_n107 )  ;
assign n19595 = state_in[119:112] ;
assign n19596 =  ( n19595 ) == ( bv_8_228_n111 )  ;
assign n19597 = state_in[119:112] ;
assign n19598 =  ( n19597 ) == ( bv_8_227_n115 )  ;
assign n19599 = state_in[119:112] ;
assign n19600 =  ( n19599 ) == ( bv_8_226_n119 )  ;
assign n19601 = state_in[119:112] ;
assign n19602 =  ( n19601 ) == ( bv_8_225_n123 )  ;
assign n19603 = state_in[119:112] ;
assign n19604 =  ( n19603 ) == ( bv_8_224_n126 )  ;
assign n19605 = state_in[119:112] ;
assign n19606 =  ( n19605 ) == ( bv_8_223_n130 )  ;
assign n19607 = state_in[119:112] ;
assign n19608 =  ( n19607 ) == ( bv_8_222_n134 )  ;
assign n19609 = state_in[119:112] ;
assign n19610 =  ( n19609 ) == ( bv_8_221_n138 )  ;
assign n19611 = state_in[119:112] ;
assign n19612 =  ( n19611 ) == ( bv_8_220_n142 )  ;
assign n19613 = state_in[119:112] ;
assign n19614 =  ( n19613 ) == ( bv_8_219_n146 )  ;
assign n19615 = state_in[119:112] ;
assign n19616 =  ( n19615 ) == ( bv_8_218_n150 )  ;
assign n19617 = state_in[119:112] ;
assign n19618 =  ( n19617 ) == ( bv_8_217_n128 )  ;
assign n19619 = state_in[119:112] ;
assign n19620 =  ( n19619 ) == ( bv_8_216_n157 )  ;
assign n19621 = state_in[119:112] ;
assign n19622 =  ( n19621 ) == ( bv_8_215_n45 )  ;
assign n19623 = state_in[119:112] ;
assign n19624 =  ( n19623 ) == ( bv_8_214_n164 )  ;
assign n19625 = state_in[119:112] ;
assign n19626 =  ( n19625 ) == ( bv_8_213_n167 )  ;
assign n19627 = state_in[119:112] ;
assign n19628 =  ( n19627 ) == ( bv_8_212_n171 )  ;
assign n19629 = state_in[119:112] ;
assign n19630 =  ( n19629 ) == ( bv_8_211_n175 )  ;
assign n19631 = state_in[119:112] ;
assign n19632 =  ( n19631 ) == ( bv_8_210_n113 )  ;
assign n19633 = state_in[119:112] ;
assign n19634 =  ( n19633 ) == ( bv_8_209_n182 )  ;
assign n19635 = state_in[119:112] ;
assign n19636 =  ( n19635 ) == ( bv_8_208_n37 )  ;
assign n19637 = state_in[119:112] ;
assign n19638 =  ( n19637 ) == ( bv_8_207_n188 )  ;
assign n19639 = state_in[119:112] ;
assign n19640 =  ( n19639 ) == ( bv_8_206_n192 )  ;
assign n19641 = state_in[119:112] ;
assign n19642 =  ( n19641 ) == ( bv_8_205_n196 )  ;
assign n19643 = state_in[119:112] ;
assign n19644 =  ( n19643 ) == ( bv_8_204_n177 )  ;
assign n19645 = state_in[119:112] ;
assign n19646 =  ( n19645 ) == ( bv_8_203_n203 )  ;
assign n19647 = state_in[119:112] ;
assign n19648 =  ( n19647 ) == ( bv_8_202_n207 )  ;
assign n19649 = state_in[119:112] ;
assign n19650 =  ( n19649 ) == ( bv_8_201_n85 )  ;
assign n19651 = state_in[119:112] ;
assign n19652 =  ( n19651 ) == ( bv_8_200_n213 )  ;
assign n19653 = state_in[119:112] ;
assign n19654 =  ( n19653 ) == ( bv_8_199_n216 )  ;
assign n19655 = state_in[119:112] ;
assign n19656 =  ( n19655 ) == ( bv_8_198_n220 )  ;
assign n19657 = state_in[119:112] ;
assign n19658 =  ( n19657 ) == ( bv_8_197_n224 )  ;
assign n19659 = state_in[119:112] ;
assign n19660 =  ( n19659 ) == ( bv_8_196_n228 )  ;
assign n19661 = state_in[119:112] ;
assign n19662 =  ( n19661 ) == ( bv_8_195_n232 )  ;
assign n19663 = state_in[119:112] ;
assign n19664 =  ( n19663 ) == ( bv_8_194_n159 )  ;
assign n19665 = state_in[119:112] ;
assign n19666 =  ( n19665 ) == ( bv_8_193_n239 )  ;
assign n19667 = state_in[119:112] ;
assign n19668 =  ( n19667 ) == ( bv_8_192_n242 )  ;
assign n19669 = state_in[119:112] ;
assign n19670 =  ( n19669 ) == ( bv_8_191_n246 )  ;
assign n19671 = state_in[119:112] ;
assign n19672 =  ( n19671 ) == ( bv_8_190_n250 )  ;
assign n19673 = state_in[119:112] ;
assign n19674 =  ( n19673 ) == ( bv_8_189_n254 )  ;
assign n19675 = state_in[119:112] ;
assign n19676 =  ( n19675 ) == ( bv_8_188_n257 )  ;
assign n19677 = state_in[119:112] ;
assign n19678 =  ( n19677 ) == ( bv_8_187_n260 )  ;
assign n19679 = state_in[119:112] ;
assign n19680 =  ( n19679 ) == ( bv_8_186_n263 )  ;
assign n19681 = state_in[119:112] ;
assign n19682 =  ( n19681 ) == ( bv_8_185_n266 )  ;
assign n19683 = state_in[119:112] ;
assign n19684 =  ( n19683 ) == ( bv_8_184_n270 )  ;
assign n19685 = state_in[119:112] ;
assign n19686 =  ( n19685 ) == ( bv_8_183_n273 )  ;
assign n19687 = state_in[119:112] ;
assign n19688 =  ( n19687 ) == ( bv_8_182_n277 )  ;
assign n19689 = state_in[119:112] ;
assign n19690 =  ( n19689 ) == ( bv_8_181_n281 )  ;
assign n19691 = state_in[119:112] ;
assign n19692 =  ( n19691 ) == ( bv_8_180_n285 )  ;
assign n19693 = state_in[119:112] ;
assign n19694 =  ( n19693 ) == ( bv_8_179_n289 )  ;
assign n19695 = state_in[119:112] ;
assign n19696 =  ( n19695 ) == ( bv_8_178_n292 )  ;
assign n19697 = state_in[119:112] ;
assign n19698 =  ( n19697 ) == ( bv_8_177_n283 )  ;
assign n19699 = state_in[119:112] ;
assign n19700 =  ( n19699 ) == ( bv_8_176_n299 )  ;
assign n19701 = state_in[119:112] ;
assign n19702 =  ( n19701 ) == ( bv_8_175_n302 )  ;
assign n19703 = state_in[119:112] ;
assign n19704 =  ( n19703 ) == ( bv_8_174_n152 )  ;
assign n19705 = state_in[119:112] ;
assign n19706 =  ( n19705 ) == ( bv_8_173_n307 )  ;
assign n19707 = state_in[119:112] ;
assign n19708 =  ( n19707 ) == ( bv_8_172_n268 )  ;
assign n19709 = state_in[119:112] ;
assign n19710 =  ( n19709 ) == ( bv_8_171_n314 )  ;
assign n19711 = state_in[119:112] ;
assign n19712 =  ( n19711 ) == ( bv_8_170_n77 )  ;
assign n19713 = state_in[119:112] ;
assign n19714 =  ( n19713 ) == ( bv_8_169_n109 )  ;
assign n19715 = state_in[119:112] ;
assign n19716 =  ( n19715 ) == ( bv_8_168_n13 )  ;
assign n19717 = state_in[119:112] ;
assign n19718 =  ( n19717 ) == ( bv_8_167_n325 )  ;
assign n19719 = state_in[119:112] ;
assign n19720 =  ( n19719 ) == ( bv_8_166_n328 )  ;
assign n19721 = state_in[119:112] ;
assign n19722 =  ( n19721 ) == ( bv_8_165_n69 )  ;
assign n19723 = state_in[119:112] ;
assign n19724 =  ( n19723 ) == ( bv_8_164_n335 )  ;
assign n19725 = state_in[119:112] ;
assign n19726 =  ( n19725 ) == ( bv_8_163_n339 )  ;
assign n19727 = state_in[119:112] ;
assign n19728 =  ( n19727 ) == ( bv_8_162_n343 )  ;
assign n19729 = state_in[119:112] ;
assign n19730 =  ( n19729 ) == ( bv_8_161_n211 )  ;
assign n19731 = state_in[119:112] ;
assign n19732 =  ( n19731 ) == ( bv_8_160_n350 )  ;
assign n19733 = state_in[119:112] ;
assign n19734 =  ( n19733 ) == ( bv_8_159_n323 )  ;
assign n19735 = state_in[119:112] ;
assign n19736 =  ( n19735 ) == ( bv_8_158_n355 )  ;
assign n19737 = state_in[119:112] ;
assign n19738 =  ( n19737 ) == ( bv_8_157_n359 )  ;
assign n19739 = state_in[119:112] ;
assign n19740 =  ( n19739 ) == ( bv_8_156_n279 )  ;
assign n19741 = state_in[119:112] ;
assign n19742 =  ( n19741 ) == ( bv_8_155_n364 )  ;
assign n19743 = state_in[119:112] ;
assign n19744 =  ( n19743 ) == ( bv_8_154_n368 )  ;
assign n19745 = state_in[119:112] ;
assign n19746 =  ( n19745 ) == ( bv_8_153_n140 )  ;
assign n19747 = state_in[119:112] ;
assign n19748 =  ( n19747 ) == ( bv_8_152_n374 )  ;
assign n19749 = state_in[119:112] ;
assign n19750 =  ( n19749 ) == ( bv_8_151_n218 )  ;
assign n19751 = state_in[119:112] ;
assign n19752 =  ( n19751 ) == ( bv_8_150_n201 )  ;
assign n19753 = state_in[119:112] ;
assign n19754 =  ( n19753 ) == ( bv_8_149_n384 )  ;
assign n19755 = state_in[119:112] ;
assign n19756 =  ( n19755 ) == ( bv_8_148_n388 )  ;
assign n19757 = state_in[119:112] ;
assign n19758 =  ( n19757 ) == ( bv_8_147_n392 )  ;
assign n19759 = state_in[119:112] ;
assign n19760 =  ( n19759 ) == ( bv_8_146_n337 )  ;
assign n19761 = state_in[119:112] ;
assign n19762 =  ( n19761 ) == ( bv_8_145_n397 )  ;
assign n19763 = state_in[119:112] ;
assign n19764 =  ( n19763 ) == ( bv_8_144_n173 )  ;
assign n19765 = state_in[119:112] ;
assign n19766 =  ( n19765 ) == ( bv_8_143_n403 )  ;
assign n19767 = state_in[119:112] ;
assign n19768 =  ( n19767 ) == ( bv_8_142_n406 )  ;
assign n19769 = state_in[119:112] ;
assign n19770 =  ( n19769 ) == ( bv_8_141_n410 )  ;
assign n19771 = state_in[119:112] ;
assign n19772 =  ( n19771 ) == ( bv_8_140_n376 )  ;
assign n19773 = state_in[119:112] ;
assign n19774 =  ( n19773 ) == ( bv_8_139_n297 )  ;
assign n19775 = state_in[119:112] ;
assign n19776 =  ( n19775 ) == ( bv_8_138_n418 )  ;
assign n19777 = state_in[119:112] ;
assign n19778 =  ( n19777 ) == ( bv_8_137_n421 )  ;
assign n19779 = state_in[119:112] ;
assign n19780 =  ( n19779 ) == ( bv_8_136_n425 )  ;
assign n19781 = state_in[119:112] ;
assign n19782 =  ( n19781 ) == ( bv_8_135_n81 )  ;
assign n19783 = state_in[119:112] ;
assign n19784 =  ( n19783 ) == ( bv_8_134_n431 )  ;
assign n19785 = state_in[119:112] ;
assign n19786 =  ( n19785 ) == ( bv_8_133_n434 )  ;
assign n19787 = state_in[119:112] ;
assign n19788 =  ( n19787 ) == ( bv_8_132_n41 )  ;
assign n19789 = state_in[119:112] ;
assign n19790 =  ( n19789 ) == ( bv_8_131_n440 )  ;
assign n19791 = state_in[119:112] ;
assign n19792 =  ( n19791 ) == ( bv_8_130_n33 )  ;
assign n19793 = state_in[119:112] ;
assign n19794 =  ( n19793 ) == ( bv_8_129_n446 )  ;
assign n19795 = state_in[119:112] ;
assign n19796 =  ( n19795 ) == ( bv_8_128_n450 )  ;
assign n19797 = state_in[119:112] ;
assign n19798 =  ( n19797 ) == ( bv_8_127_n453 )  ;
assign n19799 = state_in[119:112] ;
assign n19800 =  ( n19799 ) == ( bv_8_126_n456 )  ;
assign n19801 = state_in[119:112] ;
assign n19802 =  ( n19801 ) == ( bv_8_125_n459 )  ;
assign n19803 = state_in[119:112] ;
assign n19804 =  ( n19803 ) == ( bv_8_124_n184 )  ;
assign n19805 = state_in[119:112] ;
assign n19806 =  ( n19805 ) == ( bv_8_123_n17 )  ;
assign n19807 = state_in[119:112] ;
assign n19808 =  ( n19807 ) == ( bv_8_122_n416 )  ;
assign n19809 = state_in[119:112] ;
assign n19810 =  ( n19809 ) == ( bv_8_121_n470 )  ;
assign n19811 = state_in[119:112] ;
assign n19812 =  ( n19811 ) == ( bv_8_120_n474 )  ;
assign n19813 = state_in[119:112] ;
assign n19814 =  ( n19813 ) == ( bv_8_119_n472 )  ;
assign n19815 = state_in[119:112] ;
assign n19816 =  ( n19815 ) == ( bv_8_118_n480 )  ;
assign n19817 = state_in[119:112] ;
assign n19818 =  ( n19817 ) == ( bv_8_117_n484 )  ;
assign n19819 = state_in[119:112] ;
assign n19820 =  ( n19819 ) == ( bv_8_116_n345 )  ;
assign n19821 = state_in[119:112] ;
assign n19822 =  ( n19821 ) == ( bv_8_115_n222 )  ;
assign n19823 = state_in[119:112] ;
assign n19824 =  ( n19823 ) == ( bv_8_114_n494 )  ;
assign n19825 = state_in[119:112] ;
assign n19826 =  ( n19825 ) == ( bv_8_113_n180 )  ;
assign n19827 = state_in[119:112] ;
assign n19828 =  ( n19827 ) == ( bv_8_112_n482 )  ;
assign n19829 = state_in[119:112] ;
assign n19830 =  ( n19829 ) == ( bv_8_111_n244 )  ;
assign n19831 = state_in[119:112] ;
assign n19832 =  ( n19831 ) == ( bv_8_110_n294 )  ;
assign n19833 = state_in[119:112] ;
assign n19834 =  ( n19833 ) == ( bv_8_109_n9 )  ;
assign n19835 = state_in[119:112] ;
assign n19836 =  ( n19835 ) == ( bv_8_108_n510 )  ;
assign n19837 = state_in[119:112] ;
assign n19838 =  ( n19837 ) == ( bv_8_107_n370 )  ;
assign n19839 = state_in[119:112] ;
assign n19840 =  ( n19839 ) == ( bv_8_106_n155 )  ;
assign n19841 = state_in[119:112] ;
assign n19842 =  ( n19841 ) == ( bv_8_105_n148 )  ;
assign n19843 = state_in[119:112] ;
assign n19844 =  ( n19843 ) == ( bv_8_104_n520 )  ;
assign n19845 = state_in[119:112] ;
assign n19846 =  ( n19845 ) == ( bv_8_103_n523 )  ;
assign n19847 = state_in[119:112] ;
assign n19848 =  ( n19847 ) == ( bv_8_102_n527 )  ;
assign n19849 = state_in[119:112] ;
assign n19850 =  ( n19849 ) == ( bv_8_101_n49 )  ;
assign n19851 = state_in[119:112] ;
assign n19852 =  ( n19851 ) == ( bv_8_100_n348 )  ;
assign n19853 = state_in[119:112] ;
assign n19854 =  ( n19853 ) == ( bv_8_99_n476 )  ;
assign n19855 = state_in[119:112] ;
assign n19856 =  ( n19855 ) == ( bv_8_98_n536 )  ;
assign n19857 = state_in[119:112] ;
assign n19858 =  ( n19857 ) == ( bv_8_97_n198 )  ;
assign n19859 = state_in[119:112] ;
assign n19860 =  ( n19859 ) == ( bv_8_96_n542 )  ;
assign n19861 = state_in[119:112] ;
assign n19862 =  ( n19861 ) == ( bv_8_95_n545 )  ;
assign n19863 = state_in[119:112] ;
assign n19864 =  ( n19863 ) == ( bv_8_94_n548 )  ;
assign n19865 = state_in[119:112] ;
assign n19866 =  ( n19865 ) == ( bv_8_93_n498 )  ;
assign n19867 = state_in[119:112] ;
assign n19868 =  ( n19867 ) == ( bv_8_92_n234 )  ;
assign n19869 = state_in[119:112] ;
assign n19870 =  ( n19869 ) == ( bv_8_91_n555 )  ;
assign n19871 = state_in[119:112] ;
assign n19872 =  ( n19871 ) == ( bv_8_90_n25 )  ;
assign n19873 = state_in[119:112] ;
assign n19874 =  ( n19873 ) == ( bv_8_89_n61 )  ;
assign n19875 = state_in[119:112] ;
assign n19876 =  ( n19875 ) == ( bv_8_88_n562 )  ;
assign n19877 = state_in[119:112] ;
assign n19878 =  ( n19877 ) == ( bv_8_87_n226 )  ;
assign n19879 = state_in[119:112] ;
assign n19880 =  ( n19879 ) == ( bv_8_86_n567 )  ;
assign n19881 = state_in[119:112] ;
assign n19882 =  ( n19881 ) == ( bv_8_85_n423 )  ;
assign n19883 = state_in[119:112] ;
assign n19884 =  ( n19883 ) == ( bv_8_84_n386 )  ;
assign n19885 = state_in[119:112] ;
assign n19886 =  ( n19885 ) == ( bv_8_83_n575 )  ;
assign n19887 = state_in[119:112] ;
assign n19888 =  ( n19887 ) == ( bv_8_82_n578 )  ;
assign n19889 = state_in[119:112] ;
assign n19890 =  ( n19889 ) == ( bv_8_81_n582 )  ;
assign n19891 = state_in[119:112] ;
assign n19892 =  ( n19891 ) == ( bv_8_80_n73 )  ;
assign n19893 = state_in[119:112] ;
assign n19894 =  ( n19893 ) == ( bv_8_79_n538 )  ;
assign n19895 = state_in[119:112] ;
assign n19896 =  ( n19895 ) == ( bv_8_78_n590 )  ;
assign n19897 = state_in[119:112] ;
assign n19898 =  ( n19897 ) == ( bv_8_77_n593 )  ;
assign n19899 = state_in[119:112] ;
assign n19900 =  ( n19899 ) == ( bv_8_76_n596 )  ;
assign n19901 = state_in[119:112] ;
assign n19902 =  ( n19901 ) == ( bv_8_75_n503 )  ;
assign n19903 = state_in[119:112] ;
assign n19904 =  ( n19903 ) == ( bv_8_74_n237 )  ;
assign n19905 = state_in[119:112] ;
assign n19906 =  ( n19905 ) == ( bv_8_73_n275 )  ;
assign n19907 = state_in[119:112] ;
assign n19908 =  ( n19907 ) == ( bv_8_72_n330 )  ;
assign n19909 = state_in[119:112] ;
assign n19910 =  ( n19909 ) == ( bv_8_71_n252 )  ;
assign n19911 = state_in[119:112] ;
assign n19912 =  ( n19911 ) == ( bv_8_70_n609 )  ;
assign n19913 = state_in[119:112] ;
assign n19914 =  ( n19913 ) == ( bv_8_69_n612 )  ;
assign n19915 = state_in[119:112] ;
assign n19916 =  ( n19915 ) == ( bv_8_68_n390 )  ;
assign n19917 = state_in[119:112] ;
assign n19918 =  ( n19917 ) == ( bv_8_67_n318 )  ;
assign n19919 = state_in[119:112] ;
assign n19920 =  ( n19919 ) == ( bv_8_66_n466 )  ;
assign n19921 = state_in[119:112] ;
assign n19922 =  ( n19921 ) == ( bv_8_65_n623 )  ;
assign n19923 = state_in[119:112] ;
assign n19924 =  ( n19923 ) == ( bv_8_64_n573 )  ;
assign n19925 = state_in[119:112] ;
assign n19926 =  ( n19925 ) == ( bv_8_63_n489 )  ;
assign n19927 = state_in[119:112] ;
assign n19928 =  ( n19927 ) == ( bv_8_62_n205 )  ;
assign n19929 = state_in[119:112] ;
assign n19930 =  ( n19929 ) == ( bv_8_61_n634 )  ;
assign n19931 = state_in[119:112] ;
assign n19932 =  ( n19931 ) == ( bv_8_60_n93 )  ;
assign n19933 = state_in[119:112] ;
assign n19934 =  ( n19933 ) == ( bv_8_59_n382 )  ;
assign n19935 = state_in[119:112] ;
assign n19936 =  ( n19935 ) == ( bv_8_58_n136 )  ;
assign n19937 = state_in[119:112] ;
assign n19938 =  ( n19937 ) == ( bv_8_57_n312 )  ;
assign n19939 = state_in[119:112] ;
assign n19940 =  ( n19939 ) == ( bv_8_56_n230 )  ;
assign n19941 = state_in[119:112] ;
assign n19942 =  ( n19941 ) == ( bv_8_55_n650 )  ;
assign n19943 = state_in[119:112] ;
assign n19944 =  ( n19943 ) == ( bv_8_54_n616 )  ;
assign n19945 = state_in[119:112] ;
assign n19946 =  ( n19945 ) == ( bv_8_53_n436 )  ;
assign n19947 = state_in[119:112] ;
assign n19948 =  ( n19947 ) == ( bv_8_52_n619 )  ;
assign n19949 = state_in[119:112] ;
assign n19950 =  ( n19949 ) == ( bv_8_51_n101 )  ;
assign n19951 = state_in[119:112] ;
assign n19952 =  ( n19951 ) == ( bv_8_50_n408 )  ;
assign n19953 = state_in[119:112] ;
assign n19954 =  ( n19953 ) == ( bv_8_49_n309 )  ;
assign n19955 = state_in[119:112] ;
assign n19956 =  ( n19955 ) == ( bv_8_48_n660 )  ;
assign n19957 = state_in[119:112] ;
assign n19958 =  ( n19957 ) == ( bv_8_47_n652 )  ;
assign n19959 = state_in[119:112] ;
assign n19960 =  ( n19959 ) == ( bv_8_46_n429 )  ;
assign n19961 = state_in[119:112] ;
assign n19962 =  ( n19961 ) == ( bv_8_45_n97 )  ;
assign n19963 = state_in[119:112] ;
assign n19964 =  ( n19963 ) == ( bv_8_44_n5 )  ;
assign n19965 = state_in[119:112] ;
assign n19966 =  ( n19965 ) == ( bv_8_43_n121 )  ;
assign n19967 = state_in[119:112] ;
assign n19968 =  ( n19967 ) == ( bv_8_42_n672 )  ;
assign n19969 = state_in[119:112] ;
assign n19970 =  ( n19969 ) == ( bv_8_41_n29 )  ;
assign n19971 = state_in[119:112] ;
assign n19972 =  ( n19971 ) == ( bv_8_40_n366 )  ;
assign n19973 = state_in[119:112] ;
assign n19974 =  ( n19973 ) == ( bv_8_39_n132 )  ;
assign n19975 = state_in[119:112] ;
assign n19976 =  ( n19975 ) == ( bv_8_38_n444 )  ;
assign n19977 = state_in[119:112] ;
assign n19978 =  ( n19977 ) == ( bv_8_37_n506 )  ;
assign n19979 = state_in[119:112] ;
assign n19980 =  ( n19979 ) == ( bv_8_36_n645 )  ;
assign n19981 = state_in[119:112] ;
assign n19982 =  ( n19981 ) == ( bv_8_35_n696 )  ;
assign n19983 = state_in[119:112] ;
assign n19984 =  ( n19983 ) == ( bv_8_34_n117 )  ;
assign n19985 = state_in[119:112] ;
assign n19986 =  ( n19985 ) == ( bv_8_33_n486 )  ;
assign n19987 = state_in[119:112] ;
assign n19988 =  ( n19987 ) == ( bv_8_32_n463 )  ;
assign n19989 = state_in[119:112] ;
assign n19990 =  ( n19989 ) == ( bv_8_31_n705 )  ;
assign n19991 = state_in[119:112] ;
assign n19992 =  ( n19991 ) == ( bv_8_30_n21 )  ;
assign n19993 = state_in[119:112] ;
assign n19994 =  ( n19993 ) == ( bv_8_29_n625 )  ;
assign n19995 = state_in[119:112] ;
assign n19996 =  ( n19995 ) == ( bv_8_28_n162 )  ;
assign n19997 = state_in[119:112] ;
assign n19998 =  ( n19997 ) == ( bv_8_27_n642 )  ;
assign n19999 = state_in[119:112] ;
assign n20000 =  ( n19999 ) == ( bv_8_26_n53 )  ;
assign n20001 = state_in[119:112] ;
assign n20002 =  ( n20001 ) == ( bv_8_25_n399 )  ;
assign n20003 = state_in[119:112] ;
assign n20004 =  ( n20003 ) == ( bv_8_24_n448 )  ;
assign n20005 = state_in[119:112] ;
assign n20006 =  ( n20005 ) == ( bv_8_23_n144 )  ;
assign n20007 = state_in[119:112] ;
assign n20008 =  ( n20007 ) == ( bv_8_22_n357 )  ;
assign n20009 = state_in[119:112] ;
assign n20010 =  ( n20009 ) == ( bv_8_21_n89 )  ;
assign n20011 = state_in[119:112] ;
assign n20012 =  ( n20011 ) == ( bv_8_20_n341 )  ;
assign n20013 = state_in[119:112] ;
assign n20014 =  ( n20013 ) == ( bv_8_19_n588 )  ;
assign n20015 = state_in[119:112] ;
assign n20016 =  ( n20015 ) == ( bv_8_18_n628 )  ;
assign n20017 = state_in[119:112] ;
assign n20018 =  ( n20017 ) == ( bv_8_17_n525 )  ;
assign n20019 = state_in[119:112] ;
assign n20020 =  ( n20019 ) == ( bv_8_16_n248 )  ;
assign n20021 = state_in[119:112] ;
assign n20022 =  ( n20021 ) == ( bv_8_15_n190 )  ;
assign n20023 = state_in[119:112] ;
assign n20024 =  ( n20023 ) == ( bv_8_14_n648 )  ;
assign n20025 = state_in[119:112] ;
assign n20026 =  ( n20025 ) == ( bv_8_13_n194 )  ;
assign n20027 = state_in[119:112] ;
assign n20028 =  ( n20027 ) == ( bv_8_12_n333 )  ;
assign n20029 = state_in[119:112] ;
assign n20030 =  ( n20029 ) == ( bv_8_11_n379 )  ;
assign n20031 = state_in[119:112] ;
assign n20032 =  ( n20031 ) == ( bv_8_10_n655 )  ;
assign n20033 = state_in[119:112] ;
assign n20034 =  ( n20033 ) == ( bv_8_9_n57 )  ;
assign n20035 = state_in[119:112] ;
assign n20036 =  ( n20035 ) == ( bv_8_8_n669 )  ;
assign n20037 = state_in[119:112] ;
assign n20038 =  ( n20037 ) == ( bv_8_7_n105 )  ;
assign n20039 = state_in[119:112] ;
assign n20040 =  ( n20039 ) == ( bv_8_6_n169 )  ;
assign n20041 = state_in[119:112] ;
assign n20042 =  ( n20041 ) == ( bv_8_5_n492 )  ;
assign n20043 = state_in[119:112] ;
assign n20044 =  ( n20043 ) == ( bv_8_4_n516 )  ;
assign n20045 = state_in[119:112] ;
assign n20046 =  ( n20045 ) == ( bv_8_3_n65 )  ;
assign n20047 = state_in[119:112] ;
assign n20048 =  ( n20047 ) == ( bv_8_2_n751 )  ;
assign n20049 = state_in[119:112] ;
assign n20050 =  ( n20049 ) == ( bv_8_1_n287 )  ;
assign n20051 = state_in[119:112] ;
assign n20052 =  ( n20051 ) == ( bv_8_0_n580 )  ;
assign n20053 =  ( n20052 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n20054 =  ( n20050 ) ? ( bv_8_248_n31 ) : ( n20053 ) ;
assign n20055 =  ( n20048 ) ? ( bv_8_238_n71 ) : ( n20054 ) ;
assign n20056 =  ( n20046 ) ? ( bv_8_246_n39 ) : ( n20055 ) ;
assign n20057 =  ( n20044 ) ? ( bv_8_255_n3 ) : ( n20056 ) ;
assign n20058 =  ( n20042 ) ? ( bv_8_214_n164 ) : ( n20057 ) ;
assign n20059 =  ( n20040 ) ? ( bv_8_222_n134 ) : ( n20058 ) ;
assign n20060 =  ( n20038 ) ? ( bv_8_145_n397 ) : ( n20059 ) ;
assign n20061 =  ( n20036 ) ? ( bv_8_96_n542 ) : ( n20060 ) ;
assign n20062 =  ( n20034 ) ? ( bv_8_2_n751 ) : ( n20061 ) ;
assign n20063 =  ( n20032 ) ? ( bv_8_206_n192 ) : ( n20062 ) ;
assign n20064 =  ( n20030 ) ? ( bv_8_86_n567 ) : ( n20063 ) ;
assign n20065 =  ( n20028 ) ? ( bv_8_231_n99 ) : ( n20064 ) ;
assign n20066 =  ( n20026 ) ? ( bv_8_181_n281 ) : ( n20065 ) ;
assign n20067 =  ( n20024 ) ? ( bv_8_77_n593 ) : ( n20066 ) ;
assign n20068 =  ( n20022 ) ? ( bv_8_236_n79 ) : ( n20067 ) ;
assign n20069 =  ( n20020 ) ? ( bv_8_143_n403 ) : ( n20068 ) ;
assign n20070 =  ( n20018 ) ? ( bv_8_31_n705 ) : ( n20069 ) ;
assign n20071 =  ( n20016 ) ? ( bv_8_137_n421 ) : ( n20070 ) ;
assign n20072 =  ( n20014 ) ? ( bv_8_250_n23 ) : ( n20071 ) ;
assign n20073 =  ( n20012 ) ? ( bv_8_239_n67 ) : ( n20072 ) ;
assign n20074 =  ( n20010 ) ? ( bv_8_178_n292 ) : ( n20073 ) ;
assign n20075 =  ( n20008 ) ? ( bv_8_142_n406 ) : ( n20074 ) ;
assign n20076 =  ( n20006 ) ? ( bv_8_251_n19 ) : ( n20075 ) ;
assign n20077 =  ( n20004 ) ? ( bv_8_65_n623 ) : ( n20076 ) ;
assign n20078 =  ( n20002 ) ? ( bv_8_179_n289 ) : ( n20077 ) ;
assign n20079 =  ( n20000 ) ? ( bv_8_95_n545 ) : ( n20078 ) ;
assign n20080 =  ( n19998 ) ? ( bv_8_69_n612 ) : ( n20079 ) ;
assign n20081 =  ( n19996 ) ? ( bv_8_35_n696 ) : ( n20080 ) ;
assign n20082 =  ( n19994 ) ? ( bv_8_83_n575 ) : ( n20081 ) ;
assign n20083 =  ( n19992 ) ? ( bv_8_228_n111 ) : ( n20082 ) ;
assign n20084 =  ( n19990 ) ? ( bv_8_155_n364 ) : ( n20083 ) ;
assign n20085 =  ( n19988 ) ? ( bv_8_117_n484 ) : ( n20084 ) ;
assign n20086 =  ( n19986 ) ? ( bv_8_225_n123 ) : ( n20085 ) ;
assign n20087 =  ( n19984 ) ? ( bv_8_61_n634 ) : ( n20086 ) ;
assign n20088 =  ( n19982 ) ? ( bv_8_76_n596 ) : ( n20087 ) ;
assign n20089 =  ( n19980 ) ? ( bv_8_108_n510 ) : ( n20088 ) ;
assign n20090 =  ( n19978 ) ? ( bv_8_126_n456 ) : ( n20089 ) ;
assign n20091 =  ( n19976 ) ? ( bv_8_245_n43 ) : ( n20090 ) ;
assign n20092 =  ( n19974 ) ? ( bv_8_131_n440 ) : ( n20091 ) ;
assign n20093 =  ( n19972 ) ? ( bv_8_104_n520 ) : ( n20092 ) ;
assign n20094 =  ( n19970 ) ? ( bv_8_81_n582 ) : ( n20093 ) ;
assign n20095 =  ( n19968 ) ? ( bv_8_209_n182 ) : ( n20094 ) ;
assign n20096 =  ( n19966 ) ? ( bv_8_249_n27 ) : ( n20095 ) ;
assign n20097 =  ( n19964 ) ? ( bv_8_226_n119 ) : ( n20096 ) ;
assign n20098 =  ( n19962 ) ? ( bv_8_171_n314 ) : ( n20097 ) ;
assign n20099 =  ( n19960 ) ? ( bv_8_98_n536 ) : ( n20098 ) ;
assign n20100 =  ( n19958 ) ? ( bv_8_42_n672 ) : ( n20099 ) ;
assign n20101 =  ( n19956 ) ? ( bv_8_8_n669 ) : ( n20100 ) ;
assign n20102 =  ( n19954 ) ? ( bv_8_149_n384 ) : ( n20101 ) ;
assign n20103 =  ( n19952 ) ? ( bv_8_70_n609 ) : ( n20102 ) ;
assign n20104 =  ( n19950 ) ? ( bv_8_157_n359 ) : ( n20103 ) ;
assign n20105 =  ( n19948 ) ? ( bv_8_48_n660 ) : ( n20104 ) ;
assign n20106 =  ( n19946 ) ? ( bv_8_55_n650 ) : ( n20105 ) ;
assign n20107 =  ( n19944 ) ? ( bv_8_10_n655 ) : ( n20106 ) ;
assign n20108 =  ( n19942 ) ? ( bv_8_47_n652 ) : ( n20107 ) ;
assign n20109 =  ( n19940 ) ? ( bv_8_14_n648 ) : ( n20108 ) ;
assign n20110 =  ( n19938 ) ? ( bv_8_36_n645 ) : ( n20109 ) ;
assign n20111 =  ( n19936 ) ? ( bv_8_27_n642 ) : ( n20110 ) ;
assign n20112 =  ( n19934 ) ? ( bv_8_223_n130 ) : ( n20111 ) ;
assign n20113 =  ( n19932 ) ? ( bv_8_205_n196 ) : ( n20112 ) ;
assign n20114 =  ( n19930 ) ? ( bv_8_78_n590 ) : ( n20113 ) ;
assign n20115 =  ( n19928 ) ? ( bv_8_127_n453 ) : ( n20114 ) ;
assign n20116 =  ( n19926 ) ? ( bv_8_234_n87 ) : ( n20115 ) ;
assign n20117 =  ( n19924 ) ? ( bv_8_18_n628 ) : ( n20116 ) ;
assign n20118 =  ( n19922 ) ? ( bv_8_29_n625 ) : ( n20117 ) ;
assign n20119 =  ( n19920 ) ? ( bv_8_88_n562 ) : ( n20118 ) ;
assign n20120 =  ( n19918 ) ? ( bv_8_52_n619 ) : ( n20119 ) ;
assign n20121 =  ( n19916 ) ? ( bv_8_54_n616 ) : ( n20120 ) ;
assign n20122 =  ( n19914 ) ? ( bv_8_220_n142 ) : ( n20121 ) ;
assign n20123 =  ( n19912 ) ? ( bv_8_180_n285 ) : ( n20122 ) ;
assign n20124 =  ( n19910 ) ? ( bv_8_91_n555 ) : ( n20123 ) ;
assign n20125 =  ( n19908 ) ? ( bv_8_164_n335 ) : ( n20124 ) ;
assign n20126 =  ( n19906 ) ? ( bv_8_118_n480 ) : ( n20125 ) ;
assign n20127 =  ( n19904 ) ? ( bv_8_183_n273 ) : ( n20126 ) ;
assign n20128 =  ( n19902 ) ? ( bv_8_125_n459 ) : ( n20127 ) ;
assign n20129 =  ( n19900 ) ? ( bv_8_82_n578 ) : ( n20128 ) ;
assign n20130 =  ( n19898 ) ? ( bv_8_221_n138 ) : ( n20129 ) ;
assign n20131 =  ( n19896 ) ? ( bv_8_94_n548 ) : ( n20130 ) ;
assign n20132 =  ( n19894 ) ? ( bv_8_19_n588 ) : ( n20131 ) ;
assign n20133 =  ( n19892 ) ? ( bv_8_166_n328 ) : ( n20132 ) ;
assign n20134 =  ( n19890 ) ? ( bv_8_185_n266 ) : ( n20133 ) ;
assign n20135 =  ( n19888 ) ? ( bv_8_0_n580 ) : ( n20134 ) ;
assign n20136 =  ( n19886 ) ? ( bv_8_193_n239 ) : ( n20135 ) ;
assign n20137 =  ( n19884 ) ? ( bv_8_64_n573 ) : ( n20136 ) ;
assign n20138 =  ( n19882 ) ? ( bv_8_227_n115 ) : ( n20137 ) ;
assign n20139 =  ( n19880 ) ? ( bv_8_121_n470 ) : ( n20138 ) ;
assign n20140 =  ( n19878 ) ? ( bv_8_182_n277 ) : ( n20139 ) ;
assign n20141 =  ( n19876 ) ? ( bv_8_212_n171 ) : ( n20140 ) ;
assign n20142 =  ( n19874 ) ? ( bv_8_141_n410 ) : ( n20141 ) ;
assign n20143 =  ( n19872 ) ? ( bv_8_103_n523 ) : ( n20142 ) ;
assign n20144 =  ( n19870 ) ? ( bv_8_114_n494 ) : ( n20143 ) ;
assign n20145 =  ( n19868 ) ? ( bv_8_148_n388 ) : ( n20144 ) ;
assign n20146 =  ( n19866 ) ? ( bv_8_152_n374 ) : ( n20145 ) ;
assign n20147 =  ( n19864 ) ? ( bv_8_176_n299 ) : ( n20146 ) ;
assign n20148 =  ( n19862 ) ? ( bv_8_133_n434 ) : ( n20147 ) ;
assign n20149 =  ( n19860 ) ? ( bv_8_187_n260 ) : ( n20148 ) ;
assign n20150 =  ( n19858 ) ? ( bv_8_197_n224 ) : ( n20149 ) ;
assign n20151 =  ( n19856 ) ? ( bv_8_79_n538 ) : ( n20150 ) ;
assign n20152 =  ( n19854 ) ? ( bv_8_237_n75 ) : ( n20151 ) ;
assign n20153 =  ( n19852 ) ? ( bv_8_134_n431 ) : ( n20152 ) ;
assign n20154 =  ( n19850 ) ? ( bv_8_154_n368 ) : ( n20153 ) ;
assign n20155 =  ( n19848 ) ? ( bv_8_102_n527 ) : ( n20154 ) ;
assign n20156 =  ( n19846 ) ? ( bv_8_17_n525 ) : ( n20155 ) ;
assign n20157 =  ( n19844 ) ? ( bv_8_138_n418 ) : ( n20156 ) ;
assign n20158 =  ( n19842 ) ? ( bv_8_233_n91 ) : ( n20157 ) ;
assign n20159 =  ( n19840 ) ? ( bv_8_4_n516 ) : ( n20158 ) ;
assign n20160 =  ( n19838 ) ? ( bv_8_254_n7 ) : ( n20159 ) ;
assign n20161 =  ( n19836 ) ? ( bv_8_160_n350 ) : ( n20160 ) ;
assign n20162 =  ( n19834 ) ? ( bv_8_120_n474 ) : ( n20161 ) ;
assign n20163 =  ( n19832 ) ? ( bv_8_37_n506 ) : ( n20162 ) ;
assign n20164 =  ( n19830 ) ? ( bv_8_75_n503 ) : ( n20163 ) ;
assign n20165 =  ( n19828 ) ? ( bv_8_162_n343 ) : ( n20164 ) ;
assign n20166 =  ( n19826 ) ? ( bv_8_93_n498 ) : ( n20165 ) ;
assign n20167 =  ( n19824 ) ? ( bv_8_128_n450 ) : ( n20166 ) ;
assign n20168 =  ( n19822 ) ? ( bv_8_5_n492 ) : ( n20167 ) ;
assign n20169 =  ( n19820 ) ? ( bv_8_63_n489 ) : ( n20168 ) ;
assign n20170 =  ( n19818 ) ? ( bv_8_33_n486 ) : ( n20169 ) ;
assign n20171 =  ( n19816 ) ? ( bv_8_112_n482 ) : ( n20170 ) ;
assign n20172 =  ( n19814 ) ? ( bv_8_241_n59 ) : ( n20171 ) ;
assign n20173 =  ( n19812 ) ? ( bv_8_99_n476 ) : ( n20172 ) ;
assign n20174 =  ( n19810 ) ? ( bv_8_119_n472 ) : ( n20173 ) ;
assign n20175 =  ( n19808 ) ? ( bv_8_175_n302 ) : ( n20174 ) ;
assign n20176 =  ( n19806 ) ? ( bv_8_66_n466 ) : ( n20175 ) ;
assign n20177 =  ( n19804 ) ? ( bv_8_32_n463 ) : ( n20176 ) ;
assign n20178 =  ( n19802 ) ? ( bv_8_229_n107 ) : ( n20177 ) ;
assign n20179 =  ( n19800 ) ? ( bv_8_253_n11 ) : ( n20178 ) ;
assign n20180 =  ( n19798 ) ? ( bv_8_191_n246 ) : ( n20179 ) ;
assign n20181 =  ( n19796 ) ? ( bv_8_129_n446 ) : ( n20180 ) ;
assign n20182 =  ( n19794 ) ? ( bv_8_24_n448 ) : ( n20181 ) ;
assign n20183 =  ( n19792 ) ? ( bv_8_38_n444 ) : ( n20182 ) ;
assign n20184 =  ( n19790 ) ? ( bv_8_195_n232 ) : ( n20183 ) ;
assign n20185 =  ( n19788 ) ? ( bv_8_190_n250 ) : ( n20184 ) ;
assign n20186 =  ( n19786 ) ? ( bv_8_53_n436 ) : ( n20185 ) ;
assign n20187 =  ( n19784 ) ? ( bv_8_136_n425 ) : ( n20186 ) ;
assign n20188 =  ( n19782 ) ? ( bv_8_46_n429 ) : ( n20187 ) ;
assign n20189 =  ( n19780 ) ? ( bv_8_147_n392 ) : ( n20188 ) ;
assign n20190 =  ( n19778 ) ? ( bv_8_85_n423 ) : ( n20189 ) ;
assign n20191 =  ( n19776 ) ? ( bv_8_252_n15 ) : ( n20190 ) ;
assign n20192 =  ( n19774 ) ? ( bv_8_122_n416 ) : ( n20191 ) ;
assign n20193 =  ( n19772 ) ? ( bv_8_200_n213 ) : ( n20192 ) ;
assign n20194 =  ( n19770 ) ? ( bv_8_186_n263 ) : ( n20193 ) ;
assign n20195 =  ( n19768 ) ? ( bv_8_50_n408 ) : ( n20194 ) ;
assign n20196 =  ( n19766 ) ? ( bv_8_230_n103 ) : ( n20195 ) ;
assign n20197 =  ( n19764 ) ? ( bv_8_192_n242 ) : ( n20196 ) ;
assign n20198 =  ( n19762 ) ? ( bv_8_25_n399 ) : ( n20197 ) ;
assign n20199 =  ( n19760 ) ? ( bv_8_158_n355 ) : ( n20198 ) ;
assign n20200 =  ( n19758 ) ? ( bv_8_163_n339 ) : ( n20199 ) ;
assign n20201 =  ( n19756 ) ? ( bv_8_68_n390 ) : ( n20200 ) ;
assign n20202 =  ( n19754 ) ? ( bv_8_84_n386 ) : ( n20201 ) ;
assign n20203 =  ( n19752 ) ? ( bv_8_59_n382 ) : ( n20202 ) ;
assign n20204 =  ( n19750 ) ? ( bv_8_11_n379 ) : ( n20203 ) ;
assign n20205 =  ( n19748 ) ? ( bv_8_140_n376 ) : ( n20204 ) ;
assign n20206 =  ( n19746 ) ? ( bv_8_199_n216 ) : ( n20205 ) ;
assign n20207 =  ( n19744 ) ? ( bv_8_107_n370 ) : ( n20206 ) ;
assign n20208 =  ( n19742 ) ? ( bv_8_40_n366 ) : ( n20207 ) ;
assign n20209 =  ( n19740 ) ? ( bv_8_167_n325 ) : ( n20208 ) ;
assign n20210 =  ( n19738 ) ? ( bv_8_188_n257 ) : ( n20209 ) ;
assign n20211 =  ( n19736 ) ? ( bv_8_22_n357 ) : ( n20210 ) ;
assign n20212 =  ( n19734 ) ? ( bv_8_173_n307 ) : ( n20211 ) ;
assign n20213 =  ( n19732 ) ? ( bv_8_219_n146 ) : ( n20212 ) ;
assign n20214 =  ( n19730 ) ? ( bv_8_100_n348 ) : ( n20213 ) ;
assign n20215 =  ( n19728 ) ? ( bv_8_116_n345 ) : ( n20214 ) ;
assign n20216 =  ( n19726 ) ? ( bv_8_20_n341 ) : ( n20215 ) ;
assign n20217 =  ( n19724 ) ? ( bv_8_146_n337 ) : ( n20216 ) ;
assign n20218 =  ( n19722 ) ? ( bv_8_12_n333 ) : ( n20217 ) ;
assign n20219 =  ( n19720 ) ? ( bv_8_72_n330 ) : ( n20218 ) ;
assign n20220 =  ( n19718 ) ? ( bv_8_184_n270 ) : ( n20219 ) ;
assign n20221 =  ( n19716 ) ? ( bv_8_159_n323 ) : ( n20220 ) ;
assign n20222 =  ( n19714 ) ? ( bv_8_189_n254 ) : ( n20221 ) ;
assign n20223 =  ( n19712 ) ? ( bv_8_67_n318 ) : ( n20222 ) ;
assign n20224 =  ( n19710 ) ? ( bv_8_196_n228 ) : ( n20223 ) ;
assign n20225 =  ( n19708 ) ? ( bv_8_57_n312 ) : ( n20224 ) ;
assign n20226 =  ( n19706 ) ? ( bv_8_49_n309 ) : ( n20225 ) ;
assign n20227 =  ( n19704 ) ? ( bv_8_211_n175 ) : ( n20226 ) ;
assign n20228 =  ( n19702 ) ? ( bv_8_242_n55 ) : ( n20227 ) ;
assign n20229 =  ( n19700 ) ? ( bv_8_213_n167 ) : ( n20228 ) ;
assign n20230 =  ( n19698 ) ? ( bv_8_139_n297 ) : ( n20229 ) ;
assign n20231 =  ( n19696 ) ? ( bv_8_110_n294 ) : ( n20230 ) ;
assign n20232 =  ( n19694 ) ? ( bv_8_218_n150 ) : ( n20231 ) ;
assign n20233 =  ( n19692 ) ? ( bv_8_1_n287 ) : ( n20232 ) ;
assign n20234 =  ( n19690 ) ? ( bv_8_177_n283 ) : ( n20233 ) ;
assign n20235 =  ( n19688 ) ? ( bv_8_156_n279 ) : ( n20234 ) ;
assign n20236 =  ( n19686 ) ? ( bv_8_73_n275 ) : ( n20235 ) ;
assign n20237 =  ( n19684 ) ? ( bv_8_216_n157 ) : ( n20236 ) ;
assign n20238 =  ( n19682 ) ? ( bv_8_172_n268 ) : ( n20237 ) ;
assign n20239 =  ( n19680 ) ? ( bv_8_243_n51 ) : ( n20238 ) ;
assign n20240 =  ( n19678 ) ? ( bv_8_207_n188 ) : ( n20239 ) ;
assign n20241 =  ( n19676 ) ? ( bv_8_202_n207 ) : ( n20240 ) ;
assign n20242 =  ( n19674 ) ? ( bv_8_244_n47 ) : ( n20241 ) ;
assign n20243 =  ( n19672 ) ? ( bv_8_71_n252 ) : ( n20242 ) ;
assign n20244 =  ( n19670 ) ? ( bv_8_16_n248 ) : ( n20243 ) ;
assign n20245 =  ( n19668 ) ? ( bv_8_111_n244 ) : ( n20244 ) ;
assign n20246 =  ( n19666 ) ? ( bv_8_240_n63 ) : ( n20245 ) ;
assign n20247 =  ( n19664 ) ? ( bv_8_74_n237 ) : ( n20246 ) ;
assign n20248 =  ( n19662 ) ? ( bv_8_92_n234 ) : ( n20247 ) ;
assign n20249 =  ( n19660 ) ? ( bv_8_56_n230 ) : ( n20248 ) ;
assign n20250 =  ( n19658 ) ? ( bv_8_87_n226 ) : ( n20249 ) ;
assign n20251 =  ( n19656 ) ? ( bv_8_115_n222 ) : ( n20250 ) ;
assign n20252 =  ( n19654 ) ? ( bv_8_151_n218 ) : ( n20251 ) ;
assign n20253 =  ( n19652 ) ? ( bv_8_203_n203 ) : ( n20252 ) ;
assign n20254 =  ( n19650 ) ? ( bv_8_161_n211 ) : ( n20253 ) ;
assign n20255 =  ( n19648 ) ? ( bv_8_232_n95 ) : ( n20254 ) ;
assign n20256 =  ( n19646 ) ? ( bv_8_62_n205 ) : ( n20255 ) ;
assign n20257 =  ( n19644 ) ? ( bv_8_150_n201 ) : ( n20256 ) ;
assign n20258 =  ( n19642 ) ? ( bv_8_97_n198 ) : ( n20257 ) ;
assign n20259 =  ( n19640 ) ? ( bv_8_13_n194 ) : ( n20258 ) ;
assign n20260 =  ( n19638 ) ? ( bv_8_15_n190 ) : ( n20259 ) ;
assign n20261 =  ( n19636 ) ? ( bv_8_224_n126 ) : ( n20260 ) ;
assign n20262 =  ( n19634 ) ? ( bv_8_124_n184 ) : ( n20261 ) ;
assign n20263 =  ( n19632 ) ? ( bv_8_113_n180 ) : ( n20262 ) ;
assign n20264 =  ( n19630 ) ? ( bv_8_204_n177 ) : ( n20263 ) ;
assign n20265 =  ( n19628 ) ? ( bv_8_144_n173 ) : ( n20264 ) ;
assign n20266 =  ( n19626 ) ? ( bv_8_6_n169 ) : ( n20265 ) ;
assign n20267 =  ( n19624 ) ? ( bv_8_247_n35 ) : ( n20266 ) ;
assign n20268 =  ( n19622 ) ? ( bv_8_28_n162 ) : ( n20267 ) ;
assign n20269 =  ( n19620 ) ? ( bv_8_194_n159 ) : ( n20268 ) ;
assign n20270 =  ( n19618 ) ? ( bv_8_106_n155 ) : ( n20269 ) ;
assign n20271 =  ( n19616 ) ? ( bv_8_174_n152 ) : ( n20270 ) ;
assign n20272 =  ( n19614 ) ? ( bv_8_105_n148 ) : ( n20271 ) ;
assign n20273 =  ( n19612 ) ? ( bv_8_23_n144 ) : ( n20272 ) ;
assign n20274 =  ( n19610 ) ? ( bv_8_153_n140 ) : ( n20273 ) ;
assign n20275 =  ( n19608 ) ? ( bv_8_58_n136 ) : ( n20274 ) ;
assign n20276 =  ( n19606 ) ? ( bv_8_39_n132 ) : ( n20275 ) ;
assign n20277 =  ( n19604 ) ? ( bv_8_217_n128 ) : ( n20276 ) ;
assign n20278 =  ( n19602 ) ? ( bv_8_235_n83 ) : ( n20277 ) ;
assign n20279 =  ( n19600 ) ? ( bv_8_43_n121 ) : ( n20278 ) ;
assign n20280 =  ( n19598 ) ? ( bv_8_34_n117 ) : ( n20279 ) ;
assign n20281 =  ( n19596 ) ? ( bv_8_210_n113 ) : ( n20280 ) ;
assign n20282 =  ( n19594 ) ? ( bv_8_169_n109 ) : ( n20281 ) ;
assign n20283 =  ( n19592 ) ? ( bv_8_7_n105 ) : ( n20282 ) ;
assign n20284 =  ( n19590 ) ? ( bv_8_51_n101 ) : ( n20283 ) ;
assign n20285 =  ( n19588 ) ? ( bv_8_45_n97 ) : ( n20284 ) ;
assign n20286 =  ( n19586 ) ? ( bv_8_60_n93 ) : ( n20285 ) ;
assign n20287 =  ( n19584 ) ? ( bv_8_21_n89 ) : ( n20286 ) ;
assign n20288 =  ( n19582 ) ? ( bv_8_201_n85 ) : ( n20287 ) ;
assign n20289 =  ( n19580 ) ? ( bv_8_135_n81 ) : ( n20288 ) ;
assign n20290 =  ( n19578 ) ? ( bv_8_170_n77 ) : ( n20289 ) ;
assign n20291 =  ( n19576 ) ? ( bv_8_80_n73 ) : ( n20290 ) ;
assign n20292 =  ( n19574 ) ? ( bv_8_165_n69 ) : ( n20291 ) ;
assign n20293 =  ( n19572 ) ? ( bv_8_3_n65 ) : ( n20292 ) ;
assign n20294 =  ( n19570 ) ? ( bv_8_89_n61 ) : ( n20293 ) ;
assign n20295 =  ( n19568 ) ? ( bv_8_9_n57 ) : ( n20294 ) ;
assign n20296 =  ( n19566 ) ? ( bv_8_26_n53 ) : ( n20295 ) ;
assign n20297 =  ( n19564 ) ? ( bv_8_101_n49 ) : ( n20296 ) ;
assign n20298 =  ( n19562 ) ? ( bv_8_215_n45 ) : ( n20297 ) ;
assign n20299 =  ( n19560 ) ? ( bv_8_132_n41 ) : ( n20298 ) ;
assign n20300 =  ( n19558 ) ? ( bv_8_208_n37 ) : ( n20299 ) ;
assign n20301 =  ( n19556 ) ? ( bv_8_130_n33 ) : ( n20300 ) ;
assign n20302 =  ( n19554 ) ? ( bv_8_41_n29 ) : ( n20301 ) ;
assign n20303 =  ( n19552 ) ? ( bv_8_90_n25 ) : ( n20302 ) ;
assign n20304 =  ( n19550 ) ? ( bv_8_30_n21 ) : ( n20303 ) ;
assign n20305 =  ( n19548 ) ? ( bv_8_123_n17 ) : ( n20304 ) ;
assign n20306 =  ( n19546 ) ? ( bv_8_168_n13 ) : ( n20305 ) ;
assign n20307 =  ( n19544 ) ? ( bv_8_109_n9 ) : ( n20306 ) ;
assign n20308 =  ( n19542 ) ? ( bv_8_44_n5 ) : ( n20307 ) ;
assign n20309 =  ( n19540 ) ^ ( n20308 )  ;
assign n20310 = state_in[79:72] ;
assign n20311 =  ( n20310 ) == ( bv_8_255_n3 )  ;
assign n20312 = state_in[79:72] ;
assign n20313 =  ( n20312 ) == ( bv_8_254_n7 )  ;
assign n20314 = state_in[79:72] ;
assign n20315 =  ( n20314 ) == ( bv_8_253_n11 )  ;
assign n20316 = state_in[79:72] ;
assign n20317 =  ( n20316 ) == ( bv_8_252_n15 )  ;
assign n20318 = state_in[79:72] ;
assign n20319 =  ( n20318 ) == ( bv_8_251_n19 )  ;
assign n20320 = state_in[79:72] ;
assign n20321 =  ( n20320 ) == ( bv_8_250_n23 )  ;
assign n20322 = state_in[79:72] ;
assign n20323 =  ( n20322 ) == ( bv_8_249_n27 )  ;
assign n20324 = state_in[79:72] ;
assign n20325 =  ( n20324 ) == ( bv_8_248_n31 )  ;
assign n20326 = state_in[79:72] ;
assign n20327 =  ( n20326 ) == ( bv_8_247_n35 )  ;
assign n20328 = state_in[79:72] ;
assign n20329 =  ( n20328 ) == ( bv_8_246_n39 )  ;
assign n20330 = state_in[79:72] ;
assign n20331 =  ( n20330 ) == ( bv_8_245_n43 )  ;
assign n20332 = state_in[79:72] ;
assign n20333 =  ( n20332 ) == ( bv_8_244_n47 )  ;
assign n20334 = state_in[79:72] ;
assign n20335 =  ( n20334 ) == ( bv_8_243_n51 )  ;
assign n20336 = state_in[79:72] ;
assign n20337 =  ( n20336 ) == ( bv_8_242_n55 )  ;
assign n20338 = state_in[79:72] ;
assign n20339 =  ( n20338 ) == ( bv_8_241_n59 )  ;
assign n20340 = state_in[79:72] ;
assign n20341 =  ( n20340 ) == ( bv_8_240_n63 )  ;
assign n20342 = state_in[79:72] ;
assign n20343 =  ( n20342 ) == ( bv_8_239_n67 )  ;
assign n20344 = state_in[79:72] ;
assign n20345 =  ( n20344 ) == ( bv_8_238_n71 )  ;
assign n20346 = state_in[79:72] ;
assign n20347 =  ( n20346 ) == ( bv_8_237_n75 )  ;
assign n20348 = state_in[79:72] ;
assign n20349 =  ( n20348 ) == ( bv_8_236_n79 )  ;
assign n20350 = state_in[79:72] ;
assign n20351 =  ( n20350 ) == ( bv_8_235_n83 )  ;
assign n20352 = state_in[79:72] ;
assign n20353 =  ( n20352 ) == ( bv_8_234_n87 )  ;
assign n20354 = state_in[79:72] ;
assign n20355 =  ( n20354 ) == ( bv_8_233_n91 )  ;
assign n20356 = state_in[79:72] ;
assign n20357 =  ( n20356 ) == ( bv_8_232_n95 )  ;
assign n20358 = state_in[79:72] ;
assign n20359 =  ( n20358 ) == ( bv_8_231_n99 )  ;
assign n20360 = state_in[79:72] ;
assign n20361 =  ( n20360 ) == ( bv_8_230_n103 )  ;
assign n20362 = state_in[79:72] ;
assign n20363 =  ( n20362 ) == ( bv_8_229_n107 )  ;
assign n20364 = state_in[79:72] ;
assign n20365 =  ( n20364 ) == ( bv_8_228_n111 )  ;
assign n20366 = state_in[79:72] ;
assign n20367 =  ( n20366 ) == ( bv_8_227_n115 )  ;
assign n20368 = state_in[79:72] ;
assign n20369 =  ( n20368 ) == ( bv_8_226_n119 )  ;
assign n20370 = state_in[79:72] ;
assign n20371 =  ( n20370 ) == ( bv_8_225_n123 )  ;
assign n20372 = state_in[79:72] ;
assign n20373 =  ( n20372 ) == ( bv_8_224_n126 )  ;
assign n20374 = state_in[79:72] ;
assign n20375 =  ( n20374 ) == ( bv_8_223_n130 )  ;
assign n20376 = state_in[79:72] ;
assign n20377 =  ( n20376 ) == ( bv_8_222_n134 )  ;
assign n20378 = state_in[79:72] ;
assign n20379 =  ( n20378 ) == ( bv_8_221_n138 )  ;
assign n20380 = state_in[79:72] ;
assign n20381 =  ( n20380 ) == ( bv_8_220_n142 )  ;
assign n20382 = state_in[79:72] ;
assign n20383 =  ( n20382 ) == ( bv_8_219_n146 )  ;
assign n20384 = state_in[79:72] ;
assign n20385 =  ( n20384 ) == ( bv_8_218_n150 )  ;
assign n20386 = state_in[79:72] ;
assign n20387 =  ( n20386 ) == ( bv_8_217_n128 )  ;
assign n20388 = state_in[79:72] ;
assign n20389 =  ( n20388 ) == ( bv_8_216_n157 )  ;
assign n20390 = state_in[79:72] ;
assign n20391 =  ( n20390 ) == ( bv_8_215_n45 )  ;
assign n20392 = state_in[79:72] ;
assign n20393 =  ( n20392 ) == ( bv_8_214_n164 )  ;
assign n20394 = state_in[79:72] ;
assign n20395 =  ( n20394 ) == ( bv_8_213_n167 )  ;
assign n20396 = state_in[79:72] ;
assign n20397 =  ( n20396 ) == ( bv_8_212_n171 )  ;
assign n20398 = state_in[79:72] ;
assign n20399 =  ( n20398 ) == ( bv_8_211_n175 )  ;
assign n20400 = state_in[79:72] ;
assign n20401 =  ( n20400 ) == ( bv_8_210_n113 )  ;
assign n20402 = state_in[79:72] ;
assign n20403 =  ( n20402 ) == ( bv_8_209_n182 )  ;
assign n20404 = state_in[79:72] ;
assign n20405 =  ( n20404 ) == ( bv_8_208_n37 )  ;
assign n20406 = state_in[79:72] ;
assign n20407 =  ( n20406 ) == ( bv_8_207_n188 )  ;
assign n20408 = state_in[79:72] ;
assign n20409 =  ( n20408 ) == ( bv_8_206_n192 )  ;
assign n20410 = state_in[79:72] ;
assign n20411 =  ( n20410 ) == ( bv_8_205_n196 )  ;
assign n20412 = state_in[79:72] ;
assign n20413 =  ( n20412 ) == ( bv_8_204_n177 )  ;
assign n20414 = state_in[79:72] ;
assign n20415 =  ( n20414 ) == ( bv_8_203_n203 )  ;
assign n20416 = state_in[79:72] ;
assign n20417 =  ( n20416 ) == ( bv_8_202_n207 )  ;
assign n20418 = state_in[79:72] ;
assign n20419 =  ( n20418 ) == ( bv_8_201_n85 )  ;
assign n20420 = state_in[79:72] ;
assign n20421 =  ( n20420 ) == ( bv_8_200_n213 )  ;
assign n20422 = state_in[79:72] ;
assign n20423 =  ( n20422 ) == ( bv_8_199_n216 )  ;
assign n20424 = state_in[79:72] ;
assign n20425 =  ( n20424 ) == ( bv_8_198_n220 )  ;
assign n20426 = state_in[79:72] ;
assign n20427 =  ( n20426 ) == ( bv_8_197_n224 )  ;
assign n20428 = state_in[79:72] ;
assign n20429 =  ( n20428 ) == ( bv_8_196_n228 )  ;
assign n20430 = state_in[79:72] ;
assign n20431 =  ( n20430 ) == ( bv_8_195_n232 )  ;
assign n20432 = state_in[79:72] ;
assign n20433 =  ( n20432 ) == ( bv_8_194_n159 )  ;
assign n20434 = state_in[79:72] ;
assign n20435 =  ( n20434 ) == ( bv_8_193_n239 )  ;
assign n20436 = state_in[79:72] ;
assign n20437 =  ( n20436 ) == ( bv_8_192_n242 )  ;
assign n20438 = state_in[79:72] ;
assign n20439 =  ( n20438 ) == ( bv_8_191_n246 )  ;
assign n20440 = state_in[79:72] ;
assign n20441 =  ( n20440 ) == ( bv_8_190_n250 )  ;
assign n20442 = state_in[79:72] ;
assign n20443 =  ( n20442 ) == ( bv_8_189_n254 )  ;
assign n20444 = state_in[79:72] ;
assign n20445 =  ( n20444 ) == ( bv_8_188_n257 )  ;
assign n20446 = state_in[79:72] ;
assign n20447 =  ( n20446 ) == ( bv_8_187_n260 )  ;
assign n20448 = state_in[79:72] ;
assign n20449 =  ( n20448 ) == ( bv_8_186_n263 )  ;
assign n20450 = state_in[79:72] ;
assign n20451 =  ( n20450 ) == ( bv_8_185_n266 )  ;
assign n20452 = state_in[79:72] ;
assign n20453 =  ( n20452 ) == ( bv_8_184_n270 )  ;
assign n20454 = state_in[79:72] ;
assign n20455 =  ( n20454 ) == ( bv_8_183_n273 )  ;
assign n20456 = state_in[79:72] ;
assign n20457 =  ( n20456 ) == ( bv_8_182_n277 )  ;
assign n20458 = state_in[79:72] ;
assign n20459 =  ( n20458 ) == ( bv_8_181_n281 )  ;
assign n20460 = state_in[79:72] ;
assign n20461 =  ( n20460 ) == ( bv_8_180_n285 )  ;
assign n20462 = state_in[79:72] ;
assign n20463 =  ( n20462 ) == ( bv_8_179_n289 )  ;
assign n20464 = state_in[79:72] ;
assign n20465 =  ( n20464 ) == ( bv_8_178_n292 )  ;
assign n20466 = state_in[79:72] ;
assign n20467 =  ( n20466 ) == ( bv_8_177_n283 )  ;
assign n20468 = state_in[79:72] ;
assign n20469 =  ( n20468 ) == ( bv_8_176_n299 )  ;
assign n20470 = state_in[79:72] ;
assign n20471 =  ( n20470 ) == ( bv_8_175_n302 )  ;
assign n20472 = state_in[79:72] ;
assign n20473 =  ( n20472 ) == ( bv_8_174_n152 )  ;
assign n20474 = state_in[79:72] ;
assign n20475 =  ( n20474 ) == ( bv_8_173_n307 )  ;
assign n20476 = state_in[79:72] ;
assign n20477 =  ( n20476 ) == ( bv_8_172_n268 )  ;
assign n20478 = state_in[79:72] ;
assign n20479 =  ( n20478 ) == ( bv_8_171_n314 )  ;
assign n20480 = state_in[79:72] ;
assign n20481 =  ( n20480 ) == ( bv_8_170_n77 )  ;
assign n20482 = state_in[79:72] ;
assign n20483 =  ( n20482 ) == ( bv_8_169_n109 )  ;
assign n20484 = state_in[79:72] ;
assign n20485 =  ( n20484 ) == ( bv_8_168_n13 )  ;
assign n20486 = state_in[79:72] ;
assign n20487 =  ( n20486 ) == ( bv_8_167_n325 )  ;
assign n20488 = state_in[79:72] ;
assign n20489 =  ( n20488 ) == ( bv_8_166_n328 )  ;
assign n20490 = state_in[79:72] ;
assign n20491 =  ( n20490 ) == ( bv_8_165_n69 )  ;
assign n20492 = state_in[79:72] ;
assign n20493 =  ( n20492 ) == ( bv_8_164_n335 )  ;
assign n20494 = state_in[79:72] ;
assign n20495 =  ( n20494 ) == ( bv_8_163_n339 )  ;
assign n20496 = state_in[79:72] ;
assign n20497 =  ( n20496 ) == ( bv_8_162_n343 )  ;
assign n20498 = state_in[79:72] ;
assign n20499 =  ( n20498 ) == ( bv_8_161_n211 )  ;
assign n20500 = state_in[79:72] ;
assign n20501 =  ( n20500 ) == ( bv_8_160_n350 )  ;
assign n20502 = state_in[79:72] ;
assign n20503 =  ( n20502 ) == ( bv_8_159_n323 )  ;
assign n20504 = state_in[79:72] ;
assign n20505 =  ( n20504 ) == ( bv_8_158_n355 )  ;
assign n20506 = state_in[79:72] ;
assign n20507 =  ( n20506 ) == ( bv_8_157_n359 )  ;
assign n20508 = state_in[79:72] ;
assign n20509 =  ( n20508 ) == ( bv_8_156_n279 )  ;
assign n20510 = state_in[79:72] ;
assign n20511 =  ( n20510 ) == ( bv_8_155_n364 )  ;
assign n20512 = state_in[79:72] ;
assign n20513 =  ( n20512 ) == ( bv_8_154_n368 )  ;
assign n20514 = state_in[79:72] ;
assign n20515 =  ( n20514 ) == ( bv_8_153_n140 )  ;
assign n20516 = state_in[79:72] ;
assign n20517 =  ( n20516 ) == ( bv_8_152_n374 )  ;
assign n20518 = state_in[79:72] ;
assign n20519 =  ( n20518 ) == ( bv_8_151_n218 )  ;
assign n20520 = state_in[79:72] ;
assign n20521 =  ( n20520 ) == ( bv_8_150_n201 )  ;
assign n20522 = state_in[79:72] ;
assign n20523 =  ( n20522 ) == ( bv_8_149_n384 )  ;
assign n20524 = state_in[79:72] ;
assign n20525 =  ( n20524 ) == ( bv_8_148_n388 )  ;
assign n20526 = state_in[79:72] ;
assign n20527 =  ( n20526 ) == ( bv_8_147_n392 )  ;
assign n20528 = state_in[79:72] ;
assign n20529 =  ( n20528 ) == ( bv_8_146_n337 )  ;
assign n20530 = state_in[79:72] ;
assign n20531 =  ( n20530 ) == ( bv_8_145_n397 )  ;
assign n20532 = state_in[79:72] ;
assign n20533 =  ( n20532 ) == ( bv_8_144_n173 )  ;
assign n20534 = state_in[79:72] ;
assign n20535 =  ( n20534 ) == ( bv_8_143_n403 )  ;
assign n20536 = state_in[79:72] ;
assign n20537 =  ( n20536 ) == ( bv_8_142_n406 )  ;
assign n20538 = state_in[79:72] ;
assign n20539 =  ( n20538 ) == ( bv_8_141_n410 )  ;
assign n20540 = state_in[79:72] ;
assign n20541 =  ( n20540 ) == ( bv_8_140_n376 )  ;
assign n20542 = state_in[79:72] ;
assign n20543 =  ( n20542 ) == ( bv_8_139_n297 )  ;
assign n20544 = state_in[79:72] ;
assign n20545 =  ( n20544 ) == ( bv_8_138_n418 )  ;
assign n20546 = state_in[79:72] ;
assign n20547 =  ( n20546 ) == ( bv_8_137_n421 )  ;
assign n20548 = state_in[79:72] ;
assign n20549 =  ( n20548 ) == ( bv_8_136_n425 )  ;
assign n20550 = state_in[79:72] ;
assign n20551 =  ( n20550 ) == ( bv_8_135_n81 )  ;
assign n20552 = state_in[79:72] ;
assign n20553 =  ( n20552 ) == ( bv_8_134_n431 )  ;
assign n20554 = state_in[79:72] ;
assign n20555 =  ( n20554 ) == ( bv_8_133_n434 )  ;
assign n20556 = state_in[79:72] ;
assign n20557 =  ( n20556 ) == ( bv_8_132_n41 )  ;
assign n20558 = state_in[79:72] ;
assign n20559 =  ( n20558 ) == ( bv_8_131_n440 )  ;
assign n20560 = state_in[79:72] ;
assign n20561 =  ( n20560 ) == ( bv_8_130_n33 )  ;
assign n20562 = state_in[79:72] ;
assign n20563 =  ( n20562 ) == ( bv_8_129_n446 )  ;
assign n20564 = state_in[79:72] ;
assign n20565 =  ( n20564 ) == ( bv_8_128_n450 )  ;
assign n20566 = state_in[79:72] ;
assign n20567 =  ( n20566 ) == ( bv_8_127_n453 )  ;
assign n20568 = state_in[79:72] ;
assign n20569 =  ( n20568 ) == ( bv_8_126_n456 )  ;
assign n20570 = state_in[79:72] ;
assign n20571 =  ( n20570 ) == ( bv_8_125_n459 )  ;
assign n20572 = state_in[79:72] ;
assign n20573 =  ( n20572 ) == ( bv_8_124_n184 )  ;
assign n20574 = state_in[79:72] ;
assign n20575 =  ( n20574 ) == ( bv_8_123_n17 )  ;
assign n20576 = state_in[79:72] ;
assign n20577 =  ( n20576 ) == ( bv_8_122_n416 )  ;
assign n20578 = state_in[79:72] ;
assign n20579 =  ( n20578 ) == ( bv_8_121_n470 )  ;
assign n20580 = state_in[79:72] ;
assign n20581 =  ( n20580 ) == ( bv_8_120_n474 )  ;
assign n20582 = state_in[79:72] ;
assign n20583 =  ( n20582 ) == ( bv_8_119_n472 )  ;
assign n20584 = state_in[79:72] ;
assign n20585 =  ( n20584 ) == ( bv_8_118_n480 )  ;
assign n20586 = state_in[79:72] ;
assign n20587 =  ( n20586 ) == ( bv_8_117_n484 )  ;
assign n20588 = state_in[79:72] ;
assign n20589 =  ( n20588 ) == ( bv_8_116_n345 )  ;
assign n20590 = state_in[79:72] ;
assign n20591 =  ( n20590 ) == ( bv_8_115_n222 )  ;
assign n20592 = state_in[79:72] ;
assign n20593 =  ( n20592 ) == ( bv_8_114_n494 )  ;
assign n20594 = state_in[79:72] ;
assign n20595 =  ( n20594 ) == ( bv_8_113_n180 )  ;
assign n20596 = state_in[79:72] ;
assign n20597 =  ( n20596 ) == ( bv_8_112_n482 )  ;
assign n20598 = state_in[79:72] ;
assign n20599 =  ( n20598 ) == ( bv_8_111_n244 )  ;
assign n20600 = state_in[79:72] ;
assign n20601 =  ( n20600 ) == ( bv_8_110_n294 )  ;
assign n20602 = state_in[79:72] ;
assign n20603 =  ( n20602 ) == ( bv_8_109_n9 )  ;
assign n20604 = state_in[79:72] ;
assign n20605 =  ( n20604 ) == ( bv_8_108_n510 )  ;
assign n20606 = state_in[79:72] ;
assign n20607 =  ( n20606 ) == ( bv_8_107_n370 )  ;
assign n20608 = state_in[79:72] ;
assign n20609 =  ( n20608 ) == ( bv_8_106_n155 )  ;
assign n20610 = state_in[79:72] ;
assign n20611 =  ( n20610 ) == ( bv_8_105_n148 )  ;
assign n20612 = state_in[79:72] ;
assign n20613 =  ( n20612 ) == ( bv_8_104_n520 )  ;
assign n20614 = state_in[79:72] ;
assign n20615 =  ( n20614 ) == ( bv_8_103_n523 )  ;
assign n20616 = state_in[79:72] ;
assign n20617 =  ( n20616 ) == ( bv_8_102_n527 )  ;
assign n20618 = state_in[79:72] ;
assign n20619 =  ( n20618 ) == ( bv_8_101_n49 )  ;
assign n20620 = state_in[79:72] ;
assign n20621 =  ( n20620 ) == ( bv_8_100_n348 )  ;
assign n20622 = state_in[79:72] ;
assign n20623 =  ( n20622 ) == ( bv_8_99_n476 )  ;
assign n20624 = state_in[79:72] ;
assign n20625 =  ( n20624 ) == ( bv_8_98_n536 )  ;
assign n20626 = state_in[79:72] ;
assign n20627 =  ( n20626 ) == ( bv_8_97_n198 )  ;
assign n20628 = state_in[79:72] ;
assign n20629 =  ( n20628 ) == ( bv_8_96_n542 )  ;
assign n20630 = state_in[79:72] ;
assign n20631 =  ( n20630 ) == ( bv_8_95_n545 )  ;
assign n20632 = state_in[79:72] ;
assign n20633 =  ( n20632 ) == ( bv_8_94_n548 )  ;
assign n20634 = state_in[79:72] ;
assign n20635 =  ( n20634 ) == ( bv_8_93_n498 )  ;
assign n20636 = state_in[79:72] ;
assign n20637 =  ( n20636 ) == ( bv_8_92_n234 )  ;
assign n20638 = state_in[79:72] ;
assign n20639 =  ( n20638 ) == ( bv_8_91_n555 )  ;
assign n20640 = state_in[79:72] ;
assign n20641 =  ( n20640 ) == ( bv_8_90_n25 )  ;
assign n20642 = state_in[79:72] ;
assign n20643 =  ( n20642 ) == ( bv_8_89_n61 )  ;
assign n20644 = state_in[79:72] ;
assign n20645 =  ( n20644 ) == ( bv_8_88_n562 )  ;
assign n20646 = state_in[79:72] ;
assign n20647 =  ( n20646 ) == ( bv_8_87_n226 )  ;
assign n20648 = state_in[79:72] ;
assign n20649 =  ( n20648 ) == ( bv_8_86_n567 )  ;
assign n20650 = state_in[79:72] ;
assign n20651 =  ( n20650 ) == ( bv_8_85_n423 )  ;
assign n20652 = state_in[79:72] ;
assign n20653 =  ( n20652 ) == ( bv_8_84_n386 )  ;
assign n20654 = state_in[79:72] ;
assign n20655 =  ( n20654 ) == ( bv_8_83_n575 )  ;
assign n20656 = state_in[79:72] ;
assign n20657 =  ( n20656 ) == ( bv_8_82_n578 )  ;
assign n20658 = state_in[79:72] ;
assign n20659 =  ( n20658 ) == ( bv_8_81_n582 )  ;
assign n20660 = state_in[79:72] ;
assign n20661 =  ( n20660 ) == ( bv_8_80_n73 )  ;
assign n20662 = state_in[79:72] ;
assign n20663 =  ( n20662 ) == ( bv_8_79_n538 )  ;
assign n20664 = state_in[79:72] ;
assign n20665 =  ( n20664 ) == ( bv_8_78_n590 )  ;
assign n20666 = state_in[79:72] ;
assign n20667 =  ( n20666 ) == ( bv_8_77_n593 )  ;
assign n20668 = state_in[79:72] ;
assign n20669 =  ( n20668 ) == ( bv_8_76_n596 )  ;
assign n20670 = state_in[79:72] ;
assign n20671 =  ( n20670 ) == ( bv_8_75_n503 )  ;
assign n20672 = state_in[79:72] ;
assign n20673 =  ( n20672 ) == ( bv_8_74_n237 )  ;
assign n20674 = state_in[79:72] ;
assign n20675 =  ( n20674 ) == ( bv_8_73_n275 )  ;
assign n20676 = state_in[79:72] ;
assign n20677 =  ( n20676 ) == ( bv_8_72_n330 )  ;
assign n20678 = state_in[79:72] ;
assign n20679 =  ( n20678 ) == ( bv_8_71_n252 )  ;
assign n20680 = state_in[79:72] ;
assign n20681 =  ( n20680 ) == ( bv_8_70_n609 )  ;
assign n20682 = state_in[79:72] ;
assign n20683 =  ( n20682 ) == ( bv_8_69_n612 )  ;
assign n20684 = state_in[79:72] ;
assign n20685 =  ( n20684 ) == ( bv_8_68_n390 )  ;
assign n20686 = state_in[79:72] ;
assign n20687 =  ( n20686 ) == ( bv_8_67_n318 )  ;
assign n20688 = state_in[79:72] ;
assign n20689 =  ( n20688 ) == ( bv_8_66_n466 )  ;
assign n20690 = state_in[79:72] ;
assign n20691 =  ( n20690 ) == ( bv_8_65_n623 )  ;
assign n20692 = state_in[79:72] ;
assign n20693 =  ( n20692 ) == ( bv_8_64_n573 )  ;
assign n20694 = state_in[79:72] ;
assign n20695 =  ( n20694 ) == ( bv_8_63_n489 )  ;
assign n20696 = state_in[79:72] ;
assign n20697 =  ( n20696 ) == ( bv_8_62_n205 )  ;
assign n20698 = state_in[79:72] ;
assign n20699 =  ( n20698 ) == ( bv_8_61_n634 )  ;
assign n20700 = state_in[79:72] ;
assign n20701 =  ( n20700 ) == ( bv_8_60_n93 )  ;
assign n20702 = state_in[79:72] ;
assign n20703 =  ( n20702 ) == ( bv_8_59_n382 )  ;
assign n20704 = state_in[79:72] ;
assign n20705 =  ( n20704 ) == ( bv_8_58_n136 )  ;
assign n20706 = state_in[79:72] ;
assign n20707 =  ( n20706 ) == ( bv_8_57_n312 )  ;
assign n20708 = state_in[79:72] ;
assign n20709 =  ( n20708 ) == ( bv_8_56_n230 )  ;
assign n20710 = state_in[79:72] ;
assign n20711 =  ( n20710 ) == ( bv_8_55_n650 )  ;
assign n20712 = state_in[79:72] ;
assign n20713 =  ( n20712 ) == ( bv_8_54_n616 )  ;
assign n20714 = state_in[79:72] ;
assign n20715 =  ( n20714 ) == ( bv_8_53_n436 )  ;
assign n20716 = state_in[79:72] ;
assign n20717 =  ( n20716 ) == ( bv_8_52_n619 )  ;
assign n20718 = state_in[79:72] ;
assign n20719 =  ( n20718 ) == ( bv_8_51_n101 )  ;
assign n20720 = state_in[79:72] ;
assign n20721 =  ( n20720 ) == ( bv_8_50_n408 )  ;
assign n20722 = state_in[79:72] ;
assign n20723 =  ( n20722 ) == ( bv_8_49_n309 )  ;
assign n20724 = state_in[79:72] ;
assign n20725 =  ( n20724 ) == ( bv_8_48_n660 )  ;
assign n20726 = state_in[79:72] ;
assign n20727 =  ( n20726 ) == ( bv_8_47_n652 )  ;
assign n20728 = state_in[79:72] ;
assign n20729 =  ( n20728 ) == ( bv_8_46_n429 )  ;
assign n20730 = state_in[79:72] ;
assign n20731 =  ( n20730 ) == ( bv_8_45_n97 )  ;
assign n20732 = state_in[79:72] ;
assign n20733 =  ( n20732 ) == ( bv_8_44_n5 )  ;
assign n20734 = state_in[79:72] ;
assign n20735 =  ( n20734 ) == ( bv_8_43_n121 )  ;
assign n20736 = state_in[79:72] ;
assign n20737 =  ( n20736 ) == ( bv_8_42_n672 )  ;
assign n20738 = state_in[79:72] ;
assign n20739 =  ( n20738 ) == ( bv_8_41_n29 )  ;
assign n20740 = state_in[79:72] ;
assign n20741 =  ( n20740 ) == ( bv_8_40_n366 )  ;
assign n20742 = state_in[79:72] ;
assign n20743 =  ( n20742 ) == ( bv_8_39_n132 )  ;
assign n20744 = state_in[79:72] ;
assign n20745 =  ( n20744 ) == ( bv_8_38_n444 )  ;
assign n20746 = state_in[79:72] ;
assign n20747 =  ( n20746 ) == ( bv_8_37_n506 )  ;
assign n20748 = state_in[79:72] ;
assign n20749 =  ( n20748 ) == ( bv_8_36_n645 )  ;
assign n20750 = state_in[79:72] ;
assign n20751 =  ( n20750 ) == ( bv_8_35_n696 )  ;
assign n20752 = state_in[79:72] ;
assign n20753 =  ( n20752 ) == ( bv_8_34_n117 )  ;
assign n20754 = state_in[79:72] ;
assign n20755 =  ( n20754 ) == ( bv_8_33_n486 )  ;
assign n20756 = state_in[79:72] ;
assign n20757 =  ( n20756 ) == ( bv_8_32_n463 )  ;
assign n20758 = state_in[79:72] ;
assign n20759 =  ( n20758 ) == ( bv_8_31_n705 )  ;
assign n20760 = state_in[79:72] ;
assign n20761 =  ( n20760 ) == ( bv_8_30_n21 )  ;
assign n20762 = state_in[79:72] ;
assign n20763 =  ( n20762 ) == ( bv_8_29_n625 )  ;
assign n20764 = state_in[79:72] ;
assign n20765 =  ( n20764 ) == ( bv_8_28_n162 )  ;
assign n20766 = state_in[79:72] ;
assign n20767 =  ( n20766 ) == ( bv_8_27_n642 )  ;
assign n20768 = state_in[79:72] ;
assign n20769 =  ( n20768 ) == ( bv_8_26_n53 )  ;
assign n20770 = state_in[79:72] ;
assign n20771 =  ( n20770 ) == ( bv_8_25_n399 )  ;
assign n20772 = state_in[79:72] ;
assign n20773 =  ( n20772 ) == ( bv_8_24_n448 )  ;
assign n20774 = state_in[79:72] ;
assign n20775 =  ( n20774 ) == ( bv_8_23_n144 )  ;
assign n20776 = state_in[79:72] ;
assign n20777 =  ( n20776 ) == ( bv_8_22_n357 )  ;
assign n20778 = state_in[79:72] ;
assign n20779 =  ( n20778 ) == ( bv_8_21_n89 )  ;
assign n20780 = state_in[79:72] ;
assign n20781 =  ( n20780 ) == ( bv_8_20_n341 )  ;
assign n20782 = state_in[79:72] ;
assign n20783 =  ( n20782 ) == ( bv_8_19_n588 )  ;
assign n20784 = state_in[79:72] ;
assign n20785 =  ( n20784 ) == ( bv_8_18_n628 )  ;
assign n20786 = state_in[79:72] ;
assign n20787 =  ( n20786 ) == ( bv_8_17_n525 )  ;
assign n20788 = state_in[79:72] ;
assign n20789 =  ( n20788 ) == ( bv_8_16_n248 )  ;
assign n20790 = state_in[79:72] ;
assign n20791 =  ( n20790 ) == ( bv_8_15_n190 )  ;
assign n20792 = state_in[79:72] ;
assign n20793 =  ( n20792 ) == ( bv_8_14_n648 )  ;
assign n20794 = state_in[79:72] ;
assign n20795 =  ( n20794 ) == ( bv_8_13_n194 )  ;
assign n20796 = state_in[79:72] ;
assign n20797 =  ( n20796 ) == ( bv_8_12_n333 )  ;
assign n20798 = state_in[79:72] ;
assign n20799 =  ( n20798 ) == ( bv_8_11_n379 )  ;
assign n20800 = state_in[79:72] ;
assign n20801 =  ( n20800 ) == ( bv_8_10_n655 )  ;
assign n20802 = state_in[79:72] ;
assign n20803 =  ( n20802 ) == ( bv_8_9_n57 )  ;
assign n20804 = state_in[79:72] ;
assign n20805 =  ( n20804 ) == ( bv_8_8_n669 )  ;
assign n20806 = state_in[79:72] ;
assign n20807 =  ( n20806 ) == ( bv_8_7_n105 )  ;
assign n20808 = state_in[79:72] ;
assign n20809 =  ( n20808 ) == ( bv_8_6_n169 )  ;
assign n20810 = state_in[79:72] ;
assign n20811 =  ( n20810 ) == ( bv_8_5_n492 )  ;
assign n20812 = state_in[79:72] ;
assign n20813 =  ( n20812 ) == ( bv_8_4_n516 )  ;
assign n20814 = state_in[79:72] ;
assign n20815 =  ( n20814 ) == ( bv_8_3_n65 )  ;
assign n20816 = state_in[79:72] ;
assign n20817 =  ( n20816 ) == ( bv_8_2_n751 )  ;
assign n20818 = state_in[79:72] ;
assign n20819 =  ( n20818 ) == ( bv_8_1_n287 )  ;
assign n20820 = state_in[79:72] ;
assign n20821 =  ( n20820 ) == ( bv_8_0_n580 )  ;
assign n20822 =  ( n20821 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n20823 =  ( n20819 ) ? ( bv_8_124_n184 ) : ( n20822 ) ;
assign n20824 =  ( n20817 ) ? ( bv_8_119_n472 ) : ( n20823 ) ;
assign n20825 =  ( n20815 ) ? ( bv_8_123_n17 ) : ( n20824 ) ;
assign n20826 =  ( n20813 ) ? ( bv_8_242_n55 ) : ( n20825 ) ;
assign n20827 =  ( n20811 ) ? ( bv_8_107_n370 ) : ( n20826 ) ;
assign n20828 =  ( n20809 ) ? ( bv_8_111_n244 ) : ( n20827 ) ;
assign n20829 =  ( n20807 ) ? ( bv_8_197_n224 ) : ( n20828 ) ;
assign n20830 =  ( n20805 ) ? ( bv_8_48_n660 ) : ( n20829 ) ;
assign n20831 =  ( n20803 ) ? ( bv_8_1_n287 ) : ( n20830 ) ;
assign n20832 =  ( n20801 ) ? ( bv_8_103_n523 ) : ( n20831 ) ;
assign n20833 =  ( n20799 ) ? ( bv_8_43_n121 ) : ( n20832 ) ;
assign n20834 =  ( n20797 ) ? ( bv_8_254_n7 ) : ( n20833 ) ;
assign n20835 =  ( n20795 ) ? ( bv_8_215_n45 ) : ( n20834 ) ;
assign n20836 =  ( n20793 ) ? ( bv_8_171_n314 ) : ( n20835 ) ;
assign n20837 =  ( n20791 ) ? ( bv_8_118_n480 ) : ( n20836 ) ;
assign n20838 =  ( n20789 ) ? ( bv_8_202_n207 ) : ( n20837 ) ;
assign n20839 =  ( n20787 ) ? ( bv_8_130_n33 ) : ( n20838 ) ;
assign n20840 =  ( n20785 ) ? ( bv_8_201_n85 ) : ( n20839 ) ;
assign n20841 =  ( n20783 ) ? ( bv_8_125_n459 ) : ( n20840 ) ;
assign n20842 =  ( n20781 ) ? ( bv_8_250_n23 ) : ( n20841 ) ;
assign n20843 =  ( n20779 ) ? ( bv_8_89_n61 ) : ( n20842 ) ;
assign n20844 =  ( n20777 ) ? ( bv_8_71_n252 ) : ( n20843 ) ;
assign n20845 =  ( n20775 ) ? ( bv_8_240_n63 ) : ( n20844 ) ;
assign n20846 =  ( n20773 ) ? ( bv_8_173_n307 ) : ( n20845 ) ;
assign n20847 =  ( n20771 ) ? ( bv_8_212_n171 ) : ( n20846 ) ;
assign n20848 =  ( n20769 ) ? ( bv_8_162_n343 ) : ( n20847 ) ;
assign n20849 =  ( n20767 ) ? ( bv_8_175_n302 ) : ( n20848 ) ;
assign n20850 =  ( n20765 ) ? ( bv_8_156_n279 ) : ( n20849 ) ;
assign n20851 =  ( n20763 ) ? ( bv_8_164_n335 ) : ( n20850 ) ;
assign n20852 =  ( n20761 ) ? ( bv_8_114_n494 ) : ( n20851 ) ;
assign n20853 =  ( n20759 ) ? ( bv_8_192_n242 ) : ( n20852 ) ;
assign n20854 =  ( n20757 ) ? ( bv_8_183_n273 ) : ( n20853 ) ;
assign n20855 =  ( n20755 ) ? ( bv_8_253_n11 ) : ( n20854 ) ;
assign n20856 =  ( n20753 ) ? ( bv_8_147_n392 ) : ( n20855 ) ;
assign n20857 =  ( n20751 ) ? ( bv_8_38_n444 ) : ( n20856 ) ;
assign n20858 =  ( n20749 ) ? ( bv_8_54_n616 ) : ( n20857 ) ;
assign n20859 =  ( n20747 ) ? ( bv_8_63_n489 ) : ( n20858 ) ;
assign n20860 =  ( n20745 ) ? ( bv_8_247_n35 ) : ( n20859 ) ;
assign n20861 =  ( n20743 ) ? ( bv_8_204_n177 ) : ( n20860 ) ;
assign n20862 =  ( n20741 ) ? ( bv_8_52_n619 ) : ( n20861 ) ;
assign n20863 =  ( n20739 ) ? ( bv_8_165_n69 ) : ( n20862 ) ;
assign n20864 =  ( n20737 ) ? ( bv_8_229_n107 ) : ( n20863 ) ;
assign n20865 =  ( n20735 ) ? ( bv_8_241_n59 ) : ( n20864 ) ;
assign n20866 =  ( n20733 ) ? ( bv_8_113_n180 ) : ( n20865 ) ;
assign n20867 =  ( n20731 ) ? ( bv_8_216_n157 ) : ( n20866 ) ;
assign n20868 =  ( n20729 ) ? ( bv_8_49_n309 ) : ( n20867 ) ;
assign n20869 =  ( n20727 ) ? ( bv_8_21_n89 ) : ( n20868 ) ;
assign n20870 =  ( n20725 ) ? ( bv_8_4_n516 ) : ( n20869 ) ;
assign n20871 =  ( n20723 ) ? ( bv_8_199_n216 ) : ( n20870 ) ;
assign n20872 =  ( n20721 ) ? ( bv_8_35_n696 ) : ( n20871 ) ;
assign n20873 =  ( n20719 ) ? ( bv_8_195_n232 ) : ( n20872 ) ;
assign n20874 =  ( n20717 ) ? ( bv_8_24_n448 ) : ( n20873 ) ;
assign n20875 =  ( n20715 ) ? ( bv_8_150_n201 ) : ( n20874 ) ;
assign n20876 =  ( n20713 ) ? ( bv_8_5_n492 ) : ( n20875 ) ;
assign n20877 =  ( n20711 ) ? ( bv_8_154_n368 ) : ( n20876 ) ;
assign n20878 =  ( n20709 ) ? ( bv_8_7_n105 ) : ( n20877 ) ;
assign n20879 =  ( n20707 ) ? ( bv_8_18_n628 ) : ( n20878 ) ;
assign n20880 =  ( n20705 ) ? ( bv_8_128_n450 ) : ( n20879 ) ;
assign n20881 =  ( n20703 ) ? ( bv_8_226_n119 ) : ( n20880 ) ;
assign n20882 =  ( n20701 ) ? ( bv_8_235_n83 ) : ( n20881 ) ;
assign n20883 =  ( n20699 ) ? ( bv_8_39_n132 ) : ( n20882 ) ;
assign n20884 =  ( n20697 ) ? ( bv_8_178_n292 ) : ( n20883 ) ;
assign n20885 =  ( n20695 ) ? ( bv_8_117_n484 ) : ( n20884 ) ;
assign n20886 =  ( n20693 ) ? ( bv_8_9_n57 ) : ( n20885 ) ;
assign n20887 =  ( n20691 ) ? ( bv_8_131_n440 ) : ( n20886 ) ;
assign n20888 =  ( n20689 ) ? ( bv_8_44_n5 ) : ( n20887 ) ;
assign n20889 =  ( n20687 ) ? ( bv_8_26_n53 ) : ( n20888 ) ;
assign n20890 =  ( n20685 ) ? ( bv_8_27_n642 ) : ( n20889 ) ;
assign n20891 =  ( n20683 ) ? ( bv_8_110_n294 ) : ( n20890 ) ;
assign n20892 =  ( n20681 ) ? ( bv_8_90_n25 ) : ( n20891 ) ;
assign n20893 =  ( n20679 ) ? ( bv_8_160_n350 ) : ( n20892 ) ;
assign n20894 =  ( n20677 ) ? ( bv_8_82_n578 ) : ( n20893 ) ;
assign n20895 =  ( n20675 ) ? ( bv_8_59_n382 ) : ( n20894 ) ;
assign n20896 =  ( n20673 ) ? ( bv_8_214_n164 ) : ( n20895 ) ;
assign n20897 =  ( n20671 ) ? ( bv_8_179_n289 ) : ( n20896 ) ;
assign n20898 =  ( n20669 ) ? ( bv_8_41_n29 ) : ( n20897 ) ;
assign n20899 =  ( n20667 ) ? ( bv_8_227_n115 ) : ( n20898 ) ;
assign n20900 =  ( n20665 ) ? ( bv_8_47_n652 ) : ( n20899 ) ;
assign n20901 =  ( n20663 ) ? ( bv_8_132_n41 ) : ( n20900 ) ;
assign n20902 =  ( n20661 ) ? ( bv_8_83_n575 ) : ( n20901 ) ;
assign n20903 =  ( n20659 ) ? ( bv_8_209_n182 ) : ( n20902 ) ;
assign n20904 =  ( n20657 ) ? ( bv_8_0_n580 ) : ( n20903 ) ;
assign n20905 =  ( n20655 ) ? ( bv_8_237_n75 ) : ( n20904 ) ;
assign n20906 =  ( n20653 ) ? ( bv_8_32_n463 ) : ( n20905 ) ;
assign n20907 =  ( n20651 ) ? ( bv_8_252_n15 ) : ( n20906 ) ;
assign n20908 =  ( n20649 ) ? ( bv_8_177_n283 ) : ( n20907 ) ;
assign n20909 =  ( n20647 ) ? ( bv_8_91_n555 ) : ( n20908 ) ;
assign n20910 =  ( n20645 ) ? ( bv_8_106_n155 ) : ( n20909 ) ;
assign n20911 =  ( n20643 ) ? ( bv_8_203_n203 ) : ( n20910 ) ;
assign n20912 =  ( n20641 ) ? ( bv_8_190_n250 ) : ( n20911 ) ;
assign n20913 =  ( n20639 ) ? ( bv_8_57_n312 ) : ( n20912 ) ;
assign n20914 =  ( n20637 ) ? ( bv_8_74_n237 ) : ( n20913 ) ;
assign n20915 =  ( n20635 ) ? ( bv_8_76_n596 ) : ( n20914 ) ;
assign n20916 =  ( n20633 ) ? ( bv_8_88_n562 ) : ( n20915 ) ;
assign n20917 =  ( n20631 ) ? ( bv_8_207_n188 ) : ( n20916 ) ;
assign n20918 =  ( n20629 ) ? ( bv_8_208_n37 ) : ( n20917 ) ;
assign n20919 =  ( n20627 ) ? ( bv_8_239_n67 ) : ( n20918 ) ;
assign n20920 =  ( n20625 ) ? ( bv_8_170_n77 ) : ( n20919 ) ;
assign n20921 =  ( n20623 ) ? ( bv_8_251_n19 ) : ( n20920 ) ;
assign n20922 =  ( n20621 ) ? ( bv_8_67_n318 ) : ( n20921 ) ;
assign n20923 =  ( n20619 ) ? ( bv_8_77_n593 ) : ( n20922 ) ;
assign n20924 =  ( n20617 ) ? ( bv_8_51_n101 ) : ( n20923 ) ;
assign n20925 =  ( n20615 ) ? ( bv_8_133_n434 ) : ( n20924 ) ;
assign n20926 =  ( n20613 ) ? ( bv_8_69_n612 ) : ( n20925 ) ;
assign n20927 =  ( n20611 ) ? ( bv_8_249_n27 ) : ( n20926 ) ;
assign n20928 =  ( n20609 ) ? ( bv_8_2_n751 ) : ( n20927 ) ;
assign n20929 =  ( n20607 ) ? ( bv_8_127_n453 ) : ( n20928 ) ;
assign n20930 =  ( n20605 ) ? ( bv_8_80_n73 ) : ( n20929 ) ;
assign n20931 =  ( n20603 ) ? ( bv_8_60_n93 ) : ( n20930 ) ;
assign n20932 =  ( n20601 ) ? ( bv_8_159_n323 ) : ( n20931 ) ;
assign n20933 =  ( n20599 ) ? ( bv_8_168_n13 ) : ( n20932 ) ;
assign n20934 =  ( n20597 ) ? ( bv_8_81_n582 ) : ( n20933 ) ;
assign n20935 =  ( n20595 ) ? ( bv_8_163_n339 ) : ( n20934 ) ;
assign n20936 =  ( n20593 ) ? ( bv_8_64_n573 ) : ( n20935 ) ;
assign n20937 =  ( n20591 ) ? ( bv_8_143_n403 ) : ( n20936 ) ;
assign n20938 =  ( n20589 ) ? ( bv_8_146_n337 ) : ( n20937 ) ;
assign n20939 =  ( n20587 ) ? ( bv_8_157_n359 ) : ( n20938 ) ;
assign n20940 =  ( n20585 ) ? ( bv_8_56_n230 ) : ( n20939 ) ;
assign n20941 =  ( n20583 ) ? ( bv_8_245_n43 ) : ( n20940 ) ;
assign n20942 =  ( n20581 ) ? ( bv_8_188_n257 ) : ( n20941 ) ;
assign n20943 =  ( n20579 ) ? ( bv_8_182_n277 ) : ( n20942 ) ;
assign n20944 =  ( n20577 ) ? ( bv_8_218_n150 ) : ( n20943 ) ;
assign n20945 =  ( n20575 ) ? ( bv_8_33_n486 ) : ( n20944 ) ;
assign n20946 =  ( n20573 ) ? ( bv_8_16_n248 ) : ( n20945 ) ;
assign n20947 =  ( n20571 ) ? ( bv_8_255_n3 ) : ( n20946 ) ;
assign n20948 =  ( n20569 ) ? ( bv_8_243_n51 ) : ( n20947 ) ;
assign n20949 =  ( n20567 ) ? ( bv_8_210_n113 ) : ( n20948 ) ;
assign n20950 =  ( n20565 ) ? ( bv_8_205_n196 ) : ( n20949 ) ;
assign n20951 =  ( n20563 ) ? ( bv_8_12_n333 ) : ( n20950 ) ;
assign n20952 =  ( n20561 ) ? ( bv_8_19_n588 ) : ( n20951 ) ;
assign n20953 =  ( n20559 ) ? ( bv_8_236_n79 ) : ( n20952 ) ;
assign n20954 =  ( n20557 ) ? ( bv_8_95_n545 ) : ( n20953 ) ;
assign n20955 =  ( n20555 ) ? ( bv_8_151_n218 ) : ( n20954 ) ;
assign n20956 =  ( n20553 ) ? ( bv_8_68_n390 ) : ( n20955 ) ;
assign n20957 =  ( n20551 ) ? ( bv_8_23_n144 ) : ( n20956 ) ;
assign n20958 =  ( n20549 ) ? ( bv_8_196_n228 ) : ( n20957 ) ;
assign n20959 =  ( n20547 ) ? ( bv_8_167_n325 ) : ( n20958 ) ;
assign n20960 =  ( n20545 ) ? ( bv_8_126_n456 ) : ( n20959 ) ;
assign n20961 =  ( n20543 ) ? ( bv_8_61_n634 ) : ( n20960 ) ;
assign n20962 =  ( n20541 ) ? ( bv_8_100_n348 ) : ( n20961 ) ;
assign n20963 =  ( n20539 ) ? ( bv_8_93_n498 ) : ( n20962 ) ;
assign n20964 =  ( n20537 ) ? ( bv_8_25_n399 ) : ( n20963 ) ;
assign n20965 =  ( n20535 ) ? ( bv_8_115_n222 ) : ( n20964 ) ;
assign n20966 =  ( n20533 ) ? ( bv_8_96_n542 ) : ( n20965 ) ;
assign n20967 =  ( n20531 ) ? ( bv_8_129_n446 ) : ( n20966 ) ;
assign n20968 =  ( n20529 ) ? ( bv_8_79_n538 ) : ( n20967 ) ;
assign n20969 =  ( n20527 ) ? ( bv_8_220_n142 ) : ( n20968 ) ;
assign n20970 =  ( n20525 ) ? ( bv_8_34_n117 ) : ( n20969 ) ;
assign n20971 =  ( n20523 ) ? ( bv_8_42_n672 ) : ( n20970 ) ;
assign n20972 =  ( n20521 ) ? ( bv_8_144_n173 ) : ( n20971 ) ;
assign n20973 =  ( n20519 ) ? ( bv_8_136_n425 ) : ( n20972 ) ;
assign n20974 =  ( n20517 ) ? ( bv_8_70_n609 ) : ( n20973 ) ;
assign n20975 =  ( n20515 ) ? ( bv_8_238_n71 ) : ( n20974 ) ;
assign n20976 =  ( n20513 ) ? ( bv_8_184_n270 ) : ( n20975 ) ;
assign n20977 =  ( n20511 ) ? ( bv_8_20_n341 ) : ( n20976 ) ;
assign n20978 =  ( n20509 ) ? ( bv_8_222_n134 ) : ( n20977 ) ;
assign n20979 =  ( n20507 ) ? ( bv_8_94_n548 ) : ( n20978 ) ;
assign n20980 =  ( n20505 ) ? ( bv_8_11_n379 ) : ( n20979 ) ;
assign n20981 =  ( n20503 ) ? ( bv_8_219_n146 ) : ( n20980 ) ;
assign n20982 =  ( n20501 ) ? ( bv_8_224_n126 ) : ( n20981 ) ;
assign n20983 =  ( n20499 ) ? ( bv_8_50_n408 ) : ( n20982 ) ;
assign n20984 =  ( n20497 ) ? ( bv_8_58_n136 ) : ( n20983 ) ;
assign n20985 =  ( n20495 ) ? ( bv_8_10_n655 ) : ( n20984 ) ;
assign n20986 =  ( n20493 ) ? ( bv_8_73_n275 ) : ( n20985 ) ;
assign n20987 =  ( n20491 ) ? ( bv_8_6_n169 ) : ( n20986 ) ;
assign n20988 =  ( n20489 ) ? ( bv_8_36_n645 ) : ( n20987 ) ;
assign n20989 =  ( n20487 ) ? ( bv_8_92_n234 ) : ( n20988 ) ;
assign n20990 =  ( n20485 ) ? ( bv_8_194_n159 ) : ( n20989 ) ;
assign n20991 =  ( n20483 ) ? ( bv_8_211_n175 ) : ( n20990 ) ;
assign n20992 =  ( n20481 ) ? ( bv_8_172_n268 ) : ( n20991 ) ;
assign n20993 =  ( n20479 ) ? ( bv_8_98_n536 ) : ( n20992 ) ;
assign n20994 =  ( n20477 ) ? ( bv_8_145_n397 ) : ( n20993 ) ;
assign n20995 =  ( n20475 ) ? ( bv_8_149_n384 ) : ( n20994 ) ;
assign n20996 =  ( n20473 ) ? ( bv_8_228_n111 ) : ( n20995 ) ;
assign n20997 =  ( n20471 ) ? ( bv_8_121_n470 ) : ( n20996 ) ;
assign n20998 =  ( n20469 ) ? ( bv_8_231_n99 ) : ( n20997 ) ;
assign n20999 =  ( n20467 ) ? ( bv_8_200_n213 ) : ( n20998 ) ;
assign n21000 =  ( n20465 ) ? ( bv_8_55_n650 ) : ( n20999 ) ;
assign n21001 =  ( n20463 ) ? ( bv_8_109_n9 ) : ( n21000 ) ;
assign n21002 =  ( n20461 ) ? ( bv_8_141_n410 ) : ( n21001 ) ;
assign n21003 =  ( n20459 ) ? ( bv_8_213_n167 ) : ( n21002 ) ;
assign n21004 =  ( n20457 ) ? ( bv_8_78_n590 ) : ( n21003 ) ;
assign n21005 =  ( n20455 ) ? ( bv_8_169_n109 ) : ( n21004 ) ;
assign n21006 =  ( n20453 ) ? ( bv_8_108_n510 ) : ( n21005 ) ;
assign n21007 =  ( n20451 ) ? ( bv_8_86_n567 ) : ( n21006 ) ;
assign n21008 =  ( n20449 ) ? ( bv_8_244_n47 ) : ( n21007 ) ;
assign n21009 =  ( n20447 ) ? ( bv_8_234_n87 ) : ( n21008 ) ;
assign n21010 =  ( n20445 ) ? ( bv_8_101_n49 ) : ( n21009 ) ;
assign n21011 =  ( n20443 ) ? ( bv_8_122_n416 ) : ( n21010 ) ;
assign n21012 =  ( n20441 ) ? ( bv_8_174_n152 ) : ( n21011 ) ;
assign n21013 =  ( n20439 ) ? ( bv_8_8_n669 ) : ( n21012 ) ;
assign n21014 =  ( n20437 ) ? ( bv_8_186_n263 ) : ( n21013 ) ;
assign n21015 =  ( n20435 ) ? ( bv_8_120_n474 ) : ( n21014 ) ;
assign n21016 =  ( n20433 ) ? ( bv_8_37_n506 ) : ( n21015 ) ;
assign n21017 =  ( n20431 ) ? ( bv_8_46_n429 ) : ( n21016 ) ;
assign n21018 =  ( n20429 ) ? ( bv_8_28_n162 ) : ( n21017 ) ;
assign n21019 =  ( n20427 ) ? ( bv_8_166_n328 ) : ( n21018 ) ;
assign n21020 =  ( n20425 ) ? ( bv_8_180_n285 ) : ( n21019 ) ;
assign n21021 =  ( n20423 ) ? ( bv_8_198_n220 ) : ( n21020 ) ;
assign n21022 =  ( n20421 ) ? ( bv_8_232_n95 ) : ( n21021 ) ;
assign n21023 =  ( n20419 ) ? ( bv_8_221_n138 ) : ( n21022 ) ;
assign n21024 =  ( n20417 ) ? ( bv_8_116_n345 ) : ( n21023 ) ;
assign n21025 =  ( n20415 ) ? ( bv_8_31_n705 ) : ( n21024 ) ;
assign n21026 =  ( n20413 ) ? ( bv_8_75_n503 ) : ( n21025 ) ;
assign n21027 =  ( n20411 ) ? ( bv_8_189_n254 ) : ( n21026 ) ;
assign n21028 =  ( n20409 ) ? ( bv_8_139_n297 ) : ( n21027 ) ;
assign n21029 =  ( n20407 ) ? ( bv_8_138_n418 ) : ( n21028 ) ;
assign n21030 =  ( n20405 ) ? ( bv_8_112_n482 ) : ( n21029 ) ;
assign n21031 =  ( n20403 ) ? ( bv_8_62_n205 ) : ( n21030 ) ;
assign n21032 =  ( n20401 ) ? ( bv_8_181_n281 ) : ( n21031 ) ;
assign n21033 =  ( n20399 ) ? ( bv_8_102_n527 ) : ( n21032 ) ;
assign n21034 =  ( n20397 ) ? ( bv_8_72_n330 ) : ( n21033 ) ;
assign n21035 =  ( n20395 ) ? ( bv_8_3_n65 ) : ( n21034 ) ;
assign n21036 =  ( n20393 ) ? ( bv_8_246_n39 ) : ( n21035 ) ;
assign n21037 =  ( n20391 ) ? ( bv_8_14_n648 ) : ( n21036 ) ;
assign n21038 =  ( n20389 ) ? ( bv_8_97_n198 ) : ( n21037 ) ;
assign n21039 =  ( n20387 ) ? ( bv_8_53_n436 ) : ( n21038 ) ;
assign n21040 =  ( n20385 ) ? ( bv_8_87_n226 ) : ( n21039 ) ;
assign n21041 =  ( n20383 ) ? ( bv_8_185_n266 ) : ( n21040 ) ;
assign n21042 =  ( n20381 ) ? ( bv_8_134_n431 ) : ( n21041 ) ;
assign n21043 =  ( n20379 ) ? ( bv_8_193_n239 ) : ( n21042 ) ;
assign n21044 =  ( n20377 ) ? ( bv_8_29_n625 ) : ( n21043 ) ;
assign n21045 =  ( n20375 ) ? ( bv_8_158_n355 ) : ( n21044 ) ;
assign n21046 =  ( n20373 ) ? ( bv_8_225_n123 ) : ( n21045 ) ;
assign n21047 =  ( n20371 ) ? ( bv_8_248_n31 ) : ( n21046 ) ;
assign n21048 =  ( n20369 ) ? ( bv_8_152_n374 ) : ( n21047 ) ;
assign n21049 =  ( n20367 ) ? ( bv_8_17_n525 ) : ( n21048 ) ;
assign n21050 =  ( n20365 ) ? ( bv_8_105_n148 ) : ( n21049 ) ;
assign n21051 =  ( n20363 ) ? ( bv_8_217_n128 ) : ( n21050 ) ;
assign n21052 =  ( n20361 ) ? ( bv_8_142_n406 ) : ( n21051 ) ;
assign n21053 =  ( n20359 ) ? ( bv_8_148_n388 ) : ( n21052 ) ;
assign n21054 =  ( n20357 ) ? ( bv_8_155_n364 ) : ( n21053 ) ;
assign n21055 =  ( n20355 ) ? ( bv_8_30_n21 ) : ( n21054 ) ;
assign n21056 =  ( n20353 ) ? ( bv_8_135_n81 ) : ( n21055 ) ;
assign n21057 =  ( n20351 ) ? ( bv_8_233_n91 ) : ( n21056 ) ;
assign n21058 =  ( n20349 ) ? ( bv_8_206_n192 ) : ( n21057 ) ;
assign n21059 =  ( n20347 ) ? ( bv_8_85_n423 ) : ( n21058 ) ;
assign n21060 =  ( n20345 ) ? ( bv_8_40_n366 ) : ( n21059 ) ;
assign n21061 =  ( n20343 ) ? ( bv_8_223_n130 ) : ( n21060 ) ;
assign n21062 =  ( n20341 ) ? ( bv_8_140_n376 ) : ( n21061 ) ;
assign n21063 =  ( n20339 ) ? ( bv_8_161_n211 ) : ( n21062 ) ;
assign n21064 =  ( n20337 ) ? ( bv_8_137_n421 ) : ( n21063 ) ;
assign n21065 =  ( n20335 ) ? ( bv_8_13_n194 ) : ( n21064 ) ;
assign n21066 =  ( n20333 ) ? ( bv_8_191_n246 ) : ( n21065 ) ;
assign n21067 =  ( n20331 ) ? ( bv_8_230_n103 ) : ( n21066 ) ;
assign n21068 =  ( n20329 ) ? ( bv_8_66_n466 ) : ( n21067 ) ;
assign n21069 =  ( n20327 ) ? ( bv_8_104_n520 ) : ( n21068 ) ;
assign n21070 =  ( n20325 ) ? ( bv_8_65_n623 ) : ( n21069 ) ;
assign n21071 =  ( n20323 ) ? ( bv_8_153_n140 ) : ( n21070 ) ;
assign n21072 =  ( n20321 ) ? ( bv_8_45_n97 ) : ( n21071 ) ;
assign n21073 =  ( n20319 ) ? ( bv_8_15_n190 ) : ( n21072 ) ;
assign n21074 =  ( n20317 ) ? ( bv_8_176_n299 ) : ( n21073 ) ;
assign n21075 =  ( n20315 ) ? ( bv_8_84_n386 ) : ( n21074 ) ;
assign n21076 =  ( n20313 ) ? ( bv_8_187_n260 ) : ( n21075 ) ;
assign n21077 =  ( n20311 ) ? ( bv_8_22_n357 ) : ( n21076 ) ;
assign n21078 =  ( n20309 ) ^ ( n21077 )  ;
assign n21079 = state_in[39:32] ;
assign n21080 =  ( n21079 ) == ( bv_8_255_n3 )  ;
assign n21081 = state_in[39:32] ;
assign n21082 =  ( n21081 ) == ( bv_8_254_n7 )  ;
assign n21083 = state_in[39:32] ;
assign n21084 =  ( n21083 ) == ( bv_8_253_n11 )  ;
assign n21085 = state_in[39:32] ;
assign n21086 =  ( n21085 ) == ( bv_8_252_n15 )  ;
assign n21087 = state_in[39:32] ;
assign n21088 =  ( n21087 ) == ( bv_8_251_n19 )  ;
assign n21089 = state_in[39:32] ;
assign n21090 =  ( n21089 ) == ( bv_8_250_n23 )  ;
assign n21091 = state_in[39:32] ;
assign n21092 =  ( n21091 ) == ( bv_8_249_n27 )  ;
assign n21093 = state_in[39:32] ;
assign n21094 =  ( n21093 ) == ( bv_8_248_n31 )  ;
assign n21095 = state_in[39:32] ;
assign n21096 =  ( n21095 ) == ( bv_8_247_n35 )  ;
assign n21097 = state_in[39:32] ;
assign n21098 =  ( n21097 ) == ( bv_8_246_n39 )  ;
assign n21099 = state_in[39:32] ;
assign n21100 =  ( n21099 ) == ( bv_8_245_n43 )  ;
assign n21101 = state_in[39:32] ;
assign n21102 =  ( n21101 ) == ( bv_8_244_n47 )  ;
assign n21103 = state_in[39:32] ;
assign n21104 =  ( n21103 ) == ( bv_8_243_n51 )  ;
assign n21105 = state_in[39:32] ;
assign n21106 =  ( n21105 ) == ( bv_8_242_n55 )  ;
assign n21107 = state_in[39:32] ;
assign n21108 =  ( n21107 ) == ( bv_8_241_n59 )  ;
assign n21109 = state_in[39:32] ;
assign n21110 =  ( n21109 ) == ( bv_8_240_n63 )  ;
assign n21111 = state_in[39:32] ;
assign n21112 =  ( n21111 ) == ( bv_8_239_n67 )  ;
assign n21113 = state_in[39:32] ;
assign n21114 =  ( n21113 ) == ( bv_8_238_n71 )  ;
assign n21115 = state_in[39:32] ;
assign n21116 =  ( n21115 ) == ( bv_8_237_n75 )  ;
assign n21117 = state_in[39:32] ;
assign n21118 =  ( n21117 ) == ( bv_8_236_n79 )  ;
assign n21119 = state_in[39:32] ;
assign n21120 =  ( n21119 ) == ( bv_8_235_n83 )  ;
assign n21121 = state_in[39:32] ;
assign n21122 =  ( n21121 ) == ( bv_8_234_n87 )  ;
assign n21123 = state_in[39:32] ;
assign n21124 =  ( n21123 ) == ( bv_8_233_n91 )  ;
assign n21125 = state_in[39:32] ;
assign n21126 =  ( n21125 ) == ( bv_8_232_n95 )  ;
assign n21127 = state_in[39:32] ;
assign n21128 =  ( n21127 ) == ( bv_8_231_n99 )  ;
assign n21129 = state_in[39:32] ;
assign n21130 =  ( n21129 ) == ( bv_8_230_n103 )  ;
assign n21131 = state_in[39:32] ;
assign n21132 =  ( n21131 ) == ( bv_8_229_n107 )  ;
assign n21133 = state_in[39:32] ;
assign n21134 =  ( n21133 ) == ( bv_8_228_n111 )  ;
assign n21135 = state_in[39:32] ;
assign n21136 =  ( n21135 ) == ( bv_8_227_n115 )  ;
assign n21137 = state_in[39:32] ;
assign n21138 =  ( n21137 ) == ( bv_8_226_n119 )  ;
assign n21139 = state_in[39:32] ;
assign n21140 =  ( n21139 ) == ( bv_8_225_n123 )  ;
assign n21141 = state_in[39:32] ;
assign n21142 =  ( n21141 ) == ( bv_8_224_n126 )  ;
assign n21143 = state_in[39:32] ;
assign n21144 =  ( n21143 ) == ( bv_8_223_n130 )  ;
assign n21145 = state_in[39:32] ;
assign n21146 =  ( n21145 ) == ( bv_8_222_n134 )  ;
assign n21147 = state_in[39:32] ;
assign n21148 =  ( n21147 ) == ( bv_8_221_n138 )  ;
assign n21149 = state_in[39:32] ;
assign n21150 =  ( n21149 ) == ( bv_8_220_n142 )  ;
assign n21151 = state_in[39:32] ;
assign n21152 =  ( n21151 ) == ( bv_8_219_n146 )  ;
assign n21153 = state_in[39:32] ;
assign n21154 =  ( n21153 ) == ( bv_8_218_n150 )  ;
assign n21155 = state_in[39:32] ;
assign n21156 =  ( n21155 ) == ( bv_8_217_n128 )  ;
assign n21157 = state_in[39:32] ;
assign n21158 =  ( n21157 ) == ( bv_8_216_n157 )  ;
assign n21159 = state_in[39:32] ;
assign n21160 =  ( n21159 ) == ( bv_8_215_n45 )  ;
assign n21161 = state_in[39:32] ;
assign n21162 =  ( n21161 ) == ( bv_8_214_n164 )  ;
assign n21163 = state_in[39:32] ;
assign n21164 =  ( n21163 ) == ( bv_8_213_n167 )  ;
assign n21165 = state_in[39:32] ;
assign n21166 =  ( n21165 ) == ( bv_8_212_n171 )  ;
assign n21167 = state_in[39:32] ;
assign n21168 =  ( n21167 ) == ( bv_8_211_n175 )  ;
assign n21169 = state_in[39:32] ;
assign n21170 =  ( n21169 ) == ( bv_8_210_n113 )  ;
assign n21171 = state_in[39:32] ;
assign n21172 =  ( n21171 ) == ( bv_8_209_n182 )  ;
assign n21173 = state_in[39:32] ;
assign n21174 =  ( n21173 ) == ( bv_8_208_n37 )  ;
assign n21175 = state_in[39:32] ;
assign n21176 =  ( n21175 ) == ( bv_8_207_n188 )  ;
assign n21177 = state_in[39:32] ;
assign n21178 =  ( n21177 ) == ( bv_8_206_n192 )  ;
assign n21179 = state_in[39:32] ;
assign n21180 =  ( n21179 ) == ( bv_8_205_n196 )  ;
assign n21181 = state_in[39:32] ;
assign n21182 =  ( n21181 ) == ( bv_8_204_n177 )  ;
assign n21183 = state_in[39:32] ;
assign n21184 =  ( n21183 ) == ( bv_8_203_n203 )  ;
assign n21185 = state_in[39:32] ;
assign n21186 =  ( n21185 ) == ( bv_8_202_n207 )  ;
assign n21187 = state_in[39:32] ;
assign n21188 =  ( n21187 ) == ( bv_8_201_n85 )  ;
assign n21189 = state_in[39:32] ;
assign n21190 =  ( n21189 ) == ( bv_8_200_n213 )  ;
assign n21191 = state_in[39:32] ;
assign n21192 =  ( n21191 ) == ( bv_8_199_n216 )  ;
assign n21193 = state_in[39:32] ;
assign n21194 =  ( n21193 ) == ( bv_8_198_n220 )  ;
assign n21195 = state_in[39:32] ;
assign n21196 =  ( n21195 ) == ( bv_8_197_n224 )  ;
assign n21197 = state_in[39:32] ;
assign n21198 =  ( n21197 ) == ( bv_8_196_n228 )  ;
assign n21199 = state_in[39:32] ;
assign n21200 =  ( n21199 ) == ( bv_8_195_n232 )  ;
assign n21201 = state_in[39:32] ;
assign n21202 =  ( n21201 ) == ( bv_8_194_n159 )  ;
assign n21203 = state_in[39:32] ;
assign n21204 =  ( n21203 ) == ( bv_8_193_n239 )  ;
assign n21205 = state_in[39:32] ;
assign n21206 =  ( n21205 ) == ( bv_8_192_n242 )  ;
assign n21207 = state_in[39:32] ;
assign n21208 =  ( n21207 ) == ( bv_8_191_n246 )  ;
assign n21209 = state_in[39:32] ;
assign n21210 =  ( n21209 ) == ( bv_8_190_n250 )  ;
assign n21211 = state_in[39:32] ;
assign n21212 =  ( n21211 ) == ( bv_8_189_n254 )  ;
assign n21213 = state_in[39:32] ;
assign n21214 =  ( n21213 ) == ( bv_8_188_n257 )  ;
assign n21215 = state_in[39:32] ;
assign n21216 =  ( n21215 ) == ( bv_8_187_n260 )  ;
assign n21217 = state_in[39:32] ;
assign n21218 =  ( n21217 ) == ( bv_8_186_n263 )  ;
assign n21219 = state_in[39:32] ;
assign n21220 =  ( n21219 ) == ( bv_8_185_n266 )  ;
assign n21221 = state_in[39:32] ;
assign n21222 =  ( n21221 ) == ( bv_8_184_n270 )  ;
assign n21223 = state_in[39:32] ;
assign n21224 =  ( n21223 ) == ( bv_8_183_n273 )  ;
assign n21225 = state_in[39:32] ;
assign n21226 =  ( n21225 ) == ( bv_8_182_n277 )  ;
assign n21227 = state_in[39:32] ;
assign n21228 =  ( n21227 ) == ( bv_8_181_n281 )  ;
assign n21229 = state_in[39:32] ;
assign n21230 =  ( n21229 ) == ( bv_8_180_n285 )  ;
assign n21231 = state_in[39:32] ;
assign n21232 =  ( n21231 ) == ( bv_8_179_n289 )  ;
assign n21233 = state_in[39:32] ;
assign n21234 =  ( n21233 ) == ( bv_8_178_n292 )  ;
assign n21235 = state_in[39:32] ;
assign n21236 =  ( n21235 ) == ( bv_8_177_n283 )  ;
assign n21237 = state_in[39:32] ;
assign n21238 =  ( n21237 ) == ( bv_8_176_n299 )  ;
assign n21239 = state_in[39:32] ;
assign n21240 =  ( n21239 ) == ( bv_8_175_n302 )  ;
assign n21241 = state_in[39:32] ;
assign n21242 =  ( n21241 ) == ( bv_8_174_n152 )  ;
assign n21243 = state_in[39:32] ;
assign n21244 =  ( n21243 ) == ( bv_8_173_n307 )  ;
assign n21245 = state_in[39:32] ;
assign n21246 =  ( n21245 ) == ( bv_8_172_n268 )  ;
assign n21247 = state_in[39:32] ;
assign n21248 =  ( n21247 ) == ( bv_8_171_n314 )  ;
assign n21249 = state_in[39:32] ;
assign n21250 =  ( n21249 ) == ( bv_8_170_n77 )  ;
assign n21251 = state_in[39:32] ;
assign n21252 =  ( n21251 ) == ( bv_8_169_n109 )  ;
assign n21253 = state_in[39:32] ;
assign n21254 =  ( n21253 ) == ( bv_8_168_n13 )  ;
assign n21255 = state_in[39:32] ;
assign n21256 =  ( n21255 ) == ( bv_8_167_n325 )  ;
assign n21257 = state_in[39:32] ;
assign n21258 =  ( n21257 ) == ( bv_8_166_n328 )  ;
assign n21259 = state_in[39:32] ;
assign n21260 =  ( n21259 ) == ( bv_8_165_n69 )  ;
assign n21261 = state_in[39:32] ;
assign n21262 =  ( n21261 ) == ( bv_8_164_n335 )  ;
assign n21263 = state_in[39:32] ;
assign n21264 =  ( n21263 ) == ( bv_8_163_n339 )  ;
assign n21265 = state_in[39:32] ;
assign n21266 =  ( n21265 ) == ( bv_8_162_n343 )  ;
assign n21267 = state_in[39:32] ;
assign n21268 =  ( n21267 ) == ( bv_8_161_n211 )  ;
assign n21269 = state_in[39:32] ;
assign n21270 =  ( n21269 ) == ( bv_8_160_n350 )  ;
assign n21271 = state_in[39:32] ;
assign n21272 =  ( n21271 ) == ( bv_8_159_n323 )  ;
assign n21273 = state_in[39:32] ;
assign n21274 =  ( n21273 ) == ( bv_8_158_n355 )  ;
assign n21275 = state_in[39:32] ;
assign n21276 =  ( n21275 ) == ( bv_8_157_n359 )  ;
assign n21277 = state_in[39:32] ;
assign n21278 =  ( n21277 ) == ( bv_8_156_n279 )  ;
assign n21279 = state_in[39:32] ;
assign n21280 =  ( n21279 ) == ( bv_8_155_n364 )  ;
assign n21281 = state_in[39:32] ;
assign n21282 =  ( n21281 ) == ( bv_8_154_n368 )  ;
assign n21283 = state_in[39:32] ;
assign n21284 =  ( n21283 ) == ( bv_8_153_n140 )  ;
assign n21285 = state_in[39:32] ;
assign n21286 =  ( n21285 ) == ( bv_8_152_n374 )  ;
assign n21287 = state_in[39:32] ;
assign n21288 =  ( n21287 ) == ( bv_8_151_n218 )  ;
assign n21289 = state_in[39:32] ;
assign n21290 =  ( n21289 ) == ( bv_8_150_n201 )  ;
assign n21291 = state_in[39:32] ;
assign n21292 =  ( n21291 ) == ( bv_8_149_n384 )  ;
assign n21293 = state_in[39:32] ;
assign n21294 =  ( n21293 ) == ( bv_8_148_n388 )  ;
assign n21295 = state_in[39:32] ;
assign n21296 =  ( n21295 ) == ( bv_8_147_n392 )  ;
assign n21297 = state_in[39:32] ;
assign n21298 =  ( n21297 ) == ( bv_8_146_n337 )  ;
assign n21299 = state_in[39:32] ;
assign n21300 =  ( n21299 ) == ( bv_8_145_n397 )  ;
assign n21301 = state_in[39:32] ;
assign n21302 =  ( n21301 ) == ( bv_8_144_n173 )  ;
assign n21303 = state_in[39:32] ;
assign n21304 =  ( n21303 ) == ( bv_8_143_n403 )  ;
assign n21305 = state_in[39:32] ;
assign n21306 =  ( n21305 ) == ( bv_8_142_n406 )  ;
assign n21307 = state_in[39:32] ;
assign n21308 =  ( n21307 ) == ( bv_8_141_n410 )  ;
assign n21309 = state_in[39:32] ;
assign n21310 =  ( n21309 ) == ( bv_8_140_n376 )  ;
assign n21311 = state_in[39:32] ;
assign n21312 =  ( n21311 ) == ( bv_8_139_n297 )  ;
assign n21313 = state_in[39:32] ;
assign n21314 =  ( n21313 ) == ( bv_8_138_n418 )  ;
assign n21315 = state_in[39:32] ;
assign n21316 =  ( n21315 ) == ( bv_8_137_n421 )  ;
assign n21317 = state_in[39:32] ;
assign n21318 =  ( n21317 ) == ( bv_8_136_n425 )  ;
assign n21319 = state_in[39:32] ;
assign n21320 =  ( n21319 ) == ( bv_8_135_n81 )  ;
assign n21321 = state_in[39:32] ;
assign n21322 =  ( n21321 ) == ( bv_8_134_n431 )  ;
assign n21323 = state_in[39:32] ;
assign n21324 =  ( n21323 ) == ( bv_8_133_n434 )  ;
assign n21325 = state_in[39:32] ;
assign n21326 =  ( n21325 ) == ( bv_8_132_n41 )  ;
assign n21327 = state_in[39:32] ;
assign n21328 =  ( n21327 ) == ( bv_8_131_n440 )  ;
assign n21329 = state_in[39:32] ;
assign n21330 =  ( n21329 ) == ( bv_8_130_n33 )  ;
assign n21331 = state_in[39:32] ;
assign n21332 =  ( n21331 ) == ( bv_8_129_n446 )  ;
assign n21333 = state_in[39:32] ;
assign n21334 =  ( n21333 ) == ( bv_8_128_n450 )  ;
assign n21335 = state_in[39:32] ;
assign n21336 =  ( n21335 ) == ( bv_8_127_n453 )  ;
assign n21337 = state_in[39:32] ;
assign n21338 =  ( n21337 ) == ( bv_8_126_n456 )  ;
assign n21339 = state_in[39:32] ;
assign n21340 =  ( n21339 ) == ( bv_8_125_n459 )  ;
assign n21341 = state_in[39:32] ;
assign n21342 =  ( n21341 ) == ( bv_8_124_n184 )  ;
assign n21343 = state_in[39:32] ;
assign n21344 =  ( n21343 ) == ( bv_8_123_n17 )  ;
assign n21345 = state_in[39:32] ;
assign n21346 =  ( n21345 ) == ( bv_8_122_n416 )  ;
assign n21347 = state_in[39:32] ;
assign n21348 =  ( n21347 ) == ( bv_8_121_n470 )  ;
assign n21349 = state_in[39:32] ;
assign n21350 =  ( n21349 ) == ( bv_8_120_n474 )  ;
assign n21351 = state_in[39:32] ;
assign n21352 =  ( n21351 ) == ( bv_8_119_n472 )  ;
assign n21353 = state_in[39:32] ;
assign n21354 =  ( n21353 ) == ( bv_8_118_n480 )  ;
assign n21355 = state_in[39:32] ;
assign n21356 =  ( n21355 ) == ( bv_8_117_n484 )  ;
assign n21357 = state_in[39:32] ;
assign n21358 =  ( n21357 ) == ( bv_8_116_n345 )  ;
assign n21359 = state_in[39:32] ;
assign n21360 =  ( n21359 ) == ( bv_8_115_n222 )  ;
assign n21361 = state_in[39:32] ;
assign n21362 =  ( n21361 ) == ( bv_8_114_n494 )  ;
assign n21363 = state_in[39:32] ;
assign n21364 =  ( n21363 ) == ( bv_8_113_n180 )  ;
assign n21365 = state_in[39:32] ;
assign n21366 =  ( n21365 ) == ( bv_8_112_n482 )  ;
assign n21367 = state_in[39:32] ;
assign n21368 =  ( n21367 ) == ( bv_8_111_n244 )  ;
assign n21369 = state_in[39:32] ;
assign n21370 =  ( n21369 ) == ( bv_8_110_n294 )  ;
assign n21371 = state_in[39:32] ;
assign n21372 =  ( n21371 ) == ( bv_8_109_n9 )  ;
assign n21373 = state_in[39:32] ;
assign n21374 =  ( n21373 ) == ( bv_8_108_n510 )  ;
assign n21375 = state_in[39:32] ;
assign n21376 =  ( n21375 ) == ( bv_8_107_n370 )  ;
assign n21377 = state_in[39:32] ;
assign n21378 =  ( n21377 ) == ( bv_8_106_n155 )  ;
assign n21379 = state_in[39:32] ;
assign n21380 =  ( n21379 ) == ( bv_8_105_n148 )  ;
assign n21381 = state_in[39:32] ;
assign n21382 =  ( n21381 ) == ( bv_8_104_n520 )  ;
assign n21383 = state_in[39:32] ;
assign n21384 =  ( n21383 ) == ( bv_8_103_n523 )  ;
assign n21385 = state_in[39:32] ;
assign n21386 =  ( n21385 ) == ( bv_8_102_n527 )  ;
assign n21387 = state_in[39:32] ;
assign n21388 =  ( n21387 ) == ( bv_8_101_n49 )  ;
assign n21389 = state_in[39:32] ;
assign n21390 =  ( n21389 ) == ( bv_8_100_n348 )  ;
assign n21391 = state_in[39:32] ;
assign n21392 =  ( n21391 ) == ( bv_8_99_n476 )  ;
assign n21393 = state_in[39:32] ;
assign n21394 =  ( n21393 ) == ( bv_8_98_n536 )  ;
assign n21395 = state_in[39:32] ;
assign n21396 =  ( n21395 ) == ( bv_8_97_n198 )  ;
assign n21397 = state_in[39:32] ;
assign n21398 =  ( n21397 ) == ( bv_8_96_n542 )  ;
assign n21399 = state_in[39:32] ;
assign n21400 =  ( n21399 ) == ( bv_8_95_n545 )  ;
assign n21401 = state_in[39:32] ;
assign n21402 =  ( n21401 ) == ( bv_8_94_n548 )  ;
assign n21403 = state_in[39:32] ;
assign n21404 =  ( n21403 ) == ( bv_8_93_n498 )  ;
assign n21405 = state_in[39:32] ;
assign n21406 =  ( n21405 ) == ( bv_8_92_n234 )  ;
assign n21407 = state_in[39:32] ;
assign n21408 =  ( n21407 ) == ( bv_8_91_n555 )  ;
assign n21409 = state_in[39:32] ;
assign n21410 =  ( n21409 ) == ( bv_8_90_n25 )  ;
assign n21411 = state_in[39:32] ;
assign n21412 =  ( n21411 ) == ( bv_8_89_n61 )  ;
assign n21413 = state_in[39:32] ;
assign n21414 =  ( n21413 ) == ( bv_8_88_n562 )  ;
assign n21415 = state_in[39:32] ;
assign n21416 =  ( n21415 ) == ( bv_8_87_n226 )  ;
assign n21417 = state_in[39:32] ;
assign n21418 =  ( n21417 ) == ( bv_8_86_n567 )  ;
assign n21419 = state_in[39:32] ;
assign n21420 =  ( n21419 ) == ( bv_8_85_n423 )  ;
assign n21421 = state_in[39:32] ;
assign n21422 =  ( n21421 ) == ( bv_8_84_n386 )  ;
assign n21423 = state_in[39:32] ;
assign n21424 =  ( n21423 ) == ( bv_8_83_n575 )  ;
assign n21425 = state_in[39:32] ;
assign n21426 =  ( n21425 ) == ( bv_8_82_n578 )  ;
assign n21427 = state_in[39:32] ;
assign n21428 =  ( n21427 ) == ( bv_8_81_n582 )  ;
assign n21429 = state_in[39:32] ;
assign n21430 =  ( n21429 ) == ( bv_8_80_n73 )  ;
assign n21431 = state_in[39:32] ;
assign n21432 =  ( n21431 ) == ( bv_8_79_n538 )  ;
assign n21433 = state_in[39:32] ;
assign n21434 =  ( n21433 ) == ( bv_8_78_n590 )  ;
assign n21435 = state_in[39:32] ;
assign n21436 =  ( n21435 ) == ( bv_8_77_n593 )  ;
assign n21437 = state_in[39:32] ;
assign n21438 =  ( n21437 ) == ( bv_8_76_n596 )  ;
assign n21439 = state_in[39:32] ;
assign n21440 =  ( n21439 ) == ( bv_8_75_n503 )  ;
assign n21441 = state_in[39:32] ;
assign n21442 =  ( n21441 ) == ( bv_8_74_n237 )  ;
assign n21443 = state_in[39:32] ;
assign n21444 =  ( n21443 ) == ( bv_8_73_n275 )  ;
assign n21445 = state_in[39:32] ;
assign n21446 =  ( n21445 ) == ( bv_8_72_n330 )  ;
assign n21447 = state_in[39:32] ;
assign n21448 =  ( n21447 ) == ( bv_8_71_n252 )  ;
assign n21449 = state_in[39:32] ;
assign n21450 =  ( n21449 ) == ( bv_8_70_n609 )  ;
assign n21451 = state_in[39:32] ;
assign n21452 =  ( n21451 ) == ( bv_8_69_n612 )  ;
assign n21453 = state_in[39:32] ;
assign n21454 =  ( n21453 ) == ( bv_8_68_n390 )  ;
assign n21455 = state_in[39:32] ;
assign n21456 =  ( n21455 ) == ( bv_8_67_n318 )  ;
assign n21457 = state_in[39:32] ;
assign n21458 =  ( n21457 ) == ( bv_8_66_n466 )  ;
assign n21459 = state_in[39:32] ;
assign n21460 =  ( n21459 ) == ( bv_8_65_n623 )  ;
assign n21461 = state_in[39:32] ;
assign n21462 =  ( n21461 ) == ( bv_8_64_n573 )  ;
assign n21463 = state_in[39:32] ;
assign n21464 =  ( n21463 ) == ( bv_8_63_n489 )  ;
assign n21465 = state_in[39:32] ;
assign n21466 =  ( n21465 ) == ( bv_8_62_n205 )  ;
assign n21467 = state_in[39:32] ;
assign n21468 =  ( n21467 ) == ( bv_8_61_n634 )  ;
assign n21469 = state_in[39:32] ;
assign n21470 =  ( n21469 ) == ( bv_8_60_n93 )  ;
assign n21471 = state_in[39:32] ;
assign n21472 =  ( n21471 ) == ( bv_8_59_n382 )  ;
assign n21473 = state_in[39:32] ;
assign n21474 =  ( n21473 ) == ( bv_8_58_n136 )  ;
assign n21475 = state_in[39:32] ;
assign n21476 =  ( n21475 ) == ( bv_8_57_n312 )  ;
assign n21477 = state_in[39:32] ;
assign n21478 =  ( n21477 ) == ( bv_8_56_n230 )  ;
assign n21479 = state_in[39:32] ;
assign n21480 =  ( n21479 ) == ( bv_8_55_n650 )  ;
assign n21481 = state_in[39:32] ;
assign n21482 =  ( n21481 ) == ( bv_8_54_n616 )  ;
assign n21483 = state_in[39:32] ;
assign n21484 =  ( n21483 ) == ( bv_8_53_n436 )  ;
assign n21485 = state_in[39:32] ;
assign n21486 =  ( n21485 ) == ( bv_8_52_n619 )  ;
assign n21487 = state_in[39:32] ;
assign n21488 =  ( n21487 ) == ( bv_8_51_n101 )  ;
assign n21489 = state_in[39:32] ;
assign n21490 =  ( n21489 ) == ( bv_8_50_n408 )  ;
assign n21491 = state_in[39:32] ;
assign n21492 =  ( n21491 ) == ( bv_8_49_n309 )  ;
assign n21493 = state_in[39:32] ;
assign n21494 =  ( n21493 ) == ( bv_8_48_n660 )  ;
assign n21495 = state_in[39:32] ;
assign n21496 =  ( n21495 ) == ( bv_8_47_n652 )  ;
assign n21497 = state_in[39:32] ;
assign n21498 =  ( n21497 ) == ( bv_8_46_n429 )  ;
assign n21499 = state_in[39:32] ;
assign n21500 =  ( n21499 ) == ( bv_8_45_n97 )  ;
assign n21501 = state_in[39:32] ;
assign n21502 =  ( n21501 ) == ( bv_8_44_n5 )  ;
assign n21503 = state_in[39:32] ;
assign n21504 =  ( n21503 ) == ( bv_8_43_n121 )  ;
assign n21505 = state_in[39:32] ;
assign n21506 =  ( n21505 ) == ( bv_8_42_n672 )  ;
assign n21507 = state_in[39:32] ;
assign n21508 =  ( n21507 ) == ( bv_8_41_n29 )  ;
assign n21509 = state_in[39:32] ;
assign n21510 =  ( n21509 ) == ( bv_8_40_n366 )  ;
assign n21511 = state_in[39:32] ;
assign n21512 =  ( n21511 ) == ( bv_8_39_n132 )  ;
assign n21513 = state_in[39:32] ;
assign n21514 =  ( n21513 ) == ( bv_8_38_n444 )  ;
assign n21515 = state_in[39:32] ;
assign n21516 =  ( n21515 ) == ( bv_8_37_n506 )  ;
assign n21517 = state_in[39:32] ;
assign n21518 =  ( n21517 ) == ( bv_8_36_n645 )  ;
assign n21519 = state_in[39:32] ;
assign n21520 =  ( n21519 ) == ( bv_8_35_n696 )  ;
assign n21521 = state_in[39:32] ;
assign n21522 =  ( n21521 ) == ( bv_8_34_n117 )  ;
assign n21523 = state_in[39:32] ;
assign n21524 =  ( n21523 ) == ( bv_8_33_n486 )  ;
assign n21525 = state_in[39:32] ;
assign n21526 =  ( n21525 ) == ( bv_8_32_n463 )  ;
assign n21527 = state_in[39:32] ;
assign n21528 =  ( n21527 ) == ( bv_8_31_n705 )  ;
assign n21529 = state_in[39:32] ;
assign n21530 =  ( n21529 ) == ( bv_8_30_n21 )  ;
assign n21531 = state_in[39:32] ;
assign n21532 =  ( n21531 ) == ( bv_8_29_n625 )  ;
assign n21533 = state_in[39:32] ;
assign n21534 =  ( n21533 ) == ( bv_8_28_n162 )  ;
assign n21535 = state_in[39:32] ;
assign n21536 =  ( n21535 ) == ( bv_8_27_n642 )  ;
assign n21537 = state_in[39:32] ;
assign n21538 =  ( n21537 ) == ( bv_8_26_n53 )  ;
assign n21539 = state_in[39:32] ;
assign n21540 =  ( n21539 ) == ( bv_8_25_n399 )  ;
assign n21541 = state_in[39:32] ;
assign n21542 =  ( n21541 ) == ( bv_8_24_n448 )  ;
assign n21543 = state_in[39:32] ;
assign n21544 =  ( n21543 ) == ( bv_8_23_n144 )  ;
assign n21545 = state_in[39:32] ;
assign n21546 =  ( n21545 ) == ( bv_8_22_n357 )  ;
assign n21547 = state_in[39:32] ;
assign n21548 =  ( n21547 ) == ( bv_8_21_n89 )  ;
assign n21549 = state_in[39:32] ;
assign n21550 =  ( n21549 ) == ( bv_8_20_n341 )  ;
assign n21551 = state_in[39:32] ;
assign n21552 =  ( n21551 ) == ( bv_8_19_n588 )  ;
assign n21553 = state_in[39:32] ;
assign n21554 =  ( n21553 ) == ( bv_8_18_n628 )  ;
assign n21555 = state_in[39:32] ;
assign n21556 =  ( n21555 ) == ( bv_8_17_n525 )  ;
assign n21557 = state_in[39:32] ;
assign n21558 =  ( n21557 ) == ( bv_8_16_n248 )  ;
assign n21559 = state_in[39:32] ;
assign n21560 =  ( n21559 ) == ( bv_8_15_n190 )  ;
assign n21561 = state_in[39:32] ;
assign n21562 =  ( n21561 ) == ( bv_8_14_n648 )  ;
assign n21563 = state_in[39:32] ;
assign n21564 =  ( n21563 ) == ( bv_8_13_n194 )  ;
assign n21565 = state_in[39:32] ;
assign n21566 =  ( n21565 ) == ( bv_8_12_n333 )  ;
assign n21567 = state_in[39:32] ;
assign n21568 =  ( n21567 ) == ( bv_8_11_n379 )  ;
assign n21569 = state_in[39:32] ;
assign n21570 =  ( n21569 ) == ( bv_8_10_n655 )  ;
assign n21571 = state_in[39:32] ;
assign n21572 =  ( n21571 ) == ( bv_8_9_n57 )  ;
assign n21573 = state_in[39:32] ;
assign n21574 =  ( n21573 ) == ( bv_8_8_n669 )  ;
assign n21575 = state_in[39:32] ;
assign n21576 =  ( n21575 ) == ( bv_8_7_n105 )  ;
assign n21577 = state_in[39:32] ;
assign n21578 =  ( n21577 ) == ( bv_8_6_n169 )  ;
assign n21579 = state_in[39:32] ;
assign n21580 =  ( n21579 ) == ( bv_8_5_n492 )  ;
assign n21581 = state_in[39:32] ;
assign n21582 =  ( n21581 ) == ( bv_8_4_n516 )  ;
assign n21583 = state_in[39:32] ;
assign n21584 =  ( n21583 ) == ( bv_8_3_n65 )  ;
assign n21585 = state_in[39:32] ;
assign n21586 =  ( n21585 ) == ( bv_8_2_n751 )  ;
assign n21587 = state_in[39:32] ;
assign n21588 =  ( n21587 ) == ( bv_8_1_n287 )  ;
assign n21589 = state_in[39:32] ;
assign n21590 =  ( n21589 ) == ( bv_8_0_n580 )  ;
assign n21591 =  ( n21590 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n21592 =  ( n21588 ) ? ( bv_8_124_n184 ) : ( n21591 ) ;
assign n21593 =  ( n21586 ) ? ( bv_8_119_n472 ) : ( n21592 ) ;
assign n21594 =  ( n21584 ) ? ( bv_8_123_n17 ) : ( n21593 ) ;
assign n21595 =  ( n21582 ) ? ( bv_8_242_n55 ) : ( n21594 ) ;
assign n21596 =  ( n21580 ) ? ( bv_8_107_n370 ) : ( n21595 ) ;
assign n21597 =  ( n21578 ) ? ( bv_8_111_n244 ) : ( n21596 ) ;
assign n21598 =  ( n21576 ) ? ( bv_8_197_n224 ) : ( n21597 ) ;
assign n21599 =  ( n21574 ) ? ( bv_8_48_n660 ) : ( n21598 ) ;
assign n21600 =  ( n21572 ) ? ( bv_8_1_n287 ) : ( n21599 ) ;
assign n21601 =  ( n21570 ) ? ( bv_8_103_n523 ) : ( n21600 ) ;
assign n21602 =  ( n21568 ) ? ( bv_8_43_n121 ) : ( n21601 ) ;
assign n21603 =  ( n21566 ) ? ( bv_8_254_n7 ) : ( n21602 ) ;
assign n21604 =  ( n21564 ) ? ( bv_8_215_n45 ) : ( n21603 ) ;
assign n21605 =  ( n21562 ) ? ( bv_8_171_n314 ) : ( n21604 ) ;
assign n21606 =  ( n21560 ) ? ( bv_8_118_n480 ) : ( n21605 ) ;
assign n21607 =  ( n21558 ) ? ( bv_8_202_n207 ) : ( n21606 ) ;
assign n21608 =  ( n21556 ) ? ( bv_8_130_n33 ) : ( n21607 ) ;
assign n21609 =  ( n21554 ) ? ( bv_8_201_n85 ) : ( n21608 ) ;
assign n21610 =  ( n21552 ) ? ( bv_8_125_n459 ) : ( n21609 ) ;
assign n21611 =  ( n21550 ) ? ( bv_8_250_n23 ) : ( n21610 ) ;
assign n21612 =  ( n21548 ) ? ( bv_8_89_n61 ) : ( n21611 ) ;
assign n21613 =  ( n21546 ) ? ( bv_8_71_n252 ) : ( n21612 ) ;
assign n21614 =  ( n21544 ) ? ( bv_8_240_n63 ) : ( n21613 ) ;
assign n21615 =  ( n21542 ) ? ( bv_8_173_n307 ) : ( n21614 ) ;
assign n21616 =  ( n21540 ) ? ( bv_8_212_n171 ) : ( n21615 ) ;
assign n21617 =  ( n21538 ) ? ( bv_8_162_n343 ) : ( n21616 ) ;
assign n21618 =  ( n21536 ) ? ( bv_8_175_n302 ) : ( n21617 ) ;
assign n21619 =  ( n21534 ) ? ( bv_8_156_n279 ) : ( n21618 ) ;
assign n21620 =  ( n21532 ) ? ( bv_8_164_n335 ) : ( n21619 ) ;
assign n21621 =  ( n21530 ) ? ( bv_8_114_n494 ) : ( n21620 ) ;
assign n21622 =  ( n21528 ) ? ( bv_8_192_n242 ) : ( n21621 ) ;
assign n21623 =  ( n21526 ) ? ( bv_8_183_n273 ) : ( n21622 ) ;
assign n21624 =  ( n21524 ) ? ( bv_8_253_n11 ) : ( n21623 ) ;
assign n21625 =  ( n21522 ) ? ( bv_8_147_n392 ) : ( n21624 ) ;
assign n21626 =  ( n21520 ) ? ( bv_8_38_n444 ) : ( n21625 ) ;
assign n21627 =  ( n21518 ) ? ( bv_8_54_n616 ) : ( n21626 ) ;
assign n21628 =  ( n21516 ) ? ( bv_8_63_n489 ) : ( n21627 ) ;
assign n21629 =  ( n21514 ) ? ( bv_8_247_n35 ) : ( n21628 ) ;
assign n21630 =  ( n21512 ) ? ( bv_8_204_n177 ) : ( n21629 ) ;
assign n21631 =  ( n21510 ) ? ( bv_8_52_n619 ) : ( n21630 ) ;
assign n21632 =  ( n21508 ) ? ( bv_8_165_n69 ) : ( n21631 ) ;
assign n21633 =  ( n21506 ) ? ( bv_8_229_n107 ) : ( n21632 ) ;
assign n21634 =  ( n21504 ) ? ( bv_8_241_n59 ) : ( n21633 ) ;
assign n21635 =  ( n21502 ) ? ( bv_8_113_n180 ) : ( n21634 ) ;
assign n21636 =  ( n21500 ) ? ( bv_8_216_n157 ) : ( n21635 ) ;
assign n21637 =  ( n21498 ) ? ( bv_8_49_n309 ) : ( n21636 ) ;
assign n21638 =  ( n21496 ) ? ( bv_8_21_n89 ) : ( n21637 ) ;
assign n21639 =  ( n21494 ) ? ( bv_8_4_n516 ) : ( n21638 ) ;
assign n21640 =  ( n21492 ) ? ( bv_8_199_n216 ) : ( n21639 ) ;
assign n21641 =  ( n21490 ) ? ( bv_8_35_n696 ) : ( n21640 ) ;
assign n21642 =  ( n21488 ) ? ( bv_8_195_n232 ) : ( n21641 ) ;
assign n21643 =  ( n21486 ) ? ( bv_8_24_n448 ) : ( n21642 ) ;
assign n21644 =  ( n21484 ) ? ( bv_8_150_n201 ) : ( n21643 ) ;
assign n21645 =  ( n21482 ) ? ( bv_8_5_n492 ) : ( n21644 ) ;
assign n21646 =  ( n21480 ) ? ( bv_8_154_n368 ) : ( n21645 ) ;
assign n21647 =  ( n21478 ) ? ( bv_8_7_n105 ) : ( n21646 ) ;
assign n21648 =  ( n21476 ) ? ( bv_8_18_n628 ) : ( n21647 ) ;
assign n21649 =  ( n21474 ) ? ( bv_8_128_n450 ) : ( n21648 ) ;
assign n21650 =  ( n21472 ) ? ( bv_8_226_n119 ) : ( n21649 ) ;
assign n21651 =  ( n21470 ) ? ( bv_8_235_n83 ) : ( n21650 ) ;
assign n21652 =  ( n21468 ) ? ( bv_8_39_n132 ) : ( n21651 ) ;
assign n21653 =  ( n21466 ) ? ( bv_8_178_n292 ) : ( n21652 ) ;
assign n21654 =  ( n21464 ) ? ( bv_8_117_n484 ) : ( n21653 ) ;
assign n21655 =  ( n21462 ) ? ( bv_8_9_n57 ) : ( n21654 ) ;
assign n21656 =  ( n21460 ) ? ( bv_8_131_n440 ) : ( n21655 ) ;
assign n21657 =  ( n21458 ) ? ( bv_8_44_n5 ) : ( n21656 ) ;
assign n21658 =  ( n21456 ) ? ( bv_8_26_n53 ) : ( n21657 ) ;
assign n21659 =  ( n21454 ) ? ( bv_8_27_n642 ) : ( n21658 ) ;
assign n21660 =  ( n21452 ) ? ( bv_8_110_n294 ) : ( n21659 ) ;
assign n21661 =  ( n21450 ) ? ( bv_8_90_n25 ) : ( n21660 ) ;
assign n21662 =  ( n21448 ) ? ( bv_8_160_n350 ) : ( n21661 ) ;
assign n21663 =  ( n21446 ) ? ( bv_8_82_n578 ) : ( n21662 ) ;
assign n21664 =  ( n21444 ) ? ( bv_8_59_n382 ) : ( n21663 ) ;
assign n21665 =  ( n21442 ) ? ( bv_8_214_n164 ) : ( n21664 ) ;
assign n21666 =  ( n21440 ) ? ( bv_8_179_n289 ) : ( n21665 ) ;
assign n21667 =  ( n21438 ) ? ( bv_8_41_n29 ) : ( n21666 ) ;
assign n21668 =  ( n21436 ) ? ( bv_8_227_n115 ) : ( n21667 ) ;
assign n21669 =  ( n21434 ) ? ( bv_8_47_n652 ) : ( n21668 ) ;
assign n21670 =  ( n21432 ) ? ( bv_8_132_n41 ) : ( n21669 ) ;
assign n21671 =  ( n21430 ) ? ( bv_8_83_n575 ) : ( n21670 ) ;
assign n21672 =  ( n21428 ) ? ( bv_8_209_n182 ) : ( n21671 ) ;
assign n21673 =  ( n21426 ) ? ( bv_8_0_n580 ) : ( n21672 ) ;
assign n21674 =  ( n21424 ) ? ( bv_8_237_n75 ) : ( n21673 ) ;
assign n21675 =  ( n21422 ) ? ( bv_8_32_n463 ) : ( n21674 ) ;
assign n21676 =  ( n21420 ) ? ( bv_8_252_n15 ) : ( n21675 ) ;
assign n21677 =  ( n21418 ) ? ( bv_8_177_n283 ) : ( n21676 ) ;
assign n21678 =  ( n21416 ) ? ( bv_8_91_n555 ) : ( n21677 ) ;
assign n21679 =  ( n21414 ) ? ( bv_8_106_n155 ) : ( n21678 ) ;
assign n21680 =  ( n21412 ) ? ( bv_8_203_n203 ) : ( n21679 ) ;
assign n21681 =  ( n21410 ) ? ( bv_8_190_n250 ) : ( n21680 ) ;
assign n21682 =  ( n21408 ) ? ( bv_8_57_n312 ) : ( n21681 ) ;
assign n21683 =  ( n21406 ) ? ( bv_8_74_n237 ) : ( n21682 ) ;
assign n21684 =  ( n21404 ) ? ( bv_8_76_n596 ) : ( n21683 ) ;
assign n21685 =  ( n21402 ) ? ( bv_8_88_n562 ) : ( n21684 ) ;
assign n21686 =  ( n21400 ) ? ( bv_8_207_n188 ) : ( n21685 ) ;
assign n21687 =  ( n21398 ) ? ( bv_8_208_n37 ) : ( n21686 ) ;
assign n21688 =  ( n21396 ) ? ( bv_8_239_n67 ) : ( n21687 ) ;
assign n21689 =  ( n21394 ) ? ( bv_8_170_n77 ) : ( n21688 ) ;
assign n21690 =  ( n21392 ) ? ( bv_8_251_n19 ) : ( n21689 ) ;
assign n21691 =  ( n21390 ) ? ( bv_8_67_n318 ) : ( n21690 ) ;
assign n21692 =  ( n21388 ) ? ( bv_8_77_n593 ) : ( n21691 ) ;
assign n21693 =  ( n21386 ) ? ( bv_8_51_n101 ) : ( n21692 ) ;
assign n21694 =  ( n21384 ) ? ( bv_8_133_n434 ) : ( n21693 ) ;
assign n21695 =  ( n21382 ) ? ( bv_8_69_n612 ) : ( n21694 ) ;
assign n21696 =  ( n21380 ) ? ( bv_8_249_n27 ) : ( n21695 ) ;
assign n21697 =  ( n21378 ) ? ( bv_8_2_n751 ) : ( n21696 ) ;
assign n21698 =  ( n21376 ) ? ( bv_8_127_n453 ) : ( n21697 ) ;
assign n21699 =  ( n21374 ) ? ( bv_8_80_n73 ) : ( n21698 ) ;
assign n21700 =  ( n21372 ) ? ( bv_8_60_n93 ) : ( n21699 ) ;
assign n21701 =  ( n21370 ) ? ( bv_8_159_n323 ) : ( n21700 ) ;
assign n21702 =  ( n21368 ) ? ( bv_8_168_n13 ) : ( n21701 ) ;
assign n21703 =  ( n21366 ) ? ( bv_8_81_n582 ) : ( n21702 ) ;
assign n21704 =  ( n21364 ) ? ( bv_8_163_n339 ) : ( n21703 ) ;
assign n21705 =  ( n21362 ) ? ( bv_8_64_n573 ) : ( n21704 ) ;
assign n21706 =  ( n21360 ) ? ( bv_8_143_n403 ) : ( n21705 ) ;
assign n21707 =  ( n21358 ) ? ( bv_8_146_n337 ) : ( n21706 ) ;
assign n21708 =  ( n21356 ) ? ( bv_8_157_n359 ) : ( n21707 ) ;
assign n21709 =  ( n21354 ) ? ( bv_8_56_n230 ) : ( n21708 ) ;
assign n21710 =  ( n21352 ) ? ( bv_8_245_n43 ) : ( n21709 ) ;
assign n21711 =  ( n21350 ) ? ( bv_8_188_n257 ) : ( n21710 ) ;
assign n21712 =  ( n21348 ) ? ( bv_8_182_n277 ) : ( n21711 ) ;
assign n21713 =  ( n21346 ) ? ( bv_8_218_n150 ) : ( n21712 ) ;
assign n21714 =  ( n21344 ) ? ( bv_8_33_n486 ) : ( n21713 ) ;
assign n21715 =  ( n21342 ) ? ( bv_8_16_n248 ) : ( n21714 ) ;
assign n21716 =  ( n21340 ) ? ( bv_8_255_n3 ) : ( n21715 ) ;
assign n21717 =  ( n21338 ) ? ( bv_8_243_n51 ) : ( n21716 ) ;
assign n21718 =  ( n21336 ) ? ( bv_8_210_n113 ) : ( n21717 ) ;
assign n21719 =  ( n21334 ) ? ( bv_8_205_n196 ) : ( n21718 ) ;
assign n21720 =  ( n21332 ) ? ( bv_8_12_n333 ) : ( n21719 ) ;
assign n21721 =  ( n21330 ) ? ( bv_8_19_n588 ) : ( n21720 ) ;
assign n21722 =  ( n21328 ) ? ( bv_8_236_n79 ) : ( n21721 ) ;
assign n21723 =  ( n21326 ) ? ( bv_8_95_n545 ) : ( n21722 ) ;
assign n21724 =  ( n21324 ) ? ( bv_8_151_n218 ) : ( n21723 ) ;
assign n21725 =  ( n21322 ) ? ( bv_8_68_n390 ) : ( n21724 ) ;
assign n21726 =  ( n21320 ) ? ( bv_8_23_n144 ) : ( n21725 ) ;
assign n21727 =  ( n21318 ) ? ( bv_8_196_n228 ) : ( n21726 ) ;
assign n21728 =  ( n21316 ) ? ( bv_8_167_n325 ) : ( n21727 ) ;
assign n21729 =  ( n21314 ) ? ( bv_8_126_n456 ) : ( n21728 ) ;
assign n21730 =  ( n21312 ) ? ( bv_8_61_n634 ) : ( n21729 ) ;
assign n21731 =  ( n21310 ) ? ( bv_8_100_n348 ) : ( n21730 ) ;
assign n21732 =  ( n21308 ) ? ( bv_8_93_n498 ) : ( n21731 ) ;
assign n21733 =  ( n21306 ) ? ( bv_8_25_n399 ) : ( n21732 ) ;
assign n21734 =  ( n21304 ) ? ( bv_8_115_n222 ) : ( n21733 ) ;
assign n21735 =  ( n21302 ) ? ( bv_8_96_n542 ) : ( n21734 ) ;
assign n21736 =  ( n21300 ) ? ( bv_8_129_n446 ) : ( n21735 ) ;
assign n21737 =  ( n21298 ) ? ( bv_8_79_n538 ) : ( n21736 ) ;
assign n21738 =  ( n21296 ) ? ( bv_8_220_n142 ) : ( n21737 ) ;
assign n21739 =  ( n21294 ) ? ( bv_8_34_n117 ) : ( n21738 ) ;
assign n21740 =  ( n21292 ) ? ( bv_8_42_n672 ) : ( n21739 ) ;
assign n21741 =  ( n21290 ) ? ( bv_8_144_n173 ) : ( n21740 ) ;
assign n21742 =  ( n21288 ) ? ( bv_8_136_n425 ) : ( n21741 ) ;
assign n21743 =  ( n21286 ) ? ( bv_8_70_n609 ) : ( n21742 ) ;
assign n21744 =  ( n21284 ) ? ( bv_8_238_n71 ) : ( n21743 ) ;
assign n21745 =  ( n21282 ) ? ( bv_8_184_n270 ) : ( n21744 ) ;
assign n21746 =  ( n21280 ) ? ( bv_8_20_n341 ) : ( n21745 ) ;
assign n21747 =  ( n21278 ) ? ( bv_8_222_n134 ) : ( n21746 ) ;
assign n21748 =  ( n21276 ) ? ( bv_8_94_n548 ) : ( n21747 ) ;
assign n21749 =  ( n21274 ) ? ( bv_8_11_n379 ) : ( n21748 ) ;
assign n21750 =  ( n21272 ) ? ( bv_8_219_n146 ) : ( n21749 ) ;
assign n21751 =  ( n21270 ) ? ( bv_8_224_n126 ) : ( n21750 ) ;
assign n21752 =  ( n21268 ) ? ( bv_8_50_n408 ) : ( n21751 ) ;
assign n21753 =  ( n21266 ) ? ( bv_8_58_n136 ) : ( n21752 ) ;
assign n21754 =  ( n21264 ) ? ( bv_8_10_n655 ) : ( n21753 ) ;
assign n21755 =  ( n21262 ) ? ( bv_8_73_n275 ) : ( n21754 ) ;
assign n21756 =  ( n21260 ) ? ( bv_8_6_n169 ) : ( n21755 ) ;
assign n21757 =  ( n21258 ) ? ( bv_8_36_n645 ) : ( n21756 ) ;
assign n21758 =  ( n21256 ) ? ( bv_8_92_n234 ) : ( n21757 ) ;
assign n21759 =  ( n21254 ) ? ( bv_8_194_n159 ) : ( n21758 ) ;
assign n21760 =  ( n21252 ) ? ( bv_8_211_n175 ) : ( n21759 ) ;
assign n21761 =  ( n21250 ) ? ( bv_8_172_n268 ) : ( n21760 ) ;
assign n21762 =  ( n21248 ) ? ( bv_8_98_n536 ) : ( n21761 ) ;
assign n21763 =  ( n21246 ) ? ( bv_8_145_n397 ) : ( n21762 ) ;
assign n21764 =  ( n21244 ) ? ( bv_8_149_n384 ) : ( n21763 ) ;
assign n21765 =  ( n21242 ) ? ( bv_8_228_n111 ) : ( n21764 ) ;
assign n21766 =  ( n21240 ) ? ( bv_8_121_n470 ) : ( n21765 ) ;
assign n21767 =  ( n21238 ) ? ( bv_8_231_n99 ) : ( n21766 ) ;
assign n21768 =  ( n21236 ) ? ( bv_8_200_n213 ) : ( n21767 ) ;
assign n21769 =  ( n21234 ) ? ( bv_8_55_n650 ) : ( n21768 ) ;
assign n21770 =  ( n21232 ) ? ( bv_8_109_n9 ) : ( n21769 ) ;
assign n21771 =  ( n21230 ) ? ( bv_8_141_n410 ) : ( n21770 ) ;
assign n21772 =  ( n21228 ) ? ( bv_8_213_n167 ) : ( n21771 ) ;
assign n21773 =  ( n21226 ) ? ( bv_8_78_n590 ) : ( n21772 ) ;
assign n21774 =  ( n21224 ) ? ( bv_8_169_n109 ) : ( n21773 ) ;
assign n21775 =  ( n21222 ) ? ( bv_8_108_n510 ) : ( n21774 ) ;
assign n21776 =  ( n21220 ) ? ( bv_8_86_n567 ) : ( n21775 ) ;
assign n21777 =  ( n21218 ) ? ( bv_8_244_n47 ) : ( n21776 ) ;
assign n21778 =  ( n21216 ) ? ( bv_8_234_n87 ) : ( n21777 ) ;
assign n21779 =  ( n21214 ) ? ( bv_8_101_n49 ) : ( n21778 ) ;
assign n21780 =  ( n21212 ) ? ( bv_8_122_n416 ) : ( n21779 ) ;
assign n21781 =  ( n21210 ) ? ( bv_8_174_n152 ) : ( n21780 ) ;
assign n21782 =  ( n21208 ) ? ( bv_8_8_n669 ) : ( n21781 ) ;
assign n21783 =  ( n21206 ) ? ( bv_8_186_n263 ) : ( n21782 ) ;
assign n21784 =  ( n21204 ) ? ( bv_8_120_n474 ) : ( n21783 ) ;
assign n21785 =  ( n21202 ) ? ( bv_8_37_n506 ) : ( n21784 ) ;
assign n21786 =  ( n21200 ) ? ( bv_8_46_n429 ) : ( n21785 ) ;
assign n21787 =  ( n21198 ) ? ( bv_8_28_n162 ) : ( n21786 ) ;
assign n21788 =  ( n21196 ) ? ( bv_8_166_n328 ) : ( n21787 ) ;
assign n21789 =  ( n21194 ) ? ( bv_8_180_n285 ) : ( n21788 ) ;
assign n21790 =  ( n21192 ) ? ( bv_8_198_n220 ) : ( n21789 ) ;
assign n21791 =  ( n21190 ) ? ( bv_8_232_n95 ) : ( n21790 ) ;
assign n21792 =  ( n21188 ) ? ( bv_8_221_n138 ) : ( n21791 ) ;
assign n21793 =  ( n21186 ) ? ( bv_8_116_n345 ) : ( n21792 ) ;
assign n21794 =  ( n21184 ) ? ( bv_8_31_n705 ) : ( n21793 ) ;
assign n21795 =  ( n21182 ) ? ( bv_8_75_n503 ) : ( n21794 ) ;
assign n21796 =  ( n21180 ) ? ( bv_8_189_n254 ) : ( n21795 ) ;
assign n21797 =  ( n21178 ) ? ( bv_8_139_n297 ) : ( n21796 ) ;
assign n21798 =  ( n21176 ) ? ( bv_8_138_n418 ) : ( n21797 ) ;
assign n21799 =  ( n21174 ) ? ( bv_8_112_n482 ) : ( n21798 ) ;
assign n21800 =  ( n21172 ) ? ( bv_8_62_n205 ) : ( n21799 ) ;
assign n21801 =  ( n21170 ) ? ( bv_8_181_n281 ) : ( n21800 ) ;
assign n21802 =  ( n21168 ) ? ( bv_8_102_n527 ) : ( n21801 ) ;
assign n21803 =  ( n21166 ) ? ( bv_8_72_n330 ) : ( n21802 ) ;
assign n21804 =  ( n21164 ) ? ( bv_8_3_n65 ) : ( n21803 ) ;
assign n21805 =  ( n21162 ) ? ( bv_8_246_n39 ) : ( n21804 ) ;
assign n21806 =  ( n21160 ) ? ( bv_8_14_n648 ) : ( n21805 ) ;
assign n21807 =  ( n21158 ) ? ( bv_8_97_n198 ) : ( n21806 ) ;
assign n21808 =  ( n21156 ) ? ( bv_8_53_n436 ) : ( n21807 ) ;
assign n21809 =  ( n21154 ) ? ( bv_8_87_n226 ) : ( n21808 ) ;
assign n21810 =  ( n21152 ) ? ( bv_8_185_n266 ) : ( n21809 ) ;
assign n21811 =  ( n21150 ) ? ( bv_8_134_n431 ) : ( n21810 ) ;
assign n21812 =  ( n21148 ) ? ( bv_8_193_n239 ) : ( n21811 ) ;
assign n21813 =  ( n21146 ) ? ( bv_8_29_n625 ) : ( n21812 ) ;
assign n21814 =  ( n21144 ) ? ( bv_8_158_n355 ) : ( n21813 ) ;
assign n21815 =  ( n21142 ) ? ( bv_8_225_n123 ) : ( n21814 ) ;
assign n21816 =  ( n21140 ) ? ( bv_8_248_n31 ) : ( n21815 ) ;
assign n21817 =  ( n21138 ) ? ( bv_8_152_n374 ) : ( n21816 ) ;
assign n21818 =  ( n21136 ) ? ( bv_8_17_n525 ) : ( n21817 ) ;
assign n21819 =  ( n21134 ) ? ( bv_8_105_n148 ) : ( n21818 ) ;
assign n21820 =  ( n21132 ) ? ( bv_8_217_n128 ) : ( n21819 ) ;
assign n21821 =  ( n21130 ) ? ( bv_8_142_n406 ) : ( n21820 ) ;
assign n21822 =  ( n21128 ) ? ( bv_8_148_n388 ) : ( n21821 ) ;
assign n21823 =  ( n21126 ) ? ( bv_8_155_n364 ) : ( n21822 ) ;
assign n21824 =  ( n21124 ) ? ( bv_8_30_n21 ) : ( n21823 ) ;
assign n21825 =  ( n21122 ) ? ( bv_8_135_n81 ) : ( n21824 ) ;
assign n21826 =  ( n21120 ) ? ( bv_8_233_n91 ) : ( n21825 ) ;
assign n21827 =  ( n21118 ) ? ( bv_8_206_n192 ) : ( n21826 ) ;
assign n21828 =  ( n21116 ) ? ( bv_8_85_n423 ) : ( n21827 ) ;
assign n21829 =  ( n21114 ) ? ( bv_8_40_n366 ) : ( n21828 ) ;
assign n21830 =  ( n21112 ) ? ( bv_8_223_n130 ) : ( n21829 ) ;
assign n21831 =  ( n21110 ) ? ( bv_8_140_n376 ) : ( n21830 ) ;
assign n21832 =  ( n21108 ) ? ( bv_8_161_n211 ) : ( n21831 ) ;
assign n21833 =  ( n21106 ) ? ( bv_8_137_n421 ) : ( n21832 ) ;
assign n21834 =  ( n21104 ) ? ( bv_8_13_n194 ) : ( n21833 ) ;
assign n21835 =  ( n21102 ) ? ( bv_8_191_n246 ) : ( n21834 ) ;
assign n21836 =  ( n21100 ) ? ( bv_8_230_n103 ) : ( n21835 ) ;
assign n21837 =  ( n21098 ) ? ( bv_8_66_n466 ) : ( n21836 ) ;
assign n21838 =  ( n21096 ) ? ( bv_8_104_n520 ) : ( n21837 ) ;
assign n21839 =  ( n21094 ) ? ( bv_8_65_n623 ) : ( n21838 ) ;
assign n21840 =  ( n21092 ) ? ( bv_8_153_n140 ) : ( n21839 ) ;
assign n21841 =  ( n21090 ) ? ( bv_8_45_n97 ) : ( n21840 ) ;
assign n21842 =  ( n21088 ) ? ( bv_8_15_n190 ) : ( n21841 ) ;
assign n21843 =  ( n21086 ) ? ( bv_8_176_n299 ) : ( n21842 ) ;
assign n21844 =  ( n21084 ) ? ( bv_8_84_n386 ) : ( n21843 ) ;
assign n21845 =  ( n21082 ) ? ( bv_8_187_n260 ) : ( n21844 ) ;
assign n21846 =  ( n21080 ) ? ( bv_8_22_n357 ) : ( n21845 ) ;
assign n21847 =  ( n21078 ) ^ ( n21846 )  ;
assign n21848 = state_in[31:24] ;
assign n21849 =  ( n21848 ) == ( bv_8_255_n3 )  ;
assign n21850 = state_in[31:24] ;
assign n21851 =  ( n21850 ) == ( bv_8_254_n7 )  ;
assign n21852 = state_in[31:24] ;
assign n21853 =  ( n21852 ) == ( bv_8_253_n11 )  ;
assign n21854 = state_in[31:24] ;
assign n21855 =  ( n21854 ) == ( bv_8_252_n15 )  ;
assign n21856 = state_in[31:24] ;
assign n21857 =  ( n21856 ) == ( bv_8_251_n19 )  ;
assign n21858 = state_in[31:24] ;
assign n21859 =  ( n21858 ) == ( bv_8_250_n23 )  ;
assign n21860 = state_in[31:24] ;
assign n21861 =  ( n21860 ) == ( bv_8_249_n27 )  ;
assign n21862 = state_in[31:24] ;
assign n21863 =  ( n21862 ) == ( bv_8_248_n31 )  ;
assign n21864 = state_in[31:24] ;
assign n21865 =  ( n21864 ) == ( bv_8_247_n35 )  ;
assign n21866 = state_in[31:24] ;
assign n21867 =  ( n21866 ) == ( bv_8_246_n39 )  ;
assign n21868 = state_in[31:24] ;
assign n21869 =  ( n21868 ) == ( bv_8_245_n43 )  ;
assign n21870 = state_in[31:24] ;
assign n21871 =  ( n21870 ) == ( bv_8_244_n47 )  ;
assign n21872 = state_in[31:24] ;
assign n21873 =  ( n21872 ) == ( bv_8_243_n51 )  ;
assign n21874 = state_in[31:24] ;
assign n21875 =  ( n21874 ) == ( bv_8_242_n55 )  ;
assign n21876 = state_in[31:24] ;
assign n21877 =  ( n21876 ) == ( bv_8_241_n59 )  ;
assign n21878 = state_in[31:24] ;
assign n21879 =  ( n21878 ) == ( bv_8_240_n63 )  ;
assign n21880 = state_in[31:24] ;
assign n21881 =  ( n21880 ) == ( bv_8_239_n67 )  ;
assign n21882 = state_in[31:24] ;
assign n21883 =  ( n21882 ) == ( bv_8_238_n71 )  ;
assign n21884 = state_in[31:24] ;
assign n21885 =  ( n21884 ) == ( bv_8_237_n75 )  ;
assign n21886 = state_in[31:24] ;
assign n21887 =  ( n21886 ) == ( bv_8_236_n79 )  ;
assign n21888 = state_in[31:24] ;
assign n21889 =  ( n21888 ) == ( bv_8_235_n83 )  ;
assign n21890 = state_in[31:24] ;
assign n21891 =  ( n21890 ) == ( bv_8_234_n87 )  ;
assign n21892 = state_in[31:24] ;
assign n21893 =  ( n21892 ) == ( bv_8_233_n91 )  ;
assign n21894 = state_in[31:24] ;
assign n21895 =  ( n21894 ) == ( bv_8_232_n95 )  ;
assign n21896 = state_in[31:24] ;
assign n21897 =  ( n21896 ) == ( bv_8_231_n99 )  ;
assign n21898 = state_in[31:24] ;
assign n21899 =  ( n21898 ) == ( bv_8_230_n103 )  ;
assign n21900 = state_in[31:24] ;
assign n21901 =  ( n21900 ) == ( bv_8_229_n107 )  ;
assign n21902 = state_in[31:24] ;
assign n21903 =  ( n21902 ) == ( bv_8_228_n111 )  ;
assign n21904 = state_in[31:24] ;
assign n21905 =  ( n21904 ) == ( bv_8_227_n115 )  ;
assign n21906 = state_in[31:24] ;
assign n21907 =  ( n21906 ) == ( bv_8_226_n119 )  ;
assign n21908 = state_in[31:24] ;
assign n21909 =  ( n21908 ) == ( bv_8_225_n123 )  ;
assign n21910 = state_in[31:24] ;
assign n21911 =  ( n21910 ) == ( bv_8_224_n126 )  ;
assign n21912 = state_in[31:24] ;
assign n21913 =  ( n21912 ) == ( bv_8_223_n130 )  ;
assign n21914 = state_in[31:24] ;
assign n21915 =  ( n21914 ) == ( bv_8_222_n134 )  ;
assign n21916 = state_in[31:24] ;
assign n21917 =  ( n21916 ) == ( bv_8_221_n138 )  ;
assign n21918 = state_in[31:24] ;
assign n21919 =  ( n21918 ) == ( bv_8_220_n142 )  ;
assign n21920 = state_in[31:24] ;
assign n21921 =  ( n21920 ) == ( bv_8_219_n146 )  ;
assign n21922 = state_in[31:24] ;
assign n21923 =  ( n21922 ) == ( bv_8_218_n150 )  ;
assign n21924 = state_in[31:24] ;
assign n21925 =  ( n21924 ) == ( bv_8_217_n128 )  ;
assign n21926 = state_in[31:24] ;
assign n21927 =  ( n21926 ) == ( bv_8_216_n157 )  ;
assign n21928 = state_in[31:24] ;
assign n21929 =  ( n21928 ) == ( bv_8_215_n45 )  ;
assign n21930 = state_in[31:24] ;
assign n21931 =  ( n21930 ) == ( bv_8_214_n164 )  ;
assign n21932 = state_in[31:24] ;
assign n21933 =  ( n21932 ) == ( bv_8_213_n167 )  ;
assign n21934 = state_in[31:24] ;
assign n21935 =  ( n21934 ) == ( bv_8_212_n171 )  ;
assign n21936 = state_in[31:24] ;
assign n21937 =  ( n21936 ) == ( bv_8_211_n175 )  ;
assign n21938 = state_in[31:24] ;
assign n21939 =  ( n21938 ) == ( bv_8_210_n113 )  ;
assign n21940 = state_in[31:24] ;
assign n21941 =  ( n21940 ) == ( bv_8_209_n182 )  ;
assign n21942 = state_in[31:24] ;
assign n21943 =  ( n21942 ) == ( bv_8_208_n37 )  ;
assign n21944 = state_in[31:24] ;
assign n21945 =  ( n21944 ) == ( bv_8_207_n188 )  ;
assign n21946 = state_in[31:24] ;
assign n21947 =  ( n21946 ) == ( bv_8_206_n192 )  ;
assign n21948 = state_in[31:24] ;
assign n21949 =  ( n21948 ) == ( bv_8_205_n196 )  ;
assign n21950 = state_in[31:24] ;
assign n21951 =  ( n21950 ) == ( bv_8_204_n177 )  ;
assign n21952 = state_in[31:24] ;
assign n21953 =  ( n21952 ) == ( bv_8_203_n203 )  ;
assign n21954 = state_in[31:24] ;
assign n21955 =  ( n21954 ) == ( bv_8_202_n207 )  ;
assign n21956 = state_in[31:24] ;
assign n21957 =  ( n21956 ) == ( bv_8_201_n85 )  ;
assign n21958 = state_in[31:24] ;
assign n21959 =  ( n21958 ) == ( bv_8_200_n213 )  ;
assign n21960 = state_in[31:24] ;
assign n21961 =  ( n21960 ) == ( bv_8_199_n216 )  ;
assign n21962 = state_in[31:24] ;
assign n21963 =  ( n21962 ) == ( bv_8_198_n220 )  ;
assign n21964 = state_in[31:24] ;
assign n21965 =  ( n21964 ) == ( bv_8_197_n224 )  ;
assign n21966 = state_in[31:24] ;
assign n21967 =  ( n21966 ) == ( bv_8_196_n228 )  ;
assign n21968 = state_in[31:24] ;
assign n21969 =  ( n21968 ) == ( bv_8_195_n232 )  ;
assign n21970 = state_in[31:24] ;
assign n21971 =  ( n21970 ) == ( bv_8_194_n159 )  ;
assign n21972 = state_in[31:24] ;
assign n21973 =  ( n21972 ) == ( bv_8_193_n239 )  ;
assign n21974 = state_in[31:24] ;
assign n21975 =  ( n21974 ) == ( bv_8_192_n242 )  ;
assign n21976 = state_in[31:24] ;
assign n21977 =  ( n21976 ) == ( bv_8_191_n246 )  ;
assign n21978 = state_in[31:24] ;
assign n21979 =  ( n21978 ) == ( bv_8_190_n250 )  ;
assign n21980 = state_in[31:24] ;
assign n21981 =  ( n21980 ) == ( bv_8_189_n254 )  ;
assign n21982 = state_in[31:24] ;
assign n21983 =  ( n21982 ) == ( bv_8_188_n257 )  ;
assign n21984 = state_in[31:24] ;
assign n21985 =  ( n21984 ) == ( bv_8_187_n260 )  ;
assign n21986 = state_in[31:24] ;
assign n21987 =  ( n21986 ) == ( bv_8_186_n263 )  ;
assign n21988 = state_in[31:24] ;
assign n21989 =  ( n21988 ) == ( bv_8_185_n266 )  ;
assign n21990 = state_in[31:24] ;
assign n21991 =  ( n21990 ) == ( bv_8_184_n270 )  ;
assign n21992 = state_in[31:24] ;
assign n21993 =  ( n21992 ) == ( bv_8_183_n273 )  ;
assign n21994 = state_in[31:24] ;
assign n21995 =  ( n21994 ) == ( bv_8_182_n277 )  ;
assign n21996 = state_in[31:24] ;
assign n21997 =  ( n21996 ) == ( bv_8_181_n281 )  ;
assign n21998 = state_in[31:24] ;
assign n21999 =  ( n21998 ) == ( bv_8_180_n285 )  ;
assign n22000 = state_in[31:24] ;
assign n22001 =  ( n22000 ) == ( bv_8_179_n289 )  ;
assign n22002 = state_in[31:24] ;
assign n22003 =  ( n22002 ) == ( bv_8_178_n292 )  ;
assign n22004 = state_in[31:24] ;
assign n22005 =  ( n22004 ) == ( bv_8_177_n283 )  ;
assign n22006 = state_in[31:24] ;
assign n22007 =  ( n22006 ) == ( bv_8_176_n299 )  ;
assign n22008 = state_in[31:24] ;
assign n22009 =  ( n22008 ) == ( bv_8_175_n302 )  ;
assign n22010 = state_in[31:24] ;
assign n22011 =  ( n22010 ) == ( bv_8_174_n152 )  ;
assign n22012 = state_in[31:24] ;
assign n22013 =  ( n22012 ) == ( bv_8_173_n307 )  ;
assign n22014 = state_in[31:24] ;
assign n22015 =  ( n22014 ) == ( bv_8_172_n268 )  ;
assign n22016 = state_in[31:24] ;
assign n22017 =  ( n22016 ) == ( bv_8_171_n314 )  ;
assign n22018 = state_in[31:24] ;
assign n22019 =  ( n22018 ) == ( bv_8_170_n77 )  ;
assign n22020 = state_in[31:24] ;
assign n22021 =  ( n22020 ) == ( bv_8_169_n109 )  ;
assign n22022 = state_in[31:24] ;
assign n22023 =  ( n22022 ) == ( bv_8_168_n13 )  ;
assign n22024 = state_in[31:24] ;
assign n22025 =  ( n22024 ) == ( bv_8_167_n325 )  ;
assign n22026 = state_in[31:24] ;
assign n22027 =  ( n22026 ) == ( bv_8_166_n328 )  ;
assign n22028 = state_in[31:24] ;
assign n22029 =  ( n22028 ) == ( bv_8_165_n69 )  ;
assign n22030 = state_in[31:24] ;
assign n22031 =  ( n22030 ) == ( bv_8_164_n335 )  ;
assign n22032 = state_in[31:24] ;
assign n22033 =  ( n22032 ) == ( bv_8_163_n339 )  ;
assign n22034 = state_in[31:24] ;
assign n22035 =  ( n22034 ) == ( bv_8_162_n343 )  ;
assign n22036 = state_in[31:24] ;
assign n22037 =  ( n22036 ) == ( bv_8_161_n211 )  ;
assign n22038 = state_in[31:24] ;
assign n22039 =  ( n22038 ) == ( bv_8_160_n350 )  ;
assign n22040 = state_in[31:24] ;
assign n22041 =  ( n22040 ) == ( bv_8_159_n323 )  ;
assign n22042 = state_in[31:24] ;
assign n22043 =  ( n22042 ) == ( bv_8_158_n355 )  ;
assign n22044 = state_in[31:24] ;
assign n22045 =  ( n22044 ) == ( bv_8_157_n359 )  ;
assign n22046 = state_in[31:24] ;
assign n22047 =  ( n22046 ) == ( bv_8_156_n279 )  ;
assign n22048 = state_in[31:24] ;
assign n22049 =  ( n22048 ) == ( bv_8_155_n364 )  ;
assign n22050 = state_in[31:24] ;
assign n22051 =  ( n22050 ) == ( bv_8_154_n368 )  ;
assign n22052 = state_in[31:24] ;
assign n22053 =  ( n22052 ) == ( bv_8_153_n140 )  ;
assign n22054 = state_in[31:24] ;
assign n22055 =  ( n22054 ) == ( bv_8_152_n374 )  ;
assign n22056 = state_in[31:24] ;
assign n22057 =  ( n22056 ) == ( bv_8_151_n218 )  ;
assign n22058 = state_in[31:24] ;
assign n22059 =  ( n22058 ) == ( bv_8_150_n201 )  ;
assign n22060 = state_in[31:24] ;
assign n22061 =  ( n22060 ) == ( bv_8_149_n384 )  ;
assign n22062 = state_in[31:24] ;
assign n22063 =  ( n22062 ) == ( bv_8_148_n388 )  ;
assign n22064 = state_in[31:24] ;
assign n22065 =  ( n22064 ) == ( bv_8_147_n392 )  ;
assign n22066 = state_in[31:24] ;
assign n22067 =  ( n22066 ) == ( bv_8_146_n337 )  ;
assign n22068 = state_in[31:24] ;
assign n22069 =  ( n22068 ) == ( bv_8_145_n397 )  ;
assign n22070 = state_in[31:24] ;
assign n22071 =  ( n22070 ) == ( bv_8_144_n173 )  ;
assign n22072 = state_in[31:24] ;
assign n22073 =  ( n22072 ) == ( bv_8_143_n403 )  ;
assign n22074 = state_in[31:24] ;
assign n22075 =  ( n22074 ) == ( bv_8_142_n406 )  ;
assign n22076 = state_in[31:24] ;
assign n22077 =  ( n22076 ) == ( bv_8_141_n410 )  ;
assign n22078 = state_in[31:24] ;
assign n22079 =  ( n22078 ) == ( bv_8_140_n376 )  ;
assign n22080 = state_in[31:24] ;
assign n22081 =  ( n22080 ) == ( bv_8_139_n297 )  ;
assign n22082 = state_in[31:24] ;
assign n22083 =  ( n22082 ) == ( bv_8_138_n418 )  ;
assign n22084 = state_in[31:24] ;
assign n22085 =  ( n22084 ) == ( bv_8_137_n421 )  ;
assign n22086 = state_in[31:24] ;
assign n22087 =  ( n22086 ) == ( bv_8_136_n425 )  ;
assign n22088 = state_in[31:24] ;
assign n22089 =  ( n22088 ) == ( bv_8_135_n81 )  ;
assign n22090 = state_in[31:24] ;
assign n22091 =  ( n22090 ) == ( bv_8_134_n431 )  ;
assign n22092 = state_in[31:24] ;
assign n22093 =  ( n22092 ) == ( bv_8_133_n434 )  ;
assign n22094 = state_in[31:24] ;
assign n22095 =  ( n22094 ) == ( bv_8_132_n41 )  ;
assign n22096 = state_in[31:24] ;
assign n22097 =  ( n22096 ) == ( bv_8_131_n440 )  ;
assign n22098 = state_in[31:24] ;
assign n22099 =  ( n22098 ) == ( bv_8_130_n33 )  ;
assign n22100 = state_in[31:24] ;
assign n22101 =  ( n22100 ) == ( bv_8_129_n446 )  ;
assign n22102 = state_in[31:24] ;
assign n22103 =  ( n22102 ) == ( bv_8_128_n450 )  ;
assign n22104 = state_in[31:24] ;
assign n22105 =  ( n22104 ) == ( bv_8_127_n453 )  ;
assign n22106 = state_in[31:24] ;
assign n22107 =  ( n22106 ) == ( bv_8_126_n456 )  ;
assign n22108 = state_in[31:24] ;
assign n22109 =  ( n22108 ) == ( bv_8_125_n459 )  ;
assign n22110 = state_in[31:24] ;
assign n22111 =  ( n22110 ) == ( bv_8_124_n184 )  ;
assign n22112 = state_in[31:24] ;
assign n22113 =  ( n22112 ) == ( bv_8_123_n17 )  ;
assign n22114 = state_in[31:24] ;
assign n22115 =  ( n22114 ) == ( bv_8_122_n416 )  ;
assign n22116 = state_in[31:24] ;
assign n22117 =  ( n22116 ) == ( bv_8_121_n470 )  ;
assign n22118 = state_in[31:24] ;
assign n22119 =  ( n22118 ) == ( bv_8_120_n474 )  ;
assign n22120 = state_in[31:24] ;
assign n22121 =  ( n22120 ) == ( bv_8_119_n472 )  ;
assign n22122 = state_in[31:24] ;
assign n22123 =  ( n22122 ) == ( bv_8_118_n480 )  ;
assign n22124 = state_in[31:24] ;
assign n22125 =  ( n22124 ) == ( bv_8_117_n484 )  ;
assign n22126 = state_in[31:24] ;
assign n22127 =  ( n22126 ) == ( bv_8_116_n345 )  ;
assign n22128 = state_in[31:24] ;
assign n22129 =  ( n22128 ) == ( bv_8_115_n222 )  ;
assign n22130 = state_in[31:24] ;
assign n22131 =  ( n22130 ) == ( bv_8_114_n494 )  ;
assign n22132 = state_in[31:24] ;
assign n22133 =  ( n22132 ) == ( bv_8_113_n180 )  ;
assign n22134 = state_in[31:24] ;
assign n22135 =  ( n22134 ) == ( bv_8_112_n482 )  ;
assign n22136 = state_in[31:24] ;
assign n22137 =  ( n22136 ) == ( bv_8_111_n244 )  ;
assign n22138 = state_in[31:24] ;
assign n22139 =  ( n22138 ) == ( bv_8_110_n294 )  ;
assign n22140 = state_in[31:24] ;
assign n22141 =  ( n22140 ) == ( bv_8_109_n9 )  ;
assign n22142 = state_in[31:24] ;
assign n22143 =  ( n22142 ) == ( bv_8_108_n510 )  ;
assign n22144 = state_in[31:24] ;
assign n22145 =  ( n22144 ) == ( bv_8_107_n370 )  ;
assign n22146 = state_in[31:24] ;
assign n22147 =  ( n22146 ) == ( bv_8_106_n155 )  ;
assign n22148 = state_in[31:24] ;
assign n22149 =  ( n22148 ) == ( bv_8_105_n148 )  ;
assign n22150 = state_in[31:24] ;
assign n22151 =  ( n22150 ) == ( bv_8_104_n520 )  ;
assign n22152 = state_in[31:24] ;
assign n22153 =  ( n22152 ) == ( bv_8_103_n523 )  ;
assign n22154 = state_in[31:24] ;
assign n22155 =  ( n22154 ) == ( bv_8_102_n527 )  ;
assign n22156 = state_in[31:24] ;
assign n22157 =  ( n22156 ) == ( bv_8_101_n49 )  ;
assign n22158 = state_in[31:24] ;
assign n22159 =  ( n22158 ) == ( bv_8_100_n348 )  ;
assign n22160 = state_in[31:24] ;
assign n22161 =  ( n22160 ) == ( bv_8_99_n476 )  ;
assign n22162 = state_in[31:24] ;
assign n22163 =  ( n22162 ) == ( bv_8_98_n536 )  ;
assign n22164 = state_in[31:24] ;
assign n22165 =  ( n22164 ) == ( bv_8_97_n198 )  ;
assign n22166 = state_in[31:24] ;
assign n22167 =  ( n22166 ) == ( bv_8_96_n542 )  ;
assign n22168 = state_in[31:24] ;
assign n22169 =  ( n22168 ) == ( bv_8_95_n545 )  ;
assign n22170 = state_in[31:24] ;
assign n22171 =  ( n22170 ) == ( bv_8_94_n548 )  ;
assign n22172 = state_in[31:24] ;
assign n22173 =  ( n22172 ) == ( bv_8_93_n498 )  ;
assign n22174 = state_in[31:24] ;
assign n22175 =  ( n22174 ) == ( bv_8_92_n234 )  ;
assign n22176 = state_in[31:24] ;
assign n22177 =  ( n22176 ) == ( bv_8_91_n555 )  ;
assign n22178 = state_in[31:24] ;
assign n22179 =  ( n22178 ) == ( bv_8_90_n25 )  ;
assign n22180 = state_in[31:24] ;
assign n22181 =  ( n22180 ) == ( bv_8_89_n61 )  ;
assign n22182 = state_in[31:24] ;
assign n22183 =  ( n22182 ) == ( bv_8_88_n562 )  ;
assign n22184 = state_in[31:24] ;
assign n22185 =  ( n22184 ) == ( bv_8_87_n226 )  ;
assign n22186 = state_in[31:24] ;
assign n22187 =  ( n22186 ) == ( bv_8_86_n567 )  ;
assign n22188 = state_in[31:24] ;
assign n22189 =  ( n22188 ) == ( bv_8_85_n423 )  ;
assign n22190 = state_in[31:24] ;
assign n22191 =  ( n22190 ) == ( bv_8_84_n386 )  ;
assign n22192 = state_in[31:24] ;
assign n22193 =  ( n22192 ) == ( bv_8_83_n575 )  ;
assign n22194 = state_in[31:24] ;
assign n22195 =  ( n22194 ) == ( bv_8_82_n578 )  ;
assign n22196 = state_in[31:24] ;
assign n22197 =  ( n22196 ) == ( bv_8_81_n582 )  ;
assign n22198 = state_in[31:24] ;
assign n22199 =  ( n22198 ) == ( bv_8_80_n73 )  ;
assign n22200 = state_in[31:24] ;
assign n22201 =  ( n22200 ) == ( bv_8_79_n538 )  ;
assign n22202 = state_in[31:24] ;
assign n22203 =  ( n22202 ) == ( bv_8_78_n590 )  ;
assign n22204 = state_in[31:24] ;
assign n22205 =  ( n22204 ) == ( bv_8_77_n593 )  ;
assign n22206 = state_in[31:24] ;
assign n22207 =  ( n22206 ) == ( bv_8_76_n596 )  ;
assign n22208 = state_in[31:24] ;
assign n22209 =  ( n22208 ) == ( bv_8_75_n503 )  ;
assign n22210 = state_in[31:24] ;
assign n22211 =  ( n22210 ) == ( bv_8_74_n237 )  ;
assign n22212 = state_in[31:24] ;
assign n22213 =  ( n22212 ) == ( bv_8_73_n275 )  ;
assign n22214 = state_in[31:24] ;
assign n22215 =  ( n22214 ) == ( bv_8_72_n330 )  ;
assign n22216 = state_in[31:24] ;
assign n22217 =  ( n22216 ) == ( bv_8_71_n252 )  ;
assign n22218 = state_in[31:24] ;
assign n22219 =  ( n22218 ) == ( bv_8_70_n609 )  ;
assign n22220 = state_in[31:24] ;
assign n22221 =  ( n22220 ) == ( bv_8_69_n612 )  ;
assign n22222 = state_in[31:24] ;
assign n22223 =  ( n22222 ) == ( bv_8_68_n390 )  ;
assign n22224 = state_in[31:24] ;
assign n22225 =  ( n22224 ) == ( bv_8_67_n318 )  ;
assign n22226 = state_in[31:24] ;
assign n22227 =  ( n22226 ) == ( bv_8_66_n466 )  ;
assign n22228 = state_in[31:24] ;
assign n22229 =  ( n22228 ) == ( bv_8_65_n623 )  ;
assign n22230 = state_in[31:24] ;
assign n22231 =  ( n22230 ) == ( bv_8_64_n573 )  ;
assign n22232 = state_in[31:24] ;
assign n22233 =  ( n22232 ) == ( bv_8_63_n489 )  ;
assign n22234 = state_in[31:24] ;
assign n22235 =  ( n22234 ) == ( bv_8_62_n205 )  ;
assign n22236 = state_in[31:24] ;
assign n22237 =  ( n22236 ) == ( bv_8_61_n634 )  ;
assign n22238 = state_in[31:24] ;
assign n22239 =  ( n22238 ) == ( bv_8_60_n93 )  ;
assign n22240 = state_in[31:24] ;
assign n22241 =  ( n22240 ) == ( bv_8_59_n382 )  ;
assign n22242 = state_in[31:24] ;
assign n22243 =  ( n22242 ) == ( bv_8_58_n136 )  ;
assign n22244 = state_in[31:24] ;
assign n22245 =  ( n22244 ) == ( bv_8_57_n312 )  ;
assign n22246 = state_in[31:24] ;
assign n22247 =  ( n22246 ) == ( bv_8_56_n230 )  ;
assign n22248 = state_in[31:24] ;
assign n22249 =  ( n22248 ) == ( bv_8_55_n650 )  ;
assign n22250 = state_in[31:24] ;
assign n22251 =  ( n22250 ) == ( bv_8_54_n616 )  ;
assign n22252 = state_in[31:24] ;
assign n22253 =  ( n22252 ) == ( bv_8_53_n436 )  ;
assign n22254 = state_in[31:24] ;
assign n22255 =  ( n22254 ) == ( bv_8_52_n619 )  ;
assign n22256 = state_in[31:24] ;
assign n22257 =  ( n22256 ) == ( bv_8_51_n101 )  ;
assign n22258 = state_in[31:24] ;
assign n22259 =  ( n22258 ) == ( bv_8_50_n408 )  ;
assign n22260 = state_in[31:24] ;
assign n22261 =  ( n22260 ) == ( bv_8_49_n309 )  ;
assign n22262 = state_in[31:24] ;
assign n22263 =  ( n22262 ) == ( bv_8_48_n660 )  ;
assign n22264 = state_in[31:24] ;
assign n22265 =  ( n22264 ) == ( bv_8_47_n652 )  ;
assign n22266 = state_in[31:24] ;
assign n22267 =  ( n22266 ) == ( bv_8_46_n429 )  ;
assign n22268 = state_in[31:24] ;
assign n22269 =  ( n22268 ) == ( bv_8_45_n97 )  ;
assign n22270 = state_in[31:24] ;
assign n22271 =  ( n22270 ) == ( bv_8_44_n5 )  ;
assign n22272 = state_in[31:24] ;
assign n22273 =  ( n22272 ) == ( bv_8_43_n121 )  ;
assign n22274 = state_in[31:24] ;
assign n22275 =  ( n22274 ) == ( bv_8_42_n672 )  ;
assign n22276 = state_in[31:24] ;
assign n22277 =  ( n22276 ) == ( bv_8_41_n29 )  ;
assign n22278 = state_in[31:24] ;
assign n22279 =  ( n22278 ) == ( bv_8_40_n366 )  ;
assign n22280 = state_in[31:24] ;
assign n22281 =  ( n22280 ) == ( bv_8_39_n132 )  ;
assign n22282 = state_in[31:24] ;
assign n22283 =  ( n22282 ) == ( bv_8_38_n444 )  ;
assign n22284 = state_in[31:24] ;
assign n22285 =  ( n22284 ) == ( bv_8_37_n506 )  ;
assign n22286 = state_in[31:24] ;
assign n22287 =  ( n22286 ) == ( bv_8_36_n645 )  ;
assign n22288 = state_in[31:24] ;
assign n22289 =  ( n22288 ) == ( bv_8_35_n696 )  ;
assign n22290 = state_in[31:24] ;
assign n22291 =  ( n22290 ) == ( bv_8_34_n117 )  ;
assign n22292 = state_in[31:24] ;
assign n22293 =  ( n22292 ) == ( bv_8_33_n486 )  ;
assign n22294 = state_in[31:24] ;
assign n22295 =  ( n22294 ) == ( bv_8_32_n463 )  ;
assign n22296 = state_in[31:24] ;
assign n22297 =  ( n22296 ) == ( bv_8_31_n705 )  ;
assign n22298 = state_in[31:24] ;
assign n22299 =  ( n22298 ) == ( bv_8_30_n21 )  ;
assign n22300 = state_in[31:24] ;
assign n22301 =  ( n22300 ) == ( bv_8_29_n625 )  ;
assign n22302 = state_in[31:24] ;
assign n22303 =  ( n22302 ) == ( bv_8_28_n162 )  ;
assign n22304 = state_in[31:24] ;
assign n22305 =  ( n22304 ) == ( bv_8_27_n642 )  ;
assign n22306 = state_in[31:24] ;
assign n22307 =  ( n22306 ) == ( bv_8_26_n53 )  ;
assign n22308 = state_in[31:24] ;
assign n22309 =  ( n22308 ) == ( bv_8_25_n399 )  ;
assign n22310 = state_in[31:24] ;
assign n22311 =  ( n22310 ) == ( bv_8_24_n448 )  ;
assign n22312 = state_in[31:24] ;
assign n22313 =  ( n22312 ) == ( bv_8_23_n144 )  ;
assign n22314 = state_in[31:24] ;
assign n22315 =  ( n22314 ) == ( bv_8_22_n357 )  ;
assign n22316 = state_in[31:24] ;
assign n22317 =  ( n22316 ) == ( bv_8_21_n89 )  ;
assign n22318 = state_in[31:24] ;
assign n22319 =  ( n22318 ) == ( bv_8_20_n341 )  ;
assign n22320 = state_in[31:24] ;
assign n22321 =  ( n22320 ) == ( bv_8_19_n588 )  ;
assign n22322 = state_in[31:24] ;
assign n22323 =  ( n22322 ) == ( bv_8_18_n628 )  ;
assign n22324 = state_in[31:24] ;
assign n22325 =  ( n22324 ) == ( bv_8_17_n525 )  ;
assign n22326 = state_in[31:24] ;
assign n22327 =  ( n22326 ) == ( bv_8_16_n248 )  ;
assign n22328 = state_in[31:24] ;
assign n22329 =  ( n22328 ) == ( bv_8_15_n190 )  ;
assign n22330 = state_in[31:24] ;
assign n22331 =  ( n22330 ) == ( bv_8_14_n648 )  ;
assign n22332 = state_in[31:24] ;
assign n22333 =  ( n22332 ) == ( bv_8_13_n194 )  ;
assign n22334 = state_in[31:24] ;
assign n22335 =  ( n22334 ) == ( bv_8_12_n333 )  ;
assign n22336 = state_in[31:24] ;
assign n22337 =  ( n22336 ) == ( bv_8_11_n379 )  ;
assign n22338 = state_in[31:24] ;
assign n22339 =  ( n22338 ) == ( bv_8_10_n655 )  ;
assign n22340 = state_in[31:24] ;
assign n22341 =  ( n22340 ) == ( bv_8_9_n57 )  ;
assign n22342 = state_in[31:24] ;
assign n22343 =  ( n22342 ) == ( bv_8_8_n669 )  ;
assign n22344 = state_in[31:24] ;
assign n22345 =  ( n22344 ) == ( bv_8_7_n105 )  ;
assign n22346 = state_in[31:24] ;
assign n22347 =  ( n22346 ) == ( bv_8_6_n169 )  ;
assign n22348 = state_in[31:24] ;
assign n22349 =  ( n22348 ) == ( bv_8_5_n492 )  ;
assign n22350 = state_in[31:24] ;
assign n22351 =  ( n22350 ) == ( bv_8_4_n516 )  ;
assign n22352 = state_in[31:24] ;
assign n22353 =  ( n22352 ) == ( bv_8_3_n65 )  ;
assign n22354 = state_in[31:24] ;
assign n22355 =  ( n22354 ) == ( bv_8_2_n751 )  ;
assign n22356 = state_in[31:24] ;
assign n22357 =  ( n22356 ) == ( bv_8_1_n287 )  ;
assign n22358 = state_in[31:24] ;
assign n22359 =  ( n22358 ) == ( bv_8_0_n580 )  ;
assign n22360 =  ( n22359 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n22361 =  ( n22357 ) ? ( bv_8_248_n31 ) : ( n22360 ) ;
assign n22362 =  ( n22355 ) ? ( bv_8_238_n71 ) : ( n22361 ) ;
assign n22363 =  ( n22353 ) ? ( bv_8_246_n39 ) : ( n22362 ) ;
assign n22364 =  ( n22351 ) ? ( bv_8_255_n3 ) : ( n22363 ) ;
assign n22365 =  ( n22349 ) ? ( bv_8_214_n164 ) : ( n22364 ) ;
assign n22366 =  ( n22347 ) ? ( bv_8_222_n134 ) : ( n22365 ) ;
assign n22367 =  ( n22345 ) ? ( bv_8_145_n397 ) : ( n22366 ) ;
assign n22368 =  ( n22343 ) ? ( bv_8_96_n542 ) : ( n22367 ) ;
assign n22369 =  ( n22341 ) ? ( bv_8_2_n751 ) : ( n22368 ) ;
assign n22370 =  ( n22339 ) ? ( bv_8_206_n192 ) : ( n22369 ) ;
assign n22371 =  ( n22337 ) ? ( bv_8_86_n567 ) : ( n22370 ) ;
assign n22372 =  ( n22335 ) ? ( bv_8_231_n99 ) : ( n22371 ) ;
assign n22373 =  ( n22333 ) ? ( bv_8_181_n281 ) : ( n22372 ) ;
assign n22374 =  ( n22331 ) ? ( bv_8_77_n593 ) : ( n22373 ) ;
assign n22375 =  ( n22329 ) ? ( bv_8_236_n79 ) : ( n22374 ) ;
assign n22376 =  ( n22327 ) ? ( bv_8_143_n403 ) : ( n22375 ) ;
assign n22377 =  ( n22325 ) ? ( bv_8_31_n705 ) : ( n22376 ) ;
assign n22378 =  ( n22323 ) ? ( bv_8_137_n421 ) : ( n22377 ) ;
assign n22379 =  ( n22321 ) ? ( bv_8_250_n23 ) : ( n22378 ) ;
assign n22380 =  ( n22319 ) ? ( bv_8_239_n67 ) : ( n22379 ) ;
assign n22381 =  ( n22317 ) ? ( bv_8_178_n292 ) : ( n22380 ) ;
assign n22382 =  ( n22315 ) ? ( bv_8_142_n406 ) : ( n22381 ) ;
assign n22383 =  ( n22313 ) ? ( bv_8_251_n19 ) : ( n22382 ) ;
assign n22384 =  ( n22311 ) ? ( bv_8_65_n623 ) : ( n22383 ) ;
assign n22385 =  ( n22309 ) ? ( bv_8_179_n289 ) : ( n22384 ) ;
assign n22386 =  ( n22307 ) ? ( bv_8_95_n545 ) : ( n22385 ) ;
assign n22387 =  ( n22305 ) ? ( bv_8_69_n612 ) : ( n22386 ) ;
assign n22388 =  ( n22303 ) ? ( bv_8_35_n696 ) : ( n22387 ) ;
assign n22389 =  ( n22301 ) ? ( bv_8_83_n575 ) : ( n22388 ) ;
assign n22390 =  ( n22299 ) ? ( bv_8_228_n111 ) : ( n22389 ) ;
assign n22391 =  ( n22297 ) ? ( bv_8_155_n364 ) : ( n22390 ) ;
assign n22392 =  ( n22295 ) ? ( bv_8_117_n484 ) : ( n22391 ) ;
assign n22393 =  ( n22293 ) ? ( bv_8_225_n123 ) : ( n22392 ) ;
assign n22394 =  ( n22291 ) ? ( bv_8_61_n634 ) : ( n22393 ) ;
assign n22395 =  ( n22289 ) ? ( bv_8_76_n596 ) : ( n22394 ) ;
assign n22396 =  ( n22287 ) ? ( bv_8_108_n510 ) : ( n22395 ) ;
assign n22397 =  ( n22285 ) ? ( bv_8_126_n456 ) : ( n22396 ) ;
assign n22398 =  ( n22283 ) ? ( bv_8_245_n43 ) : ( n22397 ) ;
assign n22399 =  ( n22281 ) ? ( bv_8_131_n440 ) : ( n22398 ) ;
assign n22400 =  ( n22279 ) ? ( bv_8_104_n520 ) : ( n22399 ) ;
assign n22401 =  ( n22277 ) ? ( bv_8_81_n582 ) : ( n22400 ) ;
assign n22402 =  ( n22275 ) ? ( bv_8_209_n182 ) : ( n22401 ) ;
assign n22403 =  ( n22273 ) ? ( bv_8_249_n27 ) : ( n22402 ) ;
assign n22404 =  ( n22271 ) ? ( bv_8_226_n119 ) : ( n22403 ) ;
assign n22405 =  ( n22269 ) ? ( bv_8_171_n314 ) : ( n22404 ) ;
assign n22406 =  ( n22267 ) ? ( bv_8_98_n536 ) : ( n22405 ) ;
assign n22407 =  ( n22265 ) ? ( bv_8_42_n672 ) : ( n22406 ) ;
assign n22408 =  ( n22263 ) ? ( bv_8_8_n669 ) : ( n22407 ) ;
assign n22409 =  ( n22261 ) ? ( bv_8_149_n384 ) : ( n22408 ) ;
assign n22410 =  ( n22259 ) ? ( bv_8_70_n609 ) : ( n22409 ) ;
assign n22411 =  ( n22257 ) ? ( bv_8_157_n359 ) : ( n22410 ) ;
assign n22412 =  ( n22255 ) ? ( bv_8_48_n660 ) : ( n22411 ) ;
assign n22413 =  ( n22253 ) ? ( bv_8_55_n650 ) : ( n22412 ) ;
assign n22414 =  ( n22251 ) ? ( bv_8_10_n655 ) : ( n22413 ) ;
assign n22415 =  ( n22249 ) ? ( bv_8_47_n652 ) : ( n22414 ) ;
assign n22416 =  ( n22247 ) ? ( bv_8_14_n648 ) : ( n22415 ) ;
assign n22417 =  ( n22245 ) ? ( bv_8_36_n645 ) : ( n22416 ) ;
assign n22418 =  ( n22243 ) ? ( bv_8_27_n642 ) : ( n22417 ) ;
assign n22419 =  ( n22241 ) ? ( bv_8_223_n130 ) : ( n22418 ) ;
assign n22420 =  ( n22239 ) ? ( bv_8_205_n196 ) : ( n22419 ) ;
assign n22421 =  ( n22237 ) ? ( bv_8_78_n590 ) : ( n22420 ) ;
assign n22422 =  ( n22235 ) ? ( bv_8_127_n453 ) : ( n22421 ) ;
assign n22423 =  ( n22233 ) ? ( bv_8_234_n87 ) : ( n22422 ) ;
assign n22424 =  ( n22231 ) ? ( bv_8_18_n628 ) : ( n22423 ) ;
assign n22425 =  ( n22229 ) ? ( bv_8_29_n625 ) : ( n22424 ) ;
assign n22426 =  ( n22227 ) ? ( bv_8_88_n562 ) : ( n22425 ) ;
assign n22427 =  ( n22225 ) ? ( bv_8_52_n619 ) : ( n22426 ) ;
assign n22428 =  ( n22223 ) ? ( bv_8_54_n616 ) : ( n22427 ) ;
assign n22429 =  ( n22221 ) ? ( bv_8_220_n142 ) : ( n22428 ) ;
assign n22430 =  ( n22219 ) ? ( bv_8_180_n285 ) : ( n22429 ) ;
assign n22431 =  ( n22217 ) ? ( bv_8_91_n555 ) : ( n22430 ) ;
assign n22432 =  ( n22215 ) ? ( bv_8_164_n335 ) : ( n22431 ) ;
assign n22433 =  ( n22213 ) ? ( bv_8_118_n480 ) : ( n22432 ) ;
assign n22434 =  ( n22211 ) ? ( bv_8_183_n273 ) : ( n22433 ) ;
assign n22435 =  ( n22209 ) ? ( bv_8_125_n459 ) : ( n22434 ) ;
assign n22436 =  ( n22207 ) ? ( bv_8_82_n578 ) : ( n22435 ) ;
assign n22437 =  ( n22205 ) ? ( bv_8_221_n138 ) : ( n22436 ) ;
assign n22438 =  ( n22203 ) ? ( bv_8_94_n548 ) : ( n22437 ) ;
assign n22439 =  ( n22201 ) ? ( bv_8_19_n588 ) : ( n22438 ) ;
assign n22440 =  ( n22199 ) ? ( bv_8_166_n328 ) : ( n22439 ) ;
assign n22441 =  ( n22197 ) ? ( bv_8_185_n266 ) : ( n22440 ) ;
assign n22442 =  ( n22195 ) ? ( bv_8_0_n580 ) : ( n22441 ) ;
assign n22443 =  ( n22193 ) ? ( bv_8_193_n239 ) : ( n22442 ) ;
assign n22444 =  ( n22191 ) ? ( bv_8_64_n573 ) : ( n22443 ) ;
assign n22445 =  ( n22189 ) ? ( bv_8_227_n115 ) : ( n22444 ) ;
assign n22446 =  ( n22187 ) ? ( bv_8_121_n470 ) : ( n22445 ) ;
assign n22447 =  ( n22185 ) ? ( bv_8_182_n277 ) : ( n22446 ) ;
assign n22448 =  ( n22183 ) ? ( bv_8_212_n171 ) : ( n22447 ) ;
assign n22449 =  ( n22181 ) ? ( bv_8_141_n410 ) : ( n22448 ) ;
assign n22450 =  ( n22179 ) ? ( bv_8_103_n523 ) : ( n22449 ) ;
assign n22451 =  ( n22177 ) ? ( bv_8_114_n494 ) : ( n22450 ) ;
assign n22452 =  ( n22175 ) ? ( bv_8_148_n388 ) : ( n22451 ) ;
assign n22453 =  ( n22173 ) ? ( bv_8_152_n374 ) : ( n22452 ) ;
assign n22454 =  ( n22171 ) ? ( bv_8_176_n299 ) : ( n22453 ) ;
assign n22455 =  ( n22169 ) ? ( bv_8_133_n434 ) : ( n22454 ) ;
assign n22456 =  ( n22167 ) ? ( bv_8_187_n260 ) : ( n22455 ) ;
assign n22457 =  ( n22165 ) ? ( bv_8_197_n224 ) : ( n22456 ) ;
assign n22458 =  ( n22163 ) ? ( bv_8_79_n538 ) : ( n22457 ) ;
assign n22459 =  ( n22161 ) ? ( bv_8_237_n75 ) : ( n22458 ) ;
assign n22460 =  ( n22159 ) ? ( bv_8_134_n431 ) : ( n22459 ) ;
assign n22461 =  ( n22157 ) ? ( bv_8_154_n368 ) : ( n22460 ) ;
assign n22462 =  ( n22155 ) ? ( bv_8_102_n527 ) : ( n22461 ) ;
assign n22463 =  ( n22153 ) ? ( bv_8_17_n525 ) : ( n22462 ) ;
assign n22464 =  ( n22151 ) ? ( bv_8_138_n418 ) : ( n22463 ) ;
assign n22465 =  ( n22149 ) ? ( bv_8_233_n91 ) : ( n22464 ) ;
assign n22466 =  ( n22147 ) ? ( bv_8_4_n516 ) : ( n22465 ) ;
assign n22467 =  ( n22145 ) ? ( bv_8_254_n7 ) : ( n22466 ) ;
assign n22468 =  ( n22143 ) ? ( bv_8_160_n350 ) : ( n22467 ) ;
assign n22469 =  ( n22141 ) ? ( bv_8_120_n474 ) : ( n22468 ) ;
assign n22470 =  ( n22139 ) ? ( bv_8_37_n506 ) : ( n22469 ) ;
assign n22471 =  ( n22137 ) ? ( bv_8_75_n503 ) : ( n22470 ) ;
assign n22472 =  ( n22135 ) ? ( bv_8_162_n343 ) : ( n22471 ) ;
assign n22473 =  ( n22133 ) ? ( bv_8_93_n498 ) : ( n22472 ) ;
assign n22474 =  ( n22131 ) ? ( bv_8_128_n450 ) : ( n22473 ) ;
assign n22475 =  ( n22129 ) ? ( bv_8_5_n492 ) : ( n22474 ) ;
assign n22476 =  ( n22127 ) ? ( bv_8_63_n489 ) : ( n22475 ) ;
assign n22477 =  ( n22125 ) ? ( bv_8_33_n486 ) : ( n22476 ) ;
assign n22478 =  ( n22123 ) ? ( bv_8_112_n482 ) : ( n22477 ) ;
assign n22479 =  ( n22121 ) ? ( bv_8_241_n59 ) : ( n22478 ) ;
assign n22480 =  ( n22119 ) ? ( bv_8_99_n476 ) : ( n22479 ) ;
assign n22481 =  ( n22117 ) ? ( bv_8_119_n472 ) : ( n22480 ) ;
assign n22482 =  ( n22115 ) ? ( bv_8_175_n302 ) : ( n22481 ) ;
assign n22483 =  ( n22113 ) ? ( bv_8_66_n466 ) : ( n22482 ) ;
assign n22484 =  ( n22111 ) ? ( bv_8_32_n463 ) : ( n22483 ) ;
assign n22485 =  ( n22109 ) ? ( bv_8_229_n107 ) : ( n22484 ) ;
assign n22486 =  ( n22107 ) ? ( bv_8_253_n11 ) : ( n22485 ) ;
assign n22487 =  ( n22105 ) ? ( bv_8_191_n246 ) : ( n22486 ) ;
assign n22488 =  ( n22103 ) ? ( bv_8_129_n446 ) : ( n22487 ) ;
assign n22489 =  ( n22101 ) ? ( bv_8_24_n448 ) : ( n22488 ) ;
assign n22490 =  ( n22099 ) ? ( bv_8_38_n444 ) : ( n22489 ) ;
assign n22491 =  ( n22097 ) ? ( bv_8_195_n232 ) : ( n22490 ) ;
assign n22492 =  ( n22095 ) ? ( bv_8_190_n250 ) : ( n22491 ) ;
assign n22493 =  ( n22093 ) ? ( bv_8_53_n436 ) : ( n22492 ) ;
assign n22494 =  ( n22091 ) ? ( bv_8_136_n425 ) : ( n22493 ) ;
assign n22495 =  ( n22089 ) ? ( bv_8_46_n429 ) : ( n22494 ) ;
assign n22496 =  ( n22087 ) ? ( bv_8_147_n392 ) : ( n22495 ) ;
assign n22497 =  ( n22085 ) ? ( bv_8_85_n423 ) : ( n22496 ) ;
assign n22498 =  ( n22083 ) ? ( bv_8_252_n15 ) : ( n22497 ) ;
assign n22499 =  ( n22081 ) ? ( bv_8_122_n416 ) : ( n22498 ) ;
assign n22500 =  ( n22079 ) ? ( bv_8_200_n213 ) : ( n22499 ) ;
assign n22501 =  ( n22077 ) ? ( bv_8_186_n263 ) : ( n22500 ) ;
assign n22502 =  ( n22075 ) ? ( bv_8_50_n408 ) : ( n22501 ) ;
assign n22503 =  ( n22073 ) ? ( bv_8_230_n103 ) : ( n22502 ) ;
assign n22504 =  ( n22071 ) ? ( bv_8_192_n242 ) : ( n22503 ) ;
assign n22505 =  ( n22069 ) ? ( bv_8_25_n399 ) : ( n22504 ) ;
assign n22506 =  ( n22067 ) ? ( bv_8_158_n355 ) : ( n22505 ) ;
assign n22507 =  ( n22065 ) ? ( bv_8_163_n339 ) : ( n22506 ) ;
assign n22508 =  ( n22063 ) ? ( bv_8_68_n390 ) : ( n22507 ) ;
assign n22509 =  ( n22061 ) ? ( bv_8_84_n386 ) : ( n22508 ) ;
assign n22510 =  ( n22059 ) ? ( bv_8_59_n382 ) : ( n22509 ) ;
assign n22511 =  ( n22057 ) ? ( bv_8_11_n379 ) : ( n22510 ) ;
assign n22512 =  ( n22055 ) ? ( bv_8_140_n376 ) : ( n22511 ) ;
assign n22513 =  ( n22053 ) ? ( bv_8_199_n216 ) : ( n22512 ) ;
assign n22514 =  ( n22051 ) ? ( bv_8_107_n370 ) : ( n22513 ) ;
assign n22515 =  ( n22049 ) ? ( bv_8_40_n366 ) : ( n22514 ) ;
assign n22516 =  ( n22047 ) ? ( bv_8_167_n325 ) : ( n22515 ) ;
assign n22517 =  ( n22045 ) ? ( bv_8_188_n257 ) : ( n22516 ) ;
assign n22518 =  ( n22043 ) ? ( bv_8_22_n357 ) : ( n22517 ) ;
assign n22519 =  ( n22041 ) ? ( bv_8_173_n307 ) : ( n22518 ) ;
assign n22520 =  ( n22039 ) ? ( bv_8_219_n146 ) : ( n22519 ) ;
assign n22521 =  ( n22037 ) ? ( bv_8_100_n348 ) : ( n22520 ) ;
assign n22522 =  ( n22035 ) ? ( bv_8_116_n345 ) : ( n22521 ) ;
assign n22523 =  ( n22033 ) ? ( bv_8_20_n341 ) : ( n22522 ) ;
assign n22524 =  ( n22031 ) ? ( bv_8_146_n337 ) : ( n22523 ) ;
assign n22525 =  ( n22029 ) ? ( bv_8_12_n333 ) : ( n22524 ) ;
assign n22526 =  ( n22027 ) ? ( bv_8_72_n330 ) : ( n22525 ) ;
assign n22527 =  ( n22025 ) ? ( bv_8_184_n270 ) : ( n22526 ) ;
assign n22528 =  ( n22023 ) ? ( bv_8_159_n323 ) : ( n22527 ) ;
assign n22529 =  ( n22021 ) ? ( bv_8_189_n254 ) : ( n22528 ) ;
assign n22530 =  ( n22019 ) ? ( bv_8_67_n318 ) : ( n22529 ) ;
assign n22531 =  ( n22017 ) ? ( bv_8_196_n228 ) : ( n22530 ) ;
assign n22532 =  ( n22015 ) ? ( bv_8_57_n312 ) : ( n22531 ) ;
assign n22533 =  ( n22013 ) ? ( bv_8_49_n309 ) : ( n22532 ) ;
assign n22534 =  ( n22011 ) ? ( bv_8_211_n175 ) : ( n22533 ) ;
assign n22535 =  ( n22009 ) ? ( bv_8_242_n55 ) : ( n22534 ) ;
assign n22536 =  ( n22007 ) ? ( bv_8_213_n167 ) : ( n22535 ) ;
assign n22537 =  ( n22005 ) ? ( bv_8_139_n297 ) : ( n22536 ) ;
assign n22538 =  ( n22003 ) ? ( bv_8_110_n294 ) : ( n22537 ) ;
assign n22539 =  ( n22001 ) ? ( bv_8_218_n150 ) : ( n22538 ) ;
assign n22540 =  ( n21999 ) ? ( bv_8_1_n287 ) : ( n22539 ) ;
assign n22541 =  ( n21997 ) ? ( bv_8_177_n283 ) : ( n22540 ) ;
assign n22542 =  ( n21995 ) ? ( bv_8_156_n279 ) : ( n22541 ) ;
assign n22543 =  ( n21993 ) ? ( bv_8_73_n275 ) : ( n22542 ) ;
assign n22544 =  ( n21991 ) ? ( bv_8_216_n157 ) : ( n22543 ) ;
assign n22545 =  ( n21989 ) ? ( bv_8_172_n268 ) : ( n22544 ) ;
assign n22546 =  ( n21987 ) ? ( bv_8_243_n51 ) : ( n22545 ) ;
assign n22547 =  ( n21985 ) ? ( bv_8_207_n188 ) : ( n22546 ) ;
assign n22548 =  ( n21983 ) ? ( bv_8_202_n207 ) : ( n22547 ) ;
assign n22549 =  ( n21981 ) ? ( bv_8_244_n47 ) : ( n22548 ) ;
assign n22550 =  ( n21979 ) ? ( bv_8_71_n252 ) : ( n22549 ) ;
assign n22551 =  ( n21977 ) ? ( bv_8_16_n248 ) : ( n22550 ) ;
assign n22552 =  ( n21975 ) ? ( bv_8_111_n244 ) : ( n22551 ) ;
assign n22553 =  ( n21973 ) ? ( bv_8_240_n63 ) : ( n22552 ) ;
assign n22554 =  ( n21971 ) ? ( bv_8_74_n237 ) : ( n22553 ) ;
assign n22555 =  ( n21969 ) ? ( bv_8_92_n234 ) : ( n22554 ) ;
assign n22556 =  ( n21967 ) ? ( bv_8_56_n230 ) : ( n22555 ) ;
assign n22557 =  ( n21965 ) ? ( bv_8_87_n226 ) : ( n22556 ) ;
assign n22558 =  ( n21963 ) ? ( bv_8_115_n222 ) : ( n22557 ) ;
assign n22559 =  ( n21961 ) ? ( bv_8_151_n218 ) : ( n22558 ) ;
assign n22560 =  ( n21959 ) ? ( bv_8_203_n203 ) : ( n22559 ) ;
assign n22561 =  ( n21957 ) ? ( bv_8_161_n211 ) : ( n22560 ) ;
assign n22562 =  ( n21955 ) ? ( bv_8_232_n95 ) : ( n22561 ) ;
assign n22563 =  ( n21953 ) ? ( bv_8_62_n205 ) : ( n22562 ) ;
assign n22564 =  ( n21951 ) ? ( bv_8_150_n201 ) : ( n22563 ) ;
assign n22565 =  ( n21949 ) ? ( bv_8_97_n198 ) : ( n22564 ) ;
assign n22566 =  ( n21947 ) ? ( bv_8_13_n194 ) : ( n22565 ) ;
assign n22567 =  ( n21945 ) ? ( bv_8_15_n190 ) : ( n22566 ) ;
assign n22568 =  ( n21943 ) ? ( bv_8_224_n126 ) : ( n22567 ) ;
assign n22569 =  ( n21941 ) ? ( bv_8_124_n184 ) : ( n22568 ) ;
assign n22570 =  ( n21939 ) ? ( bv_8_113_n180 ) : ( n22569 ) ;
assign n22571 =  ( n21937 ) ? ( bv_8_204_n177 ) : ( n22570 ) ;
assign n22572 =  ( n21935 ) ? ( bv_8_144_n173 ) : ( n22571 ) ;
assign n22573 =  ( n21933 ) ? ( bv_8_6_n169 ) : ( n22572 ) ;
assign n22574 =  ( n21931 ) ? ( bv_8_247_n35 ) : ( n22573 ) ;
assign n22575 =  ( n21929 ) ? ( bv_8_28_n162 ) : ( n22574 ) ;
assign n22576 =  ( n21927 ) ? ( bv_8_194_n159 ) : ( n22575 ) ;
assign n22577 =  ( n21925 ) ? ( bv_8_106_n155 ) : ( n22576 ) ;
assign n22578 =  ( n21923 ) ? ( bv_8_174_n152 ) : ( n22577 ) ;
assign n22579 =  ( n21921 ) ? ( bv_8_105_n148 ) : ( n22578 ) ;
assign n22580 =  ( n21919 ) ? ( bv_8_23_n144 ) : ( n22579 ) ;
assign n22581 =  ( n21917 ) ? ( bv_8_153_n140 ) : ( n22580 ) ;
assign n22582 =  ( n21915 ) ? ( bv_8_58_n136 ) : ( n22581 ) ;
assign n22583 =  ( n21913 ) ? ( bv_8_39_n132 ) : ( n22582 ) ;
assign n22584 =  ( n21911 ) ? ( bv_8_217_n128 ) : ( n22583 ) ;
assign n22585 =  ( n21909 ) ? ( bv_8_235_n83 ) : ( n22584 ) ;
assign n22586 =  ( n21907 ) ? ( bv_8_43_n121 ) : ( n22585 ) ;
assign n22587 =  ( n21905 ) ? ( bv_8_34_n117 ) : ( n22586 ) ;
assign n22588 =  ( n21903 ) ? ( bv_8_210_n113 ) : ( n22587 ) ;
assign n22589 =  ( n21901 ) ? ( bv_8_169_n109 ) : ( n22588 ) ;
assign n22590 =  ( n21899 ) ? ( bv_8_7_n105 ) : ( n22589 ) ;
assign n22591 =  ( n21897 ) ? ( bv_8_51_n101 ) : ( n22590 ) ;
assign n22592 =  ( n21895 ) ? ( bv_8_45_n97 ) : ( n22591 ) ;
assign n22593 =  ( n21893 ) ? ( bv_8_60_n93 ) : ( n22592 ) ;
assign n22594 =  ( n21891 ) ? ( bv_8_21_n89 ) : ( n22593 ) ;
assign n22595 =  ( n21889 ) ? ( bv_8_201_n85 ) : ( n22594 ) ;
assign n22596 =  ( n21887 ) ? ( bv_8_135_n81 ) : ( n22595 ) ;
assign n22597 =  ( n21885 ) ? ( bv_8_170_n77 ) : ( n22596 ) ;
assign n22598 =  ( n21883 ) ? ( bv_8_80_n73 ) : ( n22597 ) ;
assign n22599 =  ( n21881 ) ? ( bv_8_165_n69 ) : ( n22598 ) ;
assign n22600 =  ( n21879 ) ? ( bv_8_3_n65 ) : ( n22599 ) ;
assign n22601 =  ( n21877 ) ? ( bv_8_89_n61 ) : ( n22600 ) ;
assign n22602 =  ( n21875 ) ? ( bv_8_9_n57 ) : ( n22601 ) ;
assign n22603 =  ( n21873 ) ? ( bv_8_26_n53 ) : ( n22602 ) ;
assign n22604 =  ( n21871 ) ? ( bv_8_101_n49 ) : ( n22603 ) ;
assign n22605 =  ( n21869 ) ? ( bv_8_215_n45 ) : ( n22604 ) ;
assign n22606 =  ( n21867 ) ? ( bv_8_132_n41 ) : ( n22605 ) ;
assign n22607 =  ( n21865 ) ? ( bv_8_208_n37 ) : ( n22606 ) ;
assign n22608 =  ( n21863 ) ? ( bv_8_130_n33 ) : ( n22607 ) ;
assign n22609 =  ( n21861 ) ? ( bv_8_41_n29 ) : ( n22608 ) ;
assign n22610 =  ( n21859 ) ? ( bv_8_90_n25 ) : ( n22609 ) ;
assign n22611 =  ( n21857 ) ? ( bv_8_30_n21 ) : ( n22610 ) ;
assign n22612 =  ( n21855 ) ? ( bv_8_123_n17 ) : ( n22611 ) ;
assign n22613 =  ( n21853 ) ? ( bv_8_168_n13 ) : ( n22612 ) ;
assign n22614 =  ( n21851 ) ? ( bv_8_109_n9 ) : ( n22613 ) ;
assign n22615 =  ( n21849 ) ? ( bv_8_44_n5 ) : ( n22614 ) ;
assign n22616 =  ( n21847 ) ^ ( n22615 )  ;
assign n22617 = key[31:24] ;
assign n22618 =  ( n22616 ) ^ ( n22617 )  ;
assign n22619 =  { ( n18772 ) , ( n22618 ) }  ;
assign n22620 =  ( n20308 ) ^ ( n21077 )  ;
assign n22621 = state_in[79:72] ;
assign n22622 =  ( n22621 ) == ( bv_8_255_n3 )  ;
assign n22623 = state_in[79:72] ;
assign n22624 =  ( n22623 ) == ( bv_8_254_n7 )  ;
assign n22625 = state_in[79:72] ;
assign n22626 =  ( n22625 ) == ( bv_8_253_n11 )  ;
assign n22627 = state_in[79:72] ;
assign n22628 =  ( n22627 ) == ( bv_8_252_n15 )  ;
assign n22629 = state_in[79:72] ;
assign n22630 =  ( n22629 ) == ( bv_8_251_n19 )  ;
assign n22631 = state_in[79:72] ;
assign n22632 =  ( n22631 ) == ( bv_8_250_n23 )  ;
assign n22633 = state_in[79:72] ;
assign n22634 =  ( n22633 ) == ( bv_8_249_n27 )  ;
assign n22635 = state_in[79:72] ;
assign n22636 =  ( n22635 ) == ( bv_8_248_n31 )  ;
assign n22637 = state_in[79:72] ;
assign n22638 =  ( n22637 ) == ( bv_8_247_n35 )  ;
assign n22639 = state_in[79:72] ;
assign n22640 =  ( n22639 ) == ( bv_8_246_n39 )  ;
assign n22641 = state_in[79:72] ;
assign n22642 =  ( n22641 ) == ( bv_8_245_n43 )  ;
assign n22643 = state_in[79:72] ;
assign n22644 =  ( n22643 ) == ( bv_8_244_n47 )  ;
assign n22645 = state_in[79:72] ;
assign n22646 =  ( n22645 ) == ( bv_8_243_n51 )  ;
assign n22647 = state_in[79:72] ;
assign n22648 =  ( n22647 ) == ( bv_8_242_n55 )  ;
assign n22649 = state_in[79:72] ;
assign n22650 =  ( n22649 ) == ( bv_8_241_n59 )  ;
assign n22651 = state_in[79:72] ;
assign n22652 =  ( n22651 ) == ( bv_8_240_n63 )  ;
assign n22653 = state_in[79:72] ;
assign n22654 =  ( n22653 ) == ( bv_8_239_n67 )  ;
assign n22655 = state_in[79:72] ;
assign n22656 =  ( n22655 ) == ( bv_8_238_n71 )  ;
assign n22657 = state_in[79:72] ;
assign n22658 =  ( n22657 ) == ( bv_8_237_n75 )  ;
assign n22659 = state_in[79:72] ;
assign n22660 =  ( n22659 ) == ( bv_8_236_n79 )  ;
assign n22661 = state_in[79:72] ;
assign n22662 =  ( n22661 ) == ( bv_8_235_n83 )  ;
assign n22663 = state_in[79:72] ;
assign n22664 =  ( n22663 ) == ( bv_8_234_n87 )  ;
assign n22665 = state_in[79:72] ;
assign n22666 =  ( n22665 ) == ( bv_8_233_n91 )  ;
assign n22667 = state_in[79:72] ;
assign n22668 =  ( n22667 ) == ( bv_8_232_n95 )  ;
assign n22669 = state_in[79:72] ;
assign n22670 =  ( n22669 ) == ( bv_8_231_n99 )  ;
assign n22671 = state_in[79:72] ;
assign n22672 =  ( n22671 ) == ( bv_8_230_n103 )  ;
assign n22673 = state_in[79:72] ;
assign n22674 =  ( n22673 ) == ( bv_8_229_n107 )  ;
assign n22675 = state_in[79:72] ;
assign n22676 =  ( n22675 ) == ( bv_8_228_n111 )  ;
assign n22677 = state_in[79:72] ;
assign n22678 =  ( n22677 ) == ( bv_8_227_n115 )  ;
assign n22679 = state_in[79:72] ;
assign n22680 =  ( n22679 ) == ( bv_8_226_n119 )  ;
assign n22681 = state_in[79:72] ;
assign n22682 =  ( n22681 ) == ( bv_8_225_n123 )  ;
assign n22683 = state_in[79:72] ;
assign n22684 =  ( n22683 ) == ( bv_8_224_n126 )  ;
assign n22685 = state_in[79:72] ;
assign n22686 =  ( n22685 ) == ( bv_8_223_n130 )  ;
assign n22687 = state_in[79:72] ;
assign n22688 =  ( n22687 ) == ( bv_8_222_n134 )  ;
assign n22689 = state_in[79:72] ;
assign n22690 =  ( n22689 ) == ( bv_8_221_n138 )  ;
assign n22691 = state_in[79:72] ;
assign n22692 =  ( n22691 ) == ( bv_8_220_n142 )  ;
assign n22693 = state_in[79:72] ;
assign n22694 =  ( n22693 ) == ( bv_8_219_n146 )  ;
assign n22695 = state_in[79:72] ;
assign n22696 =  ( n22695 ) == ( bv_8_218_n150 )  ;
assign n22697 = state_in[79:72] ;
assign n22698 =  ( n22697 ) == ( bv_8_217_n128 )  ;
assign n22699 = state_in[79:72] ;
assign n22700 =  ( n22699 ) == ( bv_8_216_n157 )  ;
assign n22701 = state_in[79:72] ;
assign n22702 =  ( n22701 ) == ( bv_8_215_n45 )  ;
assign n22703 = state_in[79:72] ;
assign n22704 =  ( n22703 ) == ( bv_8_214_n164 )  ;
assign n22705 = state_in[79:72] ;
assign n22706 =  ( n22705 ) == ( bv_8_213_n167 )  ;
assign n22707 = state_in[79:72] ;
assign n22708 =  ( n22707 ) == ( bv_8_212_n171 )  ;
assign n22709 = state_in[79:72] ;
assign n22710 =  ( n22709 ) == ( bv_8_211_n175 )  ;
assign n22711 = state_in[79:72] ;
assign n22712 =  ( n22711 ) == ( bv_8_210_n113 )  ;
assign n22713 = state_in[79:72] ;
assign n22714 =  ( n22713 ) == ( bv_8_209_n182 )  ;
assign n22715 = state_in[79:72] ;
assign n22716 =  ( n22715 ) == ( bv_8_208_n37 )  ;
assign n22717 = state_in[79:72] ;
assign n22718 =  ( n22717 ) == ( bv_8_207_n188 )  ;
assign n22719 = state_in[79:72] ;
assign n22720 =  ( n22719 ) == ( bv_8_206_n192 )  ;
assign n22721 = state_in[79:72] ;
assign n22722 =  ( n22721 ) == ( bv_8_205_n196 )  ;
assign n22723 = state_in[79:72] ;
assign n22724 =  ( n22723 ) == ( bv_8_204_n177 )  ;
assign n22725 = state_in[79:72] ;
assign n22726 =  ( n22725 ) == ( bv_8_203_n203 )  ;
assign n22727 = state_in[79:72] ;
assign n22728 =  ( n22727 ) == ( bv_8_202_n207 )  ;
assign n22729 = state_in[79:72] ;
assign n22730 =  ( n22729 ) == ( bv_8_201_n85 )  ;
assign n22731 = state_in[79:72] ;
assign n22732 =  ( n22731 ) == ( bv_8_200_n213 )  ;
assign n22733 = state_in[79:72] ;
assign n22734 =  ( n22733 ) == ( bv_8_199_n216 )  ;
assign n22735 = state_in[79:72] ;
assign n22736 =  ( n22735 ) == ( bv_8_198_n220 )  ;
assign n22737 = state_in[79:72] ;
assign n22738 =  ( n22737 ) == ( bv_8_197_n224 )  ;
assign n22739 = state_in[79:72] ;
assign n22740 =  ( n22739 ) == ( bv_8_196_n228 )  ;
assign n22741 = state_in[79:72] ;
assign n22742 =  ( n22741 ) == ( bv_8_195_n232 )  ;
assign n22743 = state_in[79:72] ;
assign n22744 =  ( n22743 ) == ( bv_8_194_n159 )  ;
assign n22745 = state_in[79:72] ;
assign n22746 =  ( n22745 ) == ( bv_8_193_n239 )  ;
assign n22747 = state_in[79:72] ;
assign n22748 =  ( n22747 ) == ( bv_8_192_n242 )  ;
assign n22749 = state_in[79:72] ;
assign n22750 =  ( n22749 ) == ( bv_8_191_n246 )  ;
assign n22751 = state_in[79:72] ;
assign n22752 =  ( n22751 ) == ( bv_8_190_n250 )  ;
assign n22753 = state_in[79:72] ;
assign n22754 =  ( n22753 ) == ( bv_8_189_n254 )  ;
assign n22755 = state_in[79:72] ;
assign n22756 =  ( n22755 ) == ( bv_8_188_n257 )  ;
assign n22757 = state_in[79:72] ;
assign n22758 =  ( n22757 ) == ( bv_8_187_n260 )  ;
assign n22759 = state_in[79:72] ;
assign n22760 =  ( n22759 ) == ( bv_8_186_n263 )  ;
assign n22761 = state_in[79:72] ;
assign n22762 =  ( n22761 ) == ( bv_8_185_n266 )  ;
assign n22763 = state_in[79:72] ;
assign n22764 =  ( n22763 ) == ( bv_8_184_n270 )  ;
assign n22765 = state_in[79:72] ;
assign n22766 =  ( n22765 ) == ( bv_8_183_n273 )  ;
assign n22767 = state_in[79:72] ;
assign n22768 =  ( n22767 ) == ( bv_8_182_n277 )  ;
assign n22769 = state_in[79:72] ;
assign n22770 =  ( n22769 ) == ( bv_8_181_n281 )  ;
assign n22771 = state_in[79:72] ;
assign n22772 =  ( n22771 ) == ( bv_8_180_n285 )  ;
assign n22773 = state_in[79:72] ;
assign n22774 =  ( n22773 ) == ( bv_8_179_n289 )  ;
assign n22775 = state_in[79:72] ;
assign n22776 =  ( n22775 ) == ( bv_8_178_n292 )  ;
assign n22777 = state_in[79:72] ;
assign n22778 =  ( n22777 ) == ( bv_8_177_n283 )  ;
assign n22779 = state_in[79:72] ;
assign n22780 =  ( n22779 ) == ( bv_8_176_n299 )  ;
assign n22781 = state_in[79:72] ;
assign n22782 =  ( n22781 ) == ( bv_8_175_n302 )  ;
assign n22783 = state_in[79:72] ;
assign n22784 =  ( n22783 ) == ( bv_8_174_n152 )  ;
assign n22785 = state_in[79:72] ;
assign n22786 =  ( n22785 ) == ( bv_8_173_n307 )  ;
assign n22787 = state_in[79:72] ;
assign n22788 =  ( n22787 ) == ( bv_8_172_n268 )  ;
assign n22789 = state_in[79:72] ;
assign n22790 =  ( n22789 ) == ( bv_8_171_n314 )  ;
assign n22791 = state_in[79:72] ;
assign n22792 =  ( n22791 ) == ( bv_8_170_n77 )  ;
assign n22793 = state_in[79:72] ;
assign n22794 =  ( n22793 ) == ( bv_8_169_n109 )  ;
assign n22795 = state_in[79:72] ;
assign n22796 =  ( n22795 ) == ( bv_8_168_n13 )  ;
assign n22797 = state_in[79:72] ;
assign n22798 =  ( n22797 ) == ( bv_8_167_n325 )  ;
assign n22799 = state_in[79:72] ;
assign n22800 =  ( n22799 ) == ( bv_8_166_n328 )  ;
assign n22801 = state_in[79:72] ;
assign n22802 =  ( n22801 ) == ( bv_8_165_n69 )  ;
assign n22803 = state_in[79:72] ;
assign n22804 =  ( n22803 ) == ( bv_8_164_n335 )  ;
assign n22805 = state_in[79:72] ;
assign n22806 =  ( n22805 ) == ( bv_8_163_n339 )  ;
assign n22807 = state_in[79:72] ;
assign n22808 =  ( n22807 ) == ( bv_8_162_n343 )  ;
assign n22809 = state_in[79:72] ;
assign n22810 =  ( n22809 ) == ( bv_8_161_n211 )  ;
assign n22811 = state_in[79:72] ;
assign n22812 =  ( n22811 ) == ( bv_8_160_n350 )  ;
assign n22813 = state_in[79:72] ;
assign n22814 =  ( n22813 ) == ( bv_8_159_n323 )  ;
assign n22815 = state_in[79:72] ;
assign n22816 =  ( n22815 ) == ( bv_8_158_n355 )  ;
assign n22817 = state_in[79:72] ;
assign n22818 =  ( n22817 ) == ( bv_8_157_n359 )  ;
assign n22819 = state_in[79:72] ;
assign n22820 =  ( n22819 ) == ( bv_8_156_n279 )  ;
assign n22821 = state_in[79:72] ;
assign n22822 =  ( n22821 ) == ( bv_8_155_n364 )  ;
assign n22823 = state_in[79:72] ;
assign n22824 =  ( n22823 ) == ( bv_8_154_n368 )  ;
assign n22825 = state_in[79:72] ;
assign n22826 =  ( n22825 ) == ( bv_8_153_n140 )  ;
assign n22827 = state_in[79:72] ;
assign n22828 =  ( n22827 ) == ( bv_8_152_n374 )  ;
assign n22829 = state_in[79:72] ;
assign n22830 =  ( n22829 ) == ( bv_8_151_n218 )  ;
assign n22831 = state_in[79:72] ;
assign n22832 =  ( n22831 ) == ( bv_8_150_n201 )  ;
assign n22833 = state_in[79:72] ;
assign n22834 =  ( n22833 ) == ( bv_8_149_n384 )  ;
assign n22835 = state_in[79:72] ;
assign n22836 =  ( n22835 ) == ( bv_8_148_n388 )  ;
assign n22837 = state_in[79:72] ;
assign n22838 =  ( n22837 ) == ( bv_8_147_n392 )  ;
assign n22839 = state_in[79:72] ;
assign n22840 =  ( n22839 ) == ( bv_8_146_n337 )  ;
assign n22841 = state_in[79:72] ;
assign n22842 =  ( n22841 ) == ( bv_8_145_n397 )  ;
assign n22843 = state_in[79:72] ;
assign n22844 =  ( n22843 ) == ( bv_8_144_n173 )  ;
assign n22845 = state_in[79:72] ;
assign n22846 =  ( n22845 ) == ( bv_8_143_n403 )  ;
assign n22847 = state_in[79:72] ;
assign n22848 =  ( n22847 ) == ( bv_8_142_n406 )  ;
assign n22849 = state_in[79:72] ;
assign n22850 =  ( n22849 ) == ( bv_8_141_n410 )  ;
assign n22851 = state_in[79:72] ;
assign n22852 =  ( n22851 ) == ( bv_8_140_n376 )  ;
assign n22853 = state_in[79:72] ;
assign n22854 =  ( n22853 ) == ( bv_8_139_n297 )  ;
assign n22855 = state_in[79:72] ;
assign n22856 =  ( n22855 ) == ( bv_8_138_n418 )  ;
assign n22857 = state_in[79:72] ;
assign n22858 =  ( n22857 ) == ( bv_8_137_n421 )  ;
assign n22859 = state_in[79:72] ;
assign n22860 =  ( n22859 ) == ( bv_8_136_n425 )  ;
assign n22861 = state_in[79:72] ;
assign n22862 =  ( n22861 ) == ( bv_8_135_n81 )  ;
assign n22863 = state_in[79:72] ;
assign n22864 =  ( n22863 ) == ( bv_8_134_n431 )  ;
assign n22865 = state_in[79:72] ;
assign n22866 =  ( n22865 ) == ( bv_8_133_n434 )  ;
assign n22867 = state_in[79:72] ;
assign n22868 =  ( n22867 ) == ( bv_8_132_n41 )  ;
assign n22869 = state_in[79:72] ;
assign n22870 =  ( n22869 ) == ( bv_8_131_n440 )  ;
assign n22871 = state_in[79:72] ;
assign n22872 =  ( n22871 ) == ( bv_8_130_n33 )  ;
assign n22873 = state_in[79:72] ;
assign n22874 =  ( n22873 ) == ( bv_8_129_n446 )  ;
assign n22875 = state_in[79:72] ;
assign n22876 =  ( n22875 ) == ( bv_8_128_n450 )  ;
assign n22877 = state_in[79:72] ;
assign n22878 =  ( n22877 ) == ( bv_8_127_n453 )  ;
assign n22879 = state_in[79:72] ;
assign n22880 =  ( n22879 ) == ( bv_8_126_n456 )  ;
assign n22881 = state_in[79:72] ;
assign n22882 =  ( n22881 ) == ( bv_8_125_n459 )  ;
assign n22883 = state_in[79:72] ;
assign n22884 =  ( n22883 ) == ( bv_8_124_n184 )  ;
assign n22885 = state_in[79:72] ;
assign n22886 =  ( n22885 ) == ( bv_8_123_n17 )  ;
assign n22887 = state_in[79:72] ;
assign n22888 =  ( n22887 ) == ( bv_8_122_n416 )  ;
assign n22889 = state_in[79:72] ;
assign n22890 =  ( n22889 ) == ( bv_8_121_n470 )  ;
assign n22891 = state_in[79:72] ;
assign n22892 =  ( n22891 ) == ( bv_8_120_n474 )  ;
assign n22893 = state_in[79:72] ;
assign n22894 =  ( n22893 ) == ( bv_8_119_n472 )  ;
assign n22895 = state_in[79:72] ;
assign n22896 =  ( n22895 ) == ( bv_8_118_n480 )  ;
assign n22897 = state_in[79:72] ;
assign n22898 =  ( n22897 ) == ( bv_8_117_n484 )  ;
assign n22899 = state_in[79:72] ;
assign n22900 =  ( n22899 ) == ( bv_8_116_n345 )  ;
assign n22901 = state_in[79:72] ;
assign n22902 =  ( n22901 ) == ( bv_8_115_n222 )  ;
assign n22903 = state_in[79:72] ;
assign n22904 =  ( n22903 ) == ( bv_8_114_n494 )  ;
assign n22905 = state_in[79:72] ;
assign n22906 =  ( n22905 ) == ( bv_8_113_n180 )  ;
assign n22907 = state_in[79:72] ;
assign n22908 =  ( n22907 ) == ( bv_8_112_n482 )  ;
assign n22909 = state_in[79:72] ;
assign n22910 =  ( n22909 ) == ( bv_8_111_n244 )  ;
assign n22911 = state_in[79:72] ;
assign n22912 =  ( n22911 ) == ( bv_8_110_n294 )  ;
assign n22913 = state_in[79:72] ;
assign n22914 =  ( n22913 ) == ( bv_8_109_n9 )  ;
assign n22915 = state_in[79:72] ;
assign n22916 =  ( n22915 ) == ( bv_8_108_n510 )  ;
assign n22917 = state_in[79:72] ;
assign n22918 =  ( n22917 ) == ( bv_8_107_n370 )  ;
assign n22919 = state_in[79:72] ;
assign n22920 =  ( n22919 ) == ( bv_8_106_n155 )  ;
assign n22921 = state_in[79:72] ;
assign n22922 =  ( n22921 ) == ( bv_8_105_n148 )  ;
assign n22923 = state_in[79:72] ;
assign n22924 =  ( n22923 ) == ( bv_8_104_n520 )  ;
assign n22925 = state_in[79:72] ;
assign n22926 =  ( n22925 ) == ( bv_8_103_n523 )  ;
assign n22927 = state_in[79:72] ;
assign n22928 =  ( n22927 ) == ( bv_8_102_n527 )  ;
assign n22929 = state_in[79:72] ;
assign n22930 =  ( n22929 ) == ( bv_8_101_n49 )  ;
assign n22931 = state_in[79:72] ;
assign n22932 =  ( n22931 ) == ( bv_8_100_n348 )  ;
assign n22933 = state_in[79:72] ;
assign n22934 =  ( n22933 ) == ( bv_8_99_n476 )  ;
assign n22935 = state_in[79:72] ;
assign n22936 =  ( n22935 ) == ( bv_8_98_n536 )  ;
assign n22937 = state_in[79:72] ;
assign n22938 =  ( n22937 ) == ( bv_8_97_n198 )  ;
assign n22939 = state_in[79:72] ;
assign n22940 =  ( n22939 ) == ( bv_8_96_n542 )  ;
assign n22941 = state_in[79:72] ;
assign n22942 =  ( n22941 ) == ( bv_8_95_n545 )  ;
assign n22943 = state_in[79:72] ;
assign n22944 =  ( n22943 ) == ( bv_8_94_n548 )  ;
assign n22945 = state_in[79:72] ;
assign n22946 =  ( n22945 ) == ( bv_8_93_n498 )  ;
assign n22947 = state_in[79:72] ;
assign n22948 =  ( n22947 ) == ( bv_8_92_n234 )  ;
assign n22949 = state_in[79:72] ;
assign n22950 =  ( n22949 ) == ( bv_8_91_n555 )  ;
assign n22951 = state_in[79:72] ;
assign n22952 =  ( n22951 ) == ( bv_8_90_n25 )  ;
assign n22953 = state_in[79:72] ;
assign n22954 =  ( n22953 ) == ( bv_8_89_n61 )  ;
assign n22955 = state_in[79:72] ;
assign n22956 =  ( n22955 ) == ( bv_8_88_n562 )  ;
assign n22957 = state_in[79:72] ;
assign n22958 =  ( n22957 ) == ( bv_8_87_n226 )  ;
assign n22959 = state_in[79:72] ;
assign n22960 =  ( n22959 ) == ( bv_8_86_n567 )  ;
assign n22961 = state_in[79:72] ;
assign n22962 =  ( n22961 ) == ( bv_8_85_n423 )  ;
assign n22963 = state_in[79:72] ;
assign n22964 =  ( n22963 ) == ( bv_8_84_n386 )  ;
assign n22965 = state_in[79:72] ;
assign n22966 =  ( n22965 ) == ( bv_8_83_n575 )  ;
assign n22967 = state_in[79:72] ;
assign n22968 =  ( n22967 ) == ( bv_8_82_n578 )  ;
assign n22969 = state_in[79:72] ;
assign n22970 =  ( n22969 ) == ( bv_8_81_n582 )  ;
assign n22971 = state_in[79:72] ;
assign n22972 =  ( n22971 ) == ( bv_8_80_n73 )  ;
assign n22973 = state_in[79:72] ;
assign n22974 =  ( n22973 ) == ( bv_8_79_n538 )  ;
assign n22975 = state_in[79:72] ;
assign n22976 =  ( n22975 ) == ( bv_8_78_n590 )  ;
assign n22977 = state_in[79:72] ;
assign n22978 =  ( n22977 ) == ( bv_8_77_n593 )  ;
assign n22979 = state_in[79:72] ;
assign n22980 =  ( n22979 ) == ( bv_8_76_n596 )  ;
assign n22981 = state_in[79:72] ;
assign n22982 =  ( n22981 ) == ( bv_8_75_n503 )  ;
assign n22983 = state_in[79:72] ;
assign n22984 =  ( n22983 ) == ( bv_8_74_n237 )  ;
assign n22985 = state_in[79:72] ;
assign n22986 =  ( n22985 ) == ( bv_8_73_n275 )  ;
assign n22987 = state_in[79:72] ;
assign n22988 =  ( n22987 ) == ( bv_8_72_n330 )  ;
assign n22989 = state_in[79:72] ;
assign n22990 =  ( n22989 ) == ( bv_8_71_n252 )  ;
assign n22991 = state_in[79:72] ;
assign n22992 =  ( n22991 ) == ( bv_8_70_n609 )  ;
assign n22993 = state_in[79:72] ;
assign n22994 =  ( n22993 ) == ( bv_8_69_n612 )  ;
assign n22995 = state_in[79:72] ;
assign n22996 =  ( n22995 ) == ( bv_8_68_n390 )  ;
assign n22997 = state_in[79:72] ;
assign n22998 =  ( n22997 ) == ( bv_8_67_n318 )  ;
assign n22999 = state_in[79:72] ;
assign n23000 =  ( n22999 ) == ( bv_8_66_n466 )  ;
assign n23001 = state_in[79:72] ;
assign n23002 =  ( n23001 ) == ( bv_8_65_n623 )  ;
assign n23003 = state_in[79:72] ;
assign n23004 =  ( n23003 ) == ( bv_8_64_n573 )  ;
assign n23005 = state_in[79:72] ;
assign n23006 =  ( n23005 ) == ( bv_8_63_n489 )  ;
assign n23007 = state_in[79:72] ;
assign n23008 =  ( n23007 ) == ( bv_8_62_n205 )  ;
assign n23009 = state_in[79:72] ;
assign n23010 =  ( n23009 ) == ( bv_8_61_n634 )  ;
assign n23011 = state_in[79:72] ;
assign n23012 =  ( n23011 ) == ( bv_8_60_n93 )  ;
assign n23013 = state_in[79:72] ;
assign n23014 =  ( n23013 ) == ( bv_8_59_n382 )  ;
assign n23015 = state_in[79:72] ;
assign n23016 =  ( n23015 ) == ( bv_8_58_n136 )  ;
assign n23017 = state_in[79:72] ;
assign n23018 =  ( n23017 ) == ( bv_8_57_n312 )  ;
assign n23019 = state_in[79:72] ;
assign n23020 =  ( n23019 ) == ( bv_8_56_n230 )  ;
assign n23021 = state_in[79:72] ;
assign n23022 =  ( n23021 ) == ( bv_8_55_n650 )  ;
assign n23023 = state_in[79:72] ;
assign n23024 =  ( n23023 ) == ( bv_8_54_n616 )  ;
assign n23025 = state_in[79:72] ;
assign n23026 =  ( n23025 ) == ( bv_8_53_n436 )  ;
assign n23027 = state_in[79:72] ;
assign n23028 =  ( n23027 ) == ( bv_8_52_n619 )  ;
assign n23029 = state_in[79:72] ;
assign n23030 =  ( n23029 ) == ( bv_8_51_n101 )  ;
assign n23031 = state_in[79:72] ;
assign n23032 =  ( n23031 ) == ( bv_8_50_n408 )  ;
assign n23033 = state_in[79:72] ;
assign n23034 =  ( n23033 ) == ( bv_8_49_n309 )  ;
assign n23035 = state_in[79:72] ;
assign n23036 =  ( n23035 ) == ( bv_8_48_n660 )  ;
assign n23037 = state_in[79:72] ;
assign n23038 =  ( n23037 ) == ( bv_8_47_n652 )  ;
assign n23039 = state_in[79:72] ;
assign n23040 =  ( n23039 ) == ( bv_8_46_n429 )  ;
assign n23041 = state_in[79:72] ;
assign n23042 =  ( n23041 ) == ( bv_8_45_n97 )  ;
assign n23043 = state_in[79:72] ;
assign n23044 =  ( n23043 ) == ( bv_8_44_n5 )  ;
assign n23045 = state_in[79:72] ;
assign n23046 =  ( n23045 ) == ( bv_8_43_n121 )  ;
assign n23047 = state_in[79:72] ;
assign n23048 =  ( n23047 ) == ( bv_8_42_n672 )  ;
assign n23049 = state_in[79:72] ;
assign n23050 =  ( n23049 ) == ( bv_8_41_n29 )  ;
assign n23051 = state_in[79:72] ;
assign n23052 =  ( n23051 ) == ( bv_8_40_n366 )  ;
assign n23053 = state_in[79:72] ;
assign n23054 =  ( n23053 ) == ( bv_8_39_n132 )  ;
assign n23055 = state_in[79:72] ;
assign n23056 =  ( n23055 ) == ( bv_8_38_n444 )  ;
assign n23057 = state_in[79:72] ;
assign n23058 =  ( n23057 ) == ( bv_8_37_n506 )  ;
assign n23059 = state_in[79:72] ;
assign n23060 =  ( n23059 ) == ( bv_8_36_n645 )  ;
assign n23061 = state_in[79:72] ;
assign n23062 =  ( n23061 ) == ( bv_8_35_n696 )  ;
assign n23063 = state_in[79:72] ;
assign n23064 =  ( n23063 ) == ( bv_8_34_n117 )  ;
assign n23065 = state_in[79:72] ;
assign n23066 =  ( n23065 ) == ( bv_8_33_n486 )  ;
assign n23067 = state_in[79:72] ;
assign n23068 =  ( n23067 ) == ( bv_8_32_n463 )  ;
assign n23069 = state_in[79:72] ;
assign n23070 =  ( n23069 ) == ( bv_8_31_n705 )  ;
assign n23071 = state_in[79:72] ;
assign n23072 =  ( n23071 ) == ( bv_8_30_n21 )  ;
assign n23073 = state_in[79:72] ;
assign n23074 =  ( n23073 ) == ( bv_8_29_n625 )  ;
assign n23075 = state_in[79:72] ;
assign n23076 =  ( n23075 ) == ( bv_8_28_n162 )  ;
assign n23077 = state_in[79:72] ;
assign n23078 =  ( n23077 ) == ( bv_8_27_n642 )  ;
assign n23079 = state_in[79:72] ;
assign n23080 =  ( n23079 ) == ( bv_8_26_n53 )  ;
assign n23081 = state_in[79:72] ;
assign n23082 =  ( n23081 ) == ( bv_8_25_n399 )  ;
assign n23083 = state_in[79:72] ;
assign n23084 =  ( n23083 ) == ( bv_8_24_n448 )  ;
assign n23085 = state_in[79:72] ;
assign n23086 =  ( n23085 ) == ( bv_8_23_n144 )  ;
assign n23087 = state_in[79:72] ;
assign n23088 =  ( n23087 ) == ( bv_8_22_n357 )  ;
assign n23089 = state_in[79:72] ;
assign n23090 =  ( n23089 ) == ( bv_8_21_n89 )  ;
assign n23091 = state_in[79:72] ;
assign n23092 =  ( n23091 ) == ( bv_8_20_n341 )  ;
assign n23093 = state_in[79:72] ;
assign n23094 =  ( n23093 ) == ( bv_8_19_n588 )  ;
assign n23095 = state_in[79:72] ;
assign n23096 =  ( n23095 ) == ( bv_8_18_n628 )  ;
assign n23097 = state_in[79:72] ;
assign n23098 =  ( n23097 ) == ( bv_8_17_n525 )  ;
assign n23099 = state_in[79:72] ;
assign n23100 =  ( n23099 ) == ( bv_8_16_n248 )  ;
assign n23101 = state_in[79:72] ;
assign n23102 =  ( n23101 ) == ( bv_8_15_n190 )  ;
assign n23103 = state_in[79:72] ;
assign n23104 =  ( n23103 ) == ( bv_8_14_n648 )  ;
assign n23105 = state_in[79:72] ;
assign n23106 =  ( n23105 ) == ( bv_8_13_n194 )  ;
assign n23107 = state_in[79:72] ;
assign n23108 =  ( n23107 ) == ( bv_8_12_n333 )  ;
assign n23109 = state_in[79:72] ;
assign n23110 =  ( n23109 ) == ( bv_8_11_n379 )  ;
assign n23111 = state_in[79:72] ;
assign n23112 =  ( n23111 ) == ( bv_8_10_n655 )  ;
assign n23113 = state_in[79:72] ;
assign n23114 =  ( n23113 ) == ( bv_8_9_n57 )  ;
assign n23115 = state_in[79:72] ;
assign n23116 =  ( n23115 ) == ( bv_8_8_n669 )  ;
assign n23117 = state_in[79:72] ;
assign n23118 =  ( n23117 ) == ( bv_8_7_n105 )  ;
assign n23119 = state_in[79:72] ;
assign n23120 =  ( n23119 ) == ( bv_8_6_n169 )  ;
assign n23121 = state_in[79:72] ;
assign n23122 =  ( n23121 ) == ( bv_8_5_n492 )  ;
assign n23123 = state_in[79:72] ;
assign n23124 =  ( n23123 ) == ( bv_8_4_n516 )  ;
assign n23125 = state_in[79:72] ;
assign n23126 =  ( n23125 ) == ( bv_8_3_n65 )  ;
assign n23127 = state_in[79:72] ;
assign n23128 =  ( n23127 ) == ( bv_8_2_n751 )  ;
assign n23129 = state_in[79:72] ;
assign n23130 =  ( n23129 ) == ( bv_8_1_n287 )  ;
assign n23131 = state_in[79:72] ;
assign n23132 =  ( n23131 ) == ( bv_8_0_n580 )  ;
assign n23133 =  ( n23132 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n23134 =  ( n23130 ) ? ( bv_8_248_n31 ) : ( n23133 ) ;
assign n23135 =  ( n23128 ) ? ( bv_8_238_n71 ) : ( n23134 ) ;
assign n23136 =  ( n23126 ) ? ( bv_8_246_n39 ) : ( n23135 ) ;
assign n23137 =  ( n23124 ) ? ( bv_8_255_n3 ) : ( n23136 ) ;
assign n23138 =  ( n23122 ) ? ( bv_8_214_n164 ) : ( n23137 ) ;
assign n23139 =  ( n23120 ) ? ( bv_8_222_n134 ) : ( n23138 ) ;
assign n23140 =  ( n23118 ) ? ( bv_8_145_n397 ) : ( n23139 ) ;
assign n23141 =  ( n23116 ) ? ( bv_8_96_n542 ) : ( n23140 ) ;
assign n23142 =  ( n23114 ) ? ( bv_8_2_n751 ) : ( n23141 ) ;
assign n23143 =  ( n23112 ) ? ( bv_8_206_n192 ) : ( n23142 ) ;
assign n23144 =  ( n23110 ) ? ( bv_8_86_n567 ) : ( n23143 ) ;
assign n23145 =  ( n23108 ) ? ( bv_8_231_n99 ) : ( n23144 ) ;
assign n23146 =  ( n23106 ) ? ( bv_8_181_n281 ) : ( n23145 ) ;
assign n23147 =  ( n23104 ) ? ( bv_8_77_n593 ) : ( n23146 ) ;
assign n23148 =  ( n23102 ) ? ( bv_8_236_n79 ) : ( n23147 ) ;
assign n23149 =  ( n23100 ) ? ( bv_8_143_n403 ) : ( n23148 ) ;
assign n23150 =  ( n23098 ) ? ( bv_8_31_n705 ) : ( n23149 ) ;
assign n23151 =  ( n23096 ) ? ( bv_8_137_n421 ) : ( n23150 ) ;
assign n23152 =  ( n23094 ) ? ( bv_8_250_n23 ) : ( n23151 ) ;
assign n23153 =  ( n23092 ) ? ( bv_8_239_n67 ) : ( n23152 ) ;
assign n23154 =  ( n23090 ) ? ( bv_8_178_n292 ) : ( n23153 ) ;
assign n23155 =  ( n23088 ) ? ( bv_8_142_n406 ) : ( n23154 ) ;
assign n23156 =  ( n23086 ) ? ( bv_8_251_n19 ) : ( n23155 ) ;
assign n23157 =  ( n23084 ) ? ( bv_8_65_n623 ) : ( n23156 ) ;
assign n23158 =  ( n23082 ) ? ( bv_8_179_n289 ) : ( n23157 ) ;
assign n23159 =  ( n23080 ) ? ( bv_8_95_n545 ) : ( n23158 ) ;
assign n23160 =  ( n23078 ) ? ( bv_8_69_n612 ) : ( n23159 ) ;
assign n23161 =  ( n23076 ) ? ( bv_8_35_n696 ) : ( n23160 ) ;
assign n23162 =  ( n23074 ) ? ( bv_8_83_n575 ) : ( n23161 ) ;
assign n23163 =  ( n23072 ) ? ( bv_8_228_n111 ) : ( n23162 ) ;
assign n23164 =  ( n23070 ) ? ( bv_8_155_n364 ) : ( n23163 ) ;
assign n23165 =  ( n23068 ) ? ( bv_8_117_n484 ) : ( n23164 ) ;
assign n23166 =  ( n23066 ) ? ( bv_8_225_n123 ) : ( n23165 ) ;
assign n23167 =  ( n23064 ) ? ( bv_8_61_n634 ) : ( n23166 ) ;
assign n23168 =  ( n23062 ) ? ( bv_8_76_n596 ) : ( n23167 ) ;
assign n23169 =  ( n23060 ) ? ( bv_8_108_n510 ) : ( n23168 ) ;
assign n23170 =  ( n23058 ) ? ( bv_8_126_n456 ) : ( n23169 ) ;
assign n23171 =  ( n23056 ) ? ( bv_8_245_n43 ) : ( n23170 ) ;
assign n23172 =  ( n23054 ) ? ( bv_8_131_n440 ) : ( n23171 ) ;
assign n23173 =  ( n23052 ) ? ( bv_8_104_n520 ) : ( n23172 ) ;
assign n23174 =  ( n23050 ) ? ( bv_8_81_n582 ) : ( n23173 ) ;
assign n23175 =  ( n23048 ) ? ( bv_8_209_n182 ) : ( n23174 ) ;
assign n23176 =  ( n23046 ) ? ( bv_8_249_n27 ) : ( n23175 ) ;
assign n23177 =  ( n23044 ) ? ( bv_8_226_n119 ) : ( n23176 ) ;
assign n23178 =  ( n23042 ) ? ( bv_8_171_n314 ) : ( n23177 ) ;
assign n23179 =  ( n23040 ) ? ( bv_8_98_n536 ) : ( n23178 ) ;
assign n23180 =  ( n23038 ) ? ( bv_8_42_n672 ) : ( n23179 ) ;
assign n23181 =  ( n23036 ) ? ( bv_8_8_n669 ) : ( n23180 ) ;
assign n23182 =  ( n23034 ) ? ( bv_8_149_n384 ) : ( n23181 ) ;
assign n23183 =  ( n23032 ) ? ( bv_8_70_n609 ) : ( n23182 ) ;
assign n23184 =  ( n23030 ) ? ( bv_8_157_n359 ) : ( n23183 ) ;
assign n23185 =  ( n23028 ) ? ( bv_8_48_n660 ) : ( n23184 ) ;
assign n23186 =  ( n23026 ) ? ( bv_8_55_n650 ) : ( n23185 ) ;
assign n23187 =  ( n23024 ) ? ( bv_8_10_n655 ) : ( n23186 ) ;
assign n23188 =  ( n23022 ) ? ( bv_8_47_n652 ) : ( n23187 ) ;
assign n23189 =  ( n23020 ) ? ( bv_8_14_n648 ) : ( n23188 ) ;
assign n23190 =  ( n23018 ) ? ( bv_8_36_n645 ) : ( n23189 ) ;
assign n23191 =  ( n23016 ) ? ( bv_8_27_n642 ) : ( n23190 ) ;
assign n23192 =  ( n23014 ) ? ( bv_8_223_n130 ) : ( n23191 ) ;
assign n23193 =  ( n23012 ) ? ( bv_8_205_n196 ) : ( n23192 ) ;
assign n23194 =  ( n23010 ) ? ( bv_8_78_n590 ) : ( n23193 ) ;
assign n23195 =  ( n23008 ) ? ( bv_8_127_n453 ) : ( n23194 ) ;
assign n23196 =  ( n23006 ) ? ( bv_8_234_n87 ) : ( n23195 ) ;
assign n23197 =  ( n23004 ) ? ( bv_8_18_n628 ) : ( n23196 ) ;
assign n23198 =  ( n23002 ) ? ( bv_8_29_n625 ) : ( n23197 ) ;
assign n23199 =  ( n23000 ) ? ( bv_8_88_n562 ) : ( n23198 ) ;
assign n23200 =  ( n22998 ) ? ( bv_8_52_n619 ) : ( n23199 ) ;
assign n23201 =  ( n22996 ) ? ( bv_8_54_n616 ) : ( n23200 ) ;
assign n23202 =  ( n22994 ) ? ( bv_8_220_n142 ) : ( n23201 ) ;
assign n23203 =  ( n22992 ) ? ( bv_8_180_n285 ) : ( n23202 ) ;
assign n23204 =  ( n22990 ) ? ( bv_8_91_n555 ) : ( n23203 ) ;
assign n23205 =  ( n22988 ) ? ( bv_8_164_n335 ) : ( n23204 ) ;
assign n23206 =  ( n22986 ) ? ( bv_8_118_n480 ) : ( n23205 ) ;
assign n23207 =  ( n22984 ) ? ( bv_8_183_n273 ) : ( n23206 ) ;
assign n23208 =  ( n22982 ) ? ( bv_8_125_n459 ) : ( n23207 ) ;
assign n23209 =  ( n22980 ) ? ( bv_8_82_n578 ) : ( n23208 ) ;
assign n23210 =  ( n22978 ) ? ( bv_8_221_n138 ) : ( n23209 ) ;
assign n23211 =  ( n22976 ) ? ( bv_8_94_n548 ) : ( n23210 ) ;
assign n23212 =  ( n22974 ) ? ( bv_8_19_n588 ) : ( n23211 ) ;
assign n23213 =  ( n22972 ) ? ( bv_8_166_n328 ) : ( n23212 ) ;
assign n23214 =  ( n22970 ) ? ( bv_8_185_n266 ) : ( n23213 ) ;
assign n23215 =  ( n22968 ) ? ( bv_8_0_n580 ) : ( n23214 ) ;
assign n23216 =  ( n22966 ) ? ( bv_8_193_n239 ) : ( n23215 ) ;
assign n23217 =  ( n22964 ) ? ( bv_8_64_n573 ) : ( n23216 ) ;
assign n23218 =  ( n22962 ) ? ( bv_8_227_n115 ) : ( n23217 ) ;
assign n23219 =  ( n22960 ) ? ( bv_8_121_n470 ) : ( n23218 ) ;
assign n23220 =  ( n22958 ) ? ( bv_8_182_n277 ) : ( n23219 ) ;
assign n23221 =  ( n22956 ) ? ( bv_8_212_n171 ) : ( n23220 ) ;
assign n23222 =  ( n22954 ) ? ( bv_8_141_n410 ) : ( n23221 ) ;
assign n23223 =  ( n22952 ) ? ( bv_8_103_n523 ) : ( n23222 ) ;
assign n23224 =  ( n22950 ) ? ( bv_8_114_n494 ) : ( n23223 ) ;
assign n23225 =  ( n22948 ) ? ( bv_8_148_n388 ) : ( n23224 ) ;
assign n23226 =  ( n22946 ) ? ( bv_8_152_n374 ) : ( n23225 ) ;
assign n23227 =  ( n22944 ) ? ( bv_8_176_n299 ) : ( n23226 ) ;
assign n23228 =  ( n22942 ) ? ( bv_8_133_n434 ) : ( n23227 ) ;
assign n23229 =  ( n22940 ) ? ( bv_8_187_n260 ) : ( n23228 ) ;
assign n23230 =  ( n22938 ) ? ( bv_8_197_n224 ) : ( n23229 ) ;
assign n23231 =  ( n22936 ) ? ( bv_8_79_n538 ) : ( n23230 ) ;
assign n23232 =  ( n22934 ) ? ( bv_8_237_n75 ) : ( n23231 ) ;
assign n23233 =  ( n22932 ) ? ( bv_8_134_n431 ) : ( n23232 ) ;
assign n23234 =  ( n22930 ) ? ( bv_8_154_n368 ) : ( n23233 ) ;
assign n23235 =  ( n22928 ) ? ( bv_8_102_n527 ) : ( n23234 ) ;
assign n23236 =  ( n22926 ) ? ( bv_8_17_n525 ) : ( n23235 ) ;
assign n23237 =  ( n22924 ) ? ( bv_8_138_n418 ) : ( n23236 ) ;
assign n23238 =  ( n22922 ) ? ( bv_8_233_n91 ) : ( n23237 ) ;
assign n23239 =  ( n22920 ) ? ( bv_8_4_n516 ) : ( n23238 ) ;
assign n23240 =  ( n22918 ) ? ( bv_8_254_n7 ) : ( n23239 ) ;
assign n23241 =  ( n22916 ) ? ( bv_8_160_n350 ) : ( n23240 ) ;
assign n23242 =  ( n22914 ) ? ( bv_8_120_n474 ) : ( n23241 ) ;
assign n23243 =  ( n22912 ) ? ( bv_8_37_n506 ) : ( n23242 ) ;
assign n23244 =  ( n22910 ) ? ( bv_8_75_n503 ) : ( n23243 ) ;
assign n23245 =  ( n22908 ) ? ( bv_8_162_n343 ) : ( n23244 ) ;
assign n23246 =  ( n22906 ) ? ( bv_8_93_n498 ) : ( n23245 ) ;
assign n23247 =  ( n22904 ) ? ( bv_8_128_n450 ) : ( n23246 ) ;
assign n23248 =  ( n22902 ) ? ( bv_8_5_n492 ) : ( n23247 ) ;
assign n23249 =  ( n22900 ) ? ( bv_8_63_n489 ) : ( n23248 ) ;
assign n23250 =  ( n22898 ) ? ( bv_8_33_n486 ) : ( n23249 ) ;
assign n23251 =  ( n22896 ) ? ( bv_8_112_n482 ) : ( n23250 ) ;
assign n23252 =  ( n22894 ) ? ( bv_8_241_n59 ) : ( n23251 ) ;
assign n23253 =  ( n22892 ) ? ( bv_8_99_n476 ) : ( n23252 ) ;
assign n23254 =  ( n22890 ) ? ( bv_8_119_n472 ) : ( n23253 ) ;
assign n23255 =  ( n22888 ) ? ( bv_8_175_n302 ) : ( n23254 ) ;
assign n23256 =  ( n22886 ) ? ( bv_8_66_n466 ) : ( n23255 ) ;
assign n23257 =  ( n22884 ) ? ( bv_8_32_n463 ) : ( n23256 ) ;
assign n23258 =  ( n22882 ) ? ( bv_8_229_n107 ) : ( n23257 ) ;
assign n23259 =  ( n22880 ) ? ( bv_8_253_n11 ) : ( n23258 ) ;
assign n23260 =  ( n22878 ) ? ( bv_8_191_n246 ) : ( n23259 ) ;
assign n23261 =  ( n22876 ) ? ( bv_8_129_n446 ) : ( n23260 ) ;
assign n23262 =  ( n22874 ) ? ( bv_8_24_n448 ) : ( n23261 ) ;
assign n23263 =  ( n22872 ) ? ( bv_8_38_n444 ) : ( n23262 ) ;
assign n23264 =  ( n22870 ) ? ( bv_8_195_n232 ) : ( n23263 ) ;
assign n23265 =  ( n22868 ) ? ( bv_8_190_n250 ) : ( n23264 ) ;
assign n23266 =  ( n22866 ) ? ( bv_8_53_n436 ) : ( n23265 ) ;
assign n23267 =  ( n22864 ) ? ( bv_8_136_n425 ) : ( n23266 ) ;
assign n23268 =  ( n22862 ) ? ( bv_8_46_n429 ) : ( n23267 ) ;
assign n23269 =  ( n22860 ) ? ( bv_8_147_n392 ) : ( n23268 ) ;
assign n23270 =  ( n22858 ) ? ( bv_8_85_n423 ) : ( n23269 ) ;
assign n23271 =  ( n22856 ) ? ( bv_8_252_n15 ) : ( n23270 ) ;
assign n23272 =  ( n22854 ) ? ( bv_8_122_n416 ) : ( n23271 ) ;
assign n23273 =  ( n22852 ) ? ( bv_8_200_n213 ) : ( n23272 ) ;
assign n23274 =  ( n22850 ) ? ( bv_8_186_n263 ) : ( n23273 ) ;
assign n23275 =  ( n22848 ) ? ( bv_8_50_n408 ) : ( n23274 ) ;
assign n23276 =  ( n22846 ) ? ( bv_8_230_n103 ) : ( n23275 ) ;
assign n23277 =  ( n22844 ) ? ( bv_8_192_n242 ) : ( n23276 ) ;
assign n23278 =  ( n22842 ) ? ( bv_8_25_n399 ) : ( n23277 ) ;
assign n23279 =  ( n22840 ) ? ( bv_8_158_n355 ) : ( n23278 ) ;
assign n23280 =  ( n22838 ) ? ( bv_8_163_n339 ) : ( n23279 ) ;
assign n23281 =  ( n22836 ) ? ( bv_8_68_n390 ) : ( n23280 ) ;
assign n23282 =  ( n22834 ) ? ( bv_8_84_n386 ) : ( n23281 ) ;
assign n23283 =  ( n22832 ) ? ( bv_8_59_n382 ) : ( n23282 ) ;
assign n23284 =  ( n22830 ) ? ( bv_8_11_n379 ) : ( n23283 ) ;
assign n23285 =  ( n22828 ) ? ( bv_8_140_n376 ) : ( n23284 ) ;
assign n23286 =  ( n22826 ) ? ( bv_8_199_n216 ) : ( n23285 ) ;
assign n23287 =  ( n22824 ) ? ( bv_8_107_n370 ) : ( n23286 ) ;
assign n23288 =  ( n22822 ) ? ( bv_8_40_n366 ) : ( n23287 ) ;
assign n23289 =  ( n22820 ) ? ( bv_8_167_n325 ) : ( n23288 ) ;
assign n23290 =  ( n22818 ) ? ( bv_8_188_n257 ) : ( n23289 ) ;
assign n23291 =  ( n22816 ) ? ( bv_8_22_n357 ) : ( n23290 ) ;
assign n23292 =  ( n22814 ) ? ( bv_8_173_n307 ) : ( n23291 ) ;
assign n23293 =  ( n22812 ) ? ( bv_8_219_n146 ) : ( n23292 ) ;
assign n23294 =  ( n22810 ) ? ( bv_8_100_n348 ) : ( n23293 ) ;
assign n23295 =  ( n22808 ) ? ( bv_8_116_n345 ) : ( n23294 ) ;
assign n23296 =  ( n22806 ) ? ( bv_8_20_n341 ) : ( n23295 ) ;
assign n23297 =  ( n22804 ) ? ( bv_8_146_n337 ) : ( n23296 ) ;
assign n23298 =  ( n22802 ) ? ( bv_8_12_n333 ) : ( n23297 ) ;
assign n23299 =  ( n22800 ) ? ( bv_8_72_n330 ) : ( n23298 ) ;
assign n23300 =  ( n22798 ) ? ( bv_8_184_n270 ) : ( n23299 ) ;
assign n23301 =  ( n22796 ) ? ( bv_8_159_n323 ) : ( n23300 ) ;
assign n23302 =  ( n22794 ) ? ( bv_8_189_n254 ) : ( n23301 ) ;
assign n23303 =  ( n22792 ) ? ( bv_8_67_n318 ) : ( n23302 ) ;
assign n23304 =  ( n22790 ) ? ( bv_8_196_n228 ) : ( n23303 ) ;
assign n23305 =  ( n22788 ) ? ( bv_8_57_n312 ) : ( n23304 ) ;
assign n23306 =  ( n22786 ) ? ( bv_8_49_n309 ) : ( n23305 ) ;
assign n23307 =  ( n22784 ) ? ( bv_8_211_n175 ) : ( n23306 ) ;
assign n23308 =  ( n22782 ) ? ( bv_8_242_n55 ) : ( n23307 ) ;
assign n23309 =  ( n22780 ) ? ( bv_8_213_n167 ) : ( n23308 ) ;
assign n23310 =  ( n22778 ) ? ( bv_8_139_n297 ) : ( n23309 ) ;
assign n23311 =  ( n22776 ) ? ( bv_8_110_n294 ) : ( n23310 ) ;
assign n23312 =  ( n22774 ) ? ( bv_8_218_n150 ) : ( n23311 ) ;
assign n23313 =  ( n22772 ) ? ( bv_8_1_n287 ) : ( n23312 ) ;
assign n23314 =  ( n22770 ) ? ( bv_8_177_n283 ) : ( n23313 ) ;
assign n23315 =  ( n22768 ) ? ( bv_8_156_n279 ) : ( n23314 ) ;
assign n23316 =  ( n22766 ) ? ( bv_8_73_n275 ) : ( n23315 ) ;
assign n23317 =  ( n22764 ) ? ( bv_8_216_n157 ) : ( n23316 ) ;
assign n23318 =  ( n22762 ) ? ( bv_8_172_n268 ) : ( n23317 ) ;
assign n23319 =  ( n22760 ) ? ( bv_8_243_n51 ) : ( n23318 ) ;
assign n23320 =  ( n22758 ) ? ( bv_8_207_n188 ) : ( n23319 ) ;
assign n23321 =  ( n22756 ) ? ( bv_8_202_n207 ) : ( n23320 ) ;
assign n23322 =  ( n22754 ) ? ( bv_8_244_n47 ) : ( n23321 ) ;
assign n23323 =  ( n22752 ) ? ( bv_8_71_n252 ) : ( n23322 ) ;
assign n23324 =  ( n22750 ) ? ( bv_8_16_n248 ) : ( n23323 ) ;
assign n23325 =  ( n22748 ) ? ( bv_8_111_n244 ) : ( n23324 ) ;
assign n23326 =  ( n22746 ) ? ( bv_8_240_n63 ) : ( n23325 ) ;
assign n23327 =  ( n22744 ) ? ( bv_8_74_n237 ) : ( n23326 ) ;
assign n23328 =  ( n22742 ) ? ( bv_8_92_n234 ) : ( n23327 ) ;
assign n23329 =  ( n22740 ) ? ( bv_8_56_n230 ) : ( n23328 ) ;
assign n23330 =  ( n22738 ) ? ( bv_8_87_n226 ) : ( n23329 ) ;
assign n23331 =  ( n22736 ) ? ( bv_8_115_n222 ) : ( n23330 ) ;
assign n23332 =  ( n22734 ) ? ( bv_8_151_n218 ) : ( n23331 ) ;
assign n23333 =  ( n22732 ) ? ( bv_8_203_n203 ) : ( n23332 ) ;
assign n23334 =  ( n22730 ) ? ( bv_8_161_n211 ) : ( n23333 ) ;
assign n23335 =  ( n22728 ) ? ( bv_8_232_n95 ) : ( n23334 ) ;
assign n23336 =  ( n22726 ) ? ( bv_8_62_n205 ) : ( n23335 ) ;
assign n23337 =  ( n22724 ) ? ( bv_8_150_n201 ) : ( n23336 ) ;
assign n23338 =  ( n22722 ) ? ( bv_8_97_n198 ) : ( n23337 ) ;
assign n23339 =  ( n22720 ) ? ( bv_8_13_n194 ) : ( n23338 ) ;
assign n23340 =  ( n22718 ) ? ( bv_8_15_n190 ) : ( n23339 ) ;
assign n23341 =  ( n22716 ) ? ( bv_8_224_n126 ) : ( n23340 ) ;
assign n23342 =  ( n22714 ) ? ( bv_8_124_n184 ) : ( n23341 ) ;
assign n23343 =  ( n22712 ) ? ( bv_8_113_n180 ) : ( n23342 ) ;
assign n23344 =  ( n22710 ) ? ( bv_8_204_n177 ) : ( n23343 ) ;
assign n23345 =  ( n22708 ) ? ( bv_8_144_n173 ) : ( n23344 ) ;
assign n23346 =  ( n22706 ) ? ( bv_8_6_n169 ) : ( n23345 ) ;
assign n23347 =  ( n22704 ) ? ( bv_8_247_n35 ) : ( n23346 ) ;
assign n23348 =  ( n22702 ) ? ( bv_8_28_n162 ) : ( n23347 ) ;
assign n23349 =  ( n22700 ) ? ( bv_8_194_n159 ) : ( n23348 ) ;
assign n23350 =  ( n22698 ) ? ( bv_8_106_n155 ) : ( n23349 ) ;
assign n23351 =  ( n22696 ) ? ( bv_8_174_n152 ) : ( n23350 ) ;
assign n23352 =  ( n22694 ) ? ( bv_8_105_n148 ) : ( n23351 ) ;
assign n23353 =  ( n22692 ) ? ( bv_8_23_n144 ) : ( n23352 ) ;
assign n23354 =  ( n22690 ) ? ( bv_8_153_n140 ) : ( n23353 ) ;
assign n23355 =  ( n22688 ) ? ( bv_8_58_n136 ) : ( n23354 ) ;
assign n23356 =  ( n22686 ) ? ( bv_8_39_n132 ) : ( n23355 ) ;
assign n23357 =  ( n22684 ) ? ( bv_8_217_n128 ) : ( n23356 ) ;
assign n23358 =  ( n22682 ) ? ( bv_8_235_n83 ) : ( n23357 ) ;
assign n23359 =  ( n22680 ) ? ( bv_8_43_n121 ) : ( n23358 ) ;
assign n23360 =  ( n22678 ) ? ( bv_8_34_n117 ) : ( n23359 ) ;
assign n23361 =  ( n22676 ) ? ( bv_8_210_n113 ) : ( n23360 ) ;
assign n23362 =  ( n22674 ) ? ( bv_8_169_n109 ) : ( n23361 ) ;
assign n23363 =  ( n22672 ) ? ( bv_8_7_n105 ) : ( n23362 ) ;
assign n23364 =  ( n22670 ) ? ( bv_8_51_n101 ) : ( n23363 ) ;
assign n23365 =  ( n22668 ) ? ( bv_8_45_n97 ) : ( n23364 ) ;
assign n23366 =  ( n22666 ) ? ( bv_8_60_n93 ) : ( n23365 ) ;
assign n23367 =  ( n22664 ) ? ( bv_8_21_n89 ) : ( n23366 ) ;
assign n23368 =  ( n22662 ) ? ( bv_8_201_n85 ) : ( n23367 ) ;
assign n23369 =  ( n22660 ) ? ( bv_8_135_n81 ) : ( n23368 ) ;
assign n23370 =  ( n22658 ) ? ( bv_8_170_n77 ) : ( n23369 ) ;
assign n23371 =  ( n22656 ) ? ( bv_8_80_n73 ) : ( n23370 ) ;
assign n23372 =  ( n22654 ) ? ( bv_8_165_n69 ) : ( n23371 ) ;
assign n23373 =  ( n22652 ) ? ( bv_8_3_n65 ) : ( n23372 ) ;
assign n23374 =  ( n22650 ) ? ( bv_8_89_n61 ) : ( n23373 ) ;
assign n23375 =  ( n22648 ) ? ( bv_8_9_n57 ) : ( n23374 ) ;
assign n23376 =  ( n22646 ) ? ( bv_8_26_n53 ) : ( n23375 ) ;
assign n23377 =  ( n22644 ) ? ( bv_8_101_n49 ) : ( n23376 ) ;
assign n23378 =  ( n22642 ) ? ( bv_8_215_n45 ) : ( n23377 ) ;
assign n23379 =  ( n22640 ) ? ( bv_8_132_n41 ) : ( n23378 ) ;
assign n23380 =  ( n22638 ) ? ( bv_8_208_n37 ) : ( n23379 ) ;
assign n23381 =  ( n22636 ) ? ( bv_8_130_n33 ) : ( n23380 ) ;
assign n23382 =  ( n22634 ) ? ( bv_8_41_n29 ) : ( n23381 ) ;
assign n23383 =  ( n22632 ) ? ( bv_8_90_n25 ) : ( n23382 ) ;
assign n23384 =  ( n22630 ) ? ( bv_8_30_n21 ) : ( n23383 ) ;
assign n23385 =  ( n22628 ) ? ( bv_8_123_n17 ) : ( n23384 ) ;
assign n23386 =  ( n22626 ) ? ( bv_8_168_n13 ) : ( n23385 ) ;
assign n23387 =  ( n22624 ) ? ( bv_8_109_n9 ) : ( n23386 ) ;
assign n23388 =  ( n22622 ) ? ( bv_8_44_n5 ) : ( n23387 ) ;
assign n23389 =  ( n22620 ) ^ ( n23388 )  ;
assign n23390 =  ( n23389 ) ^ ( n21846 )  ;
assign n23391 = state_in[31:24] ;
assign n23392 =  ( n23391 ) == ( bv_8_255_n3 )  ;
assign n23393 = state_in[31:24] ;
assign n23394 =  ( n23393 ) == ( bv_8_254_n7 )  ;
assign n23395 = state_in[31:24] ;
assign n23396 =  ( n23395 ) == ( bv_8_253_n11 )  ;
assign n23397 = state_in[31:24] ;
assign n23398 =  ( n23397 ) == ( bv_8_252_n15 )  ;
assign n23399 = state_in[31:24] ;
assign n23400 =  ( n23399 ) == ( bv_8_251_n19 )  ;
assign n23401 = state_in[31:24] ;
assign n23402 =  ( n23401 ) == ( bv_8_250_n23 )  ;
assign n23403 = state_in[31:24] ;
assign n23404 =  ( n23403 ) == ( bv_8_249_n27 )  ;
assign n23405 = state_in[31:24] ;
assign n23406 =  ( n23405 ) == ( bv_8_248_n31 )  ;
assign n23407 = state_in[31:24] ;
assign n23408 =  ( n23407 ) == ( bv_8_247_n35 )  ;
assign n23409 = state_in[31:24] ;
assign n23410 =  ( n23409 ) == ( bv_8_246_n39 )  ;
assign n23411 = state_in[31:24] ;
assign n23412 =  ( n23411 ) == ( bv_8_245_n43 )  ;
assign n23413 = state_in[31:24] ;
assign n23414 =  ( n23413 ) == ( bv_8_244_n47 )  ;
assign n23415 = state_in[31:24] ;
assign n23416 =  ( n23415 ) == ( bv_8_243_n51 )  ;
assign n23417 = state_in[31:24] ;
assign n23418 =  ( n23417 ) == ( bv_8_242_n55 )  ;
assign n23419 = state_in[31:24] ;
assign n23420 =  ( n23419 ) == ( bv_8_241_n59 )  ;
assign n23421 = state_in[31:24] ;
assign n23422 =  ( n23421 ) == ( bv_8_240_n63 )  ;
assign n23423 = state_in[31:24] ;
assign n23424 =  ( n23423 ) == ( bv_8_239_n67 )  ;
assign n23425 = state_in[31:24] ;
assign n23426 =  ( n23425 ) == ( bv_8_238_n71 )  ;
assign n23427 = state_in[31:24] ;
assign n23428 =  ( n23427 ) == ( bv_8_237_n75 )  ;
assign n23429 = state_in[31:24] ;
assign n23430 =  ( n23429 ) == ( bv_8_236_n79 )  ;
assign n23431 = state_in[31:24] ;
assign n23432 =  ( n23431 ) == ( bv_8_235_n83 )  ;
assign n23433 = state_in[31:24] ;
assign n23434 =  ( n23433 ) == ( bv_8_234_n87 )  ;
assign n23435 = state_in[31:24] ;
assign n23436 =  ( n23435 ) == ( bv_8_233_n91 )  ;
assign n23437 = state_in[31:24] ;
assign n23438 =  ( n23437 ) == ( bv_8_232_n95 )  ;
assign n23439 = state_in[31:24] ;
assign n23440 =  ( n23439 ) == ( bv_8_231_n99 )  ;
assign n23441 = state_in[31:24] ;
assign n23442 =  ( n23441 ) == ( bv_8_230_n103 )  ;
assign n23443 = state_in[31:24] ;
assign n23444 =  ( n23443 ) == ( bv_8_229_n107 )  ;
assign n23445 = state_in[31:24] ;
assign n23446 =  ( n23445 ) == ( bv_8_228_n111 )  ;
assign n23447 = state_in[31:24] ;
assign n23448 =  ( n23447 ) == ( bv_8_227_n115 )  ;
assign n23449 = state_in[31:24] ;
assign n23450 =  ( n23449 ) == ( bv_8_226_n119 )  ;
assign n23451 = state_in[31:24] ;
assign n23452 =  ( n23451 ) == ( bv_8_225_n123 )  ;
assign n23453 = state_in[31:24] ;
assign n23454 =  ( n23453 ) == ( bv_8_224_n126 )  ;
assign n23455 = state_in[31:24] ;
assign n23456 =  ( n23455 ) == ( bv_8_223_n130 )  ;
assign n23457 = state_in[31:24] ;
assign n23458 =  ( n23457 ) == ( bv_8_222_n134 )  ;
assign n23459 = state_in[31:24] ;
assign n23460 =  ( n23459 ) == ( bv_8_221_n138 )  ;
assign n23461 = state_in[31:24] ;
assign n23462 =  ( n23461 ) == ( bv_8_220_n142 )  ;
assign n23463 = state_in[31:24] ;
assign n23464 =  ( n23463 ) == ( bv_8_219_n146 )  ;
assign n23465 = state_in[31:24] ;
assign n23466 =  ( n23465 ) == ( bv_8_218_n150 )  ;
assign n23467 = state_in[31:24] ;
assign n23468 =  ( n23467 ) == ( bv_8_217_n128 )  ;
assign n23469 = state_in[31:24] ;
assign n23470 =  ( n23469 ) == ( bv_8_216_n157 )  ;
assign n23471 = state_in[31:24] ;
assign n23472 =  ( n23471 ) == ( bv_8_215_n45 )  ;
assign n23473 = state_in[31:24] ;
assign n23474 =  ( n23473 ) == ( bv_8_214_n164 )  ;
assign n23475 = state_in[31:24] ;
assign n23476 =  ( n23475 ) == ( bv_8_213_n167 )  ;
assign n23477 = state_in[31:24] ;
assign n23478 =  ( n23477 ) == ( bv_8_212_n171 )  ;
assign n23479 = state_in[31:24] ;
assign n23480 =  ( n23479 ) == ( bv_8_211_n175 )  ;
assign n23481 = state_in[31:24] ;
assign n23482 =  ( n23481 ) == ( bv_8_210_n113 )  ;
assign n23483 = state_in[31:24] ;
assign n23484 =  ( n23483 ) == ( bv_8_209_n182 )  ;
assign n23485 = state_in[31:24] ;
assign n23486 =  ( n23485 ) == ( bv_8_208_n37 )  ;
assign n23487 = state_in[31:24] ;
assign n23488 =  ( n23487 ) == ( bv_8_207_n188 )  ;
assign n23489 = state_in[31:24] ;
assign n23490 =  ( n23489 ) == ( bv_8_206_n192 )  ;
assign n23491 = state_in[31:24] ;
assign n23492 =  ( n23491 ) == ( bv_8_205_n196 )  ;
assign n23493 = state_in[31:24] ;
assign n23494 =  ( n23493 ) == ( bv_8_204_n177 )  ;
assign n23495 = state_in[31:24] ;
assign n23496 =  ( n23495 ) == ( bv_8_203_n203 )  ;
assign n23497 = state_in[31:24] ;
assign n23498 =  ( n23497 ) == ( bv_8_202_n207 )  ;
assign n23499 = state_in[31:24] ;
assign n23500 =  ( n23499 ) == ( bv_8_201_n85 )  ;
assign n23501 = state_in[31:24] ;
assign n23502 =  ( n23501 ) == ( bv_8_200_n213 )  ;
assign n23503 = state_in[31:24] ;
assign n23504 =  ( n23503 ) == ( bv_8_199_n216 )  ;
assign n23505 = state_in[31:24] ;
assign n23506 =  ( n23505 ) == ( bv_8_198_n220 )  ;
assign n23507 = state_in[31:24] ;
assign n23508 =  ( n23507 ) == ( bv_8_197_n224 )  ;
assign n23509 = state_in[31:24] ;
assign n23510 =  ( n23509 ) == ( bv_8_196_n228 )  ;
assign n23511 = state_in[31:24] ;
assign n23512 =  ( n23511 ) == ( bv_8_195_n232 )  ;
assign n23513 = state_in[31:24] ;
assign n23514 =  ( n23513 ) == ( bv_8_194_n159 )  ;
assign n23515 = state_in[31:24] ;
assign n23516 =  ( n23515 ) == ( bv_8_193_n239 )  ;
assign n23517 = state_in[31:24] ;
assign n23518 =  ( n23517 ) == ( bv_8_192_n242 )  ;
assign n23519 = state_in[31:24] ;
assign n23520 =  ( n23519 ) == ( bv_8_191_n246 )  ;
assign n23521 = state_in[31:24] ;
assign n23522 =  ( n23521 ) == ( bv_8_190_n250 )  ;
assign n23523 = state_in[31:24] ;
assign n23524 =  ( n23523 ) == ( bv_8_189_n254 )  ;
assign n23525 = state_in[31:24] ;
assign n23526 =  ( n23525 ) == ( bv_8_188_n257 )  ;
assign n23527 = state_in[31:24] ;
assign n23528 =  ( n23527 ) == ( bv_8_187_n260 )  ;
assign n23529 = state_in[31:24] ;
assign n23530 =  ( n23529 ) == ( bv_8_186_n263 )  ;
assign n23531 = state_in[31:24] ;
assign n23532 =  ( n23531 ) == ( bv_8_185_n266 )  ;
assign n23533 = state_in[31:24] ;
assign n23534 =  ( n23533 ) == ( bv_8_184_n270 )  ;
assign n23535 = state_in[31:24] ;
assign n23536 =  ( n23535 ) == ( bv_8_183_n273 )  ;
assign n23537 = state_in[31:24] ;
assign n23538 =  ( n23537 ) == ( bv_8_182_n277 )  ;
assign n23539 = state_in[31:24] ;
assign n23540 =  ( n23539 ) == ( bv_8_181_n281 )  ;
assign n23541 = state_in[31:24] ;
assign n23542 =  ( n23541 ) == ( bv_8_180_n285 )  ;
assign n23543 = state_in[31:24] ;
assign n23544 =  ( n23543 ) == ( bv_8_179_n289 )  ;
assign n23545 = state_in[31:24] ;
assign n23546 =  ( n23545 ) == ( bv_8_178_n292 )  ;
assign n23547 = state_in[31:24] ;
assign n23548 =  ( n23547 ) == ( bv_8_177_n283 )  ;
assign n23549 = state_in[31:24] ;
assign n23550 =  ( n23549 ) == ( bv_8_176_n299 )  ;
assign n23551 = state_in[31:24] ;
assign n23552 =  ( n23551 ) == ( bv_8_175_n302 )  ;
assign n23553 = state_in[31:24] ;
assign n23554 =  ( n23553 ) == ( bv_8_174_n152 )  ;
assign n23555 = state_in[31:24] ;
assign n23556 =  ( n23555 ) == ( bv_8_173_n307 )  ;
assign n23557 = state_in[31:24] ;
assign n23558 =  ( n23557 ) == ( bv_8_172_n268 )  ;
assign n23559 = state_in[31:24] ;
assign n23560 =  ( n23559 ) == ( bv_8_171_n314 )  ;
assign n23561 = state_in[31:24] ;
assign n23562 =  ( n23561 ) == ( bv_8_170_n77 )  ;
assign n23563 = state_in[31:24] ;
assign n23564 =  ( n23563 ) == ( bv_8_169_n109 )  ;
assign n23565 = state_in[31:24] ;
assign n23566 =  ( n23565 ) == ( bv_8_168_n13 )  ;
assign n23567 = state_in[31:24] ;
assign n23568 =  ( n23567 ) == ( bv_8_167_n325 )  ;
assign n23569 = state_in[31:24] ;
assign n23570 =  ( n23569 ) == ( bv_8_166_n328 )  ;
assign n23571 = state_in[31:24] ;
assign n23572 =  ( n23571 ) == ( bv_8_165_n69 )  ;
assign n23573 = state_in[31:24] ;
assign n23574 =  ( n23573 ) == ( bv_8_164_n335 )  ;
assign n23575 = state_in[31:24] ;
assign n23576 =  ( n23575 ) == ( bv_8_163_n339 )  ;
assign n23577 = state_in[31:24] ;
assign n23578 =  ( n23577 ) == ( bv_8_162_n343 )  ;
assign n23579 = state_in[31:24] ;
assign n23580 =  ( n23579 ) == ( bv_8_161_n211 )  ;
assign n23581 = state_in[31:24] ;
assign n23582 =  ( n23581 ) == ( bv_8_160_n350 )  ;
assign n23583 = state_in[31:24] ;
assign n23584 =  ( n23583 ) == ( bv_8_159_n323 )  ;
assign n23585 = state_in[31:24] ;
assign n23586 =  ( n23585 ) == ( bv_8_158_n355 )  ;
assign n23587 = state_in[31:24] ;
assign n23588 =  ( n23587 ) == ( bv_8_157_n359 )  ;
assign n23589 = state_in[31:24] ;
assign n23590 =  ( n23589 ) == ( bv_8_156_n279 )  ;
assign n23591 = state_in[31:24] ;
assign n23592 =  ( n23591 ) == ( bv_8_155_n364 )  ;
assign n23593 = state_in[31:24] ;
assign n23594 =  ( n23593 ) == ( bv_8_154_n368 )  ;
assign n23595 = state_in[31:24] ;
assign n23596 =  ( n23595 ) == ( bv_8_153_n140 )  ;
assign n23597 = state_in[31:24] ;
assign n23598 =  ( n23597 ) == ( bv_8_152_n374 )  ;
assign n23599 = state_in[31:24] ;
assign n23600 =  ( n23599 ) == ( bv_8_151_n218 )  ;
assign n23601 = state_in[31:24] ;
assign n23602 =  ( n23601 ) == ( bv_8_150_n201 )  ;
assign n23603 = state_in[31:24] ;
assign n23604 =  ( n23603 ) == ( bv_8_149_n384 )  ;
assign n23605 = state_in[31:24] ;
assign n23606 =  ( n23605 ) == ( bv_8_148_n388 )  ;
assign n23607 = state_in[31:24] ;
assign n23608 =  ( n23607 ) == ( bv_8_147_n392 )  ;
assign n23609 = state_in[31:24] ;
assign n23610 =  ( n23609 ) == ( bv_8_146_n337 )  ;
assign n23611 = state_in[31:24] ;
assign n23612 =  ( n23611 ) == ( bv_8_145_n397 )  ;
assign n23613 = state_in[31:24] ;
assign n23614 =  ( n23613 ) == ( bv_8_144_n173 )  ;
assign n23615 = state_in[31:24] ;
assign n23616 =  ( n23615 ) == ( bv_8_143_n403 )  ;
assign n23617 = state_in[31:24] ;
assign n23618 =  ( n23617 ) == ( bv_8_142_n406 )  ;
assign n23619 = state_in[31:24] ;
assign n23620 =  ( n23619 ) == ( bv_8_141_n410 )  ;
assign n23621 = state_in[31:24] ;
assign n23622 =  ( n23621 ) == ( bv_8_140_n376 )  ;
assign n23623 = state_in[31:24] ;
assign n23624 =  ( n23623 ) == ( bv_8_139_n297 )  ;
assign n23625 = state_in[31:24] ;
assign n23626 =  ( n23625 ) == ( bv_8_138_n418 )  ;
assign n23627 = state_in[31:24] ;
assign n23628 =  ( n23627 ) == ( bv_8_137_n421 )  ;
assign n23629 = state_in[31:24] ;
assign n23630 =  ( n23629 ) == ( bv_8_136_n425 )  ;
assign n23631 = state_in[31:24] ;
assign n23632 =  ( n23631 ) == ( bv_8_135_n81 )  ;
assign n23633 = state_in[31:24] ;
assign n23634 =  ( n23633 ) == ( bv_8_134_n431 )  ;
assign n23635 = state_in[31:24] ;
assign n23636 =  ( n23635 ) == ( bv_8_133_n434 )  ;
assign n23637 = state_in[31:24] ;
assign n23638 =  ( n23637 ) == ( bv_8_132_n41 )  ;
assign n23639 = state_in[31:24] ;
assign n23640 =  ( n23639 ) == ( bv_8_131_n440 )  ;
assign n23641 = state_in[31:24] ;
assign n23642 =  ( n23641 ) == ( bv_8_130_n33 )  ;
assign n23643 = state_in[31:24] ;
assign n23644 =  ( n23643 ) == ( bv_8_129_n446 )  ;
assign n23645 = state_in[31:24] ;
assign n23646 =  ( n23645 ) == ( bv_8_128_n450 )  ;
assign n23647 = state_in[31:24] ;
assign n23648 =  ( n23647 ) == ( bv_8_127_n453 )  ;
assign n23649 = state_in[31:24] ;
assign n23650 =  ( n23649 ) == ( bv_8_126_n456 )  ;
assign n23651 = state_in[31:24] ;
assign n23652 =  ( n23651 ) == ( bv_8_125_n459 )  ;
assign n23653 = state_in[31:24] ;
assign n23654 =  ( n23653 ) == ( bv_8_124_n184 )  ;
assign n23655 = state_in[31:24] ;
assign n23656 =  ( n23655 ) == ( bv_8_123_n17 )  ;
assign n23657 = state_in[31:24] ;
assign n23658 =  ( n23657 ) == ( bv_8_122_n416 )  ;
assign n23659 = state_in[31:24] ;
assign n23660 =  ( n23659 ) == ( bv_8_121_n470 )  ;
assign n23661 = state_in[31:24] ;
assign n23662 =  ( n23661 ) == ( bv_8_120_n474 )  ;
assign n23663 = state_in[31:24] ;
assign n23664 =  ( n23663 ) == ( bv_8_119_n472 )  ;
assign n23665 = state_in[31:24] ;
assign n23666 =  ( n23665 ) == ( bv_8_118_n480 )  ;
assign n23667 = state_in[31:24] ;
assign n23668 =  ( n23667 ) == ( bv_8_117_n484 )  ;
assign n23669 = state_in[31:24] ;
assign n23670 =  ( n23669 ) == ( bv_8_116_n345 )  ;
assign n23671 = state_in[31:24] ;
assign n23672 =  ( n23671 ) == ( bv_8_115_n222 )  ;
assign n23673 = state_in[31:24] ;
assign n23674 =  ( n23673 ) == ( bv_8_114_n494 )  ;
assign n23675 = state_in[31:24] ;
assign n23676 =  ( n23675 ) == ( bv_8_113_n180 )  ;
assign n23677 = state_in[31:24] ;
assign n23678 =  ( n23677 ) == ( bv_8_112_n482 )  ;
assign n23679 = state_in[31:24] ;
assign n23680 =  ( n23679 ) == ( bv_8_111_n244 )  ;
assign n23681 = state_in[31:24] ;
assign n23682 =  ( n23681 ) == ( bv_8_110_n294 )  ;
assign n23683 = state_in[31:24] ;
assign n23684 =  ( n23683 ) == ( bv_8_109_n9 )  ;
assign n23685 = state_in[31:24] ;
assign n23686 =  ( n23685 ) == ( bv_8_108_n510 )  ;
assign n23687 = state_in[31:24] ;
assign n23688 =  ( n23687 ) == ( bv_8_107_n370 )  ;
assign n23689 = state_in[31:24] ;
assign n23690 =  ( n23689 ) == ( bv_8_106_n155 )  ;
assign n23691 = state_in[31:24] ;
assign n23692 =  ( n23691 ) == ( bv_8_105_n148 )  ;
assign n23693 = state_in[31:24] ;
assign n23694 =  ( n23693 ) == ( bv_8_104_n520 )  ;
assign n23695 = state_in[31:24] ;
assign n23696 =  ( n23695 ) == ( bv_8_103_n523 )  ;
assign n23697 = state_in[31:24] ;
assign n23698 =  ( n23697 ) == ( bv_8_102_n527 )  ;
assign n23699 = state_in[31:24] ;
assign n23700 =  ( n23699 ) == ( bv_8_101_n49 )  ;
assign n23701 = state_in[31:24] ;
assign n23702 =  ( n23701 ) == ( bv_8_100_n348 )  ;
assign n23703 = state_in[31:24] ;
assign n23704 =  ( n23703 ) == ( bv_8_99_n476 )  ;
assign n23705 = state_in[31:24] ;
assign n23706 =  ( n23705 ) == ( bv_8_98_n536 )  ;
assign n23707 = state_in[31:24] ;
assign n23708 =  ( n23707 ) == ( bv_8_97_n198 )  ;
assign n23709 = state_in[31:24] ;
assign n23710 =  ( n23709 ) == ( bv_8_96_n542 )  ;
assign n23711 = state_in[31:24] ;
assign n23712 =  ( n23711 ) == ( bv_8_95_n545 )  ;
assign n23713 = state_in[31:24] ;
assign n23714 =  ( n23713 ) == ( bv_8_94_n548 )  ;
assign n23715 = state_in[31:24] ;
assign n23716 =  ( n23715 ) == ( bv_8_93_n498 )  ;
assign n23717 = state_in[31:24] ;
assign n23718 =  ( n23717 ) == ( bv_8_92_n234 )  ;
assign n23719 = state_in[31:24] ;
assign n23720 =  ( n23719 ) == ( bv_8_91_n555 )  ;
assign n23721 = state_in[31:24] ;
assign n23722 =  ( n23721 ) == ( bv_8_90_n25 )  ;
assign n23723 = state_in[31:24] ;
assign n23724 =  ( n23723 ) == ( bv_8_89_n61 )  ;
assign n23725 = state_in[31:24] ;
assign n23726 =  ( n23725 ) == ( bv_8_88_n562 )  ;
assign n23727 = state_in[31:24] ;
assign n23728 =  ( n23727 ) == ( bv_8_87_n226 )  ;
assign n23729 = state_in[31:24] ;
assign n23730 =  ( n23729 ) == ( bv_8_86_n567 )  ;
assign n23731 = state_in[31:24] ;
assign n23732 =  ( n23731 ) == ( bv_8_85_n423 )  ;
assign n23733 = state_in[31:24] ;
assign n23734 =  ( n23733 ) == ( bv_8_84_n386 )  ;
assign n23735 = state_in[31:24] ;
assign n23736 =  ( n23735 ) == ( bv_8_83_n575 )  ;
assign n23737 = state_in[31:24] ;
assign n23738 =  ( n23737 ) == ( bv_8_82_n578 )  ;
assign n23739 = state_in[31:24] ;
assign n23740 =  ( n23739 ) == ( bv_8_81_n582 )  ;
assign n23741 = state_in[31:24] ;
assign n23742 =  ( n23741 ) == ( bv_8_80_n73 )  ;
assign n23743 = state_in[31:24] ;
assign n23744 =  ( n23743 ) == ( bv_8_79_n538 )  ;
assign n23745 = state_in[31:24] ;
assign n23746 =  ( n23745 ) == ( bv_8_78_n590 )  ;
assign n23747 = state_in[31:24] ;
assign n23748 =  ( n23747 ) == ( bv_8_77_n593 )  ;
assign n23749 = state_in[31:24] ;
assign n23750 =  ( n23749 ) == ( bv_8_76_n596 )  ;
assign n23751 = state_in[31:24] ;
assign n23752 =  ( n23751 ) == ( bv_8_75_n503 )  ;
assign n23753 = state_in[31:24] ;
assign n23754 =  ( n23753 ) == ( bv_8_74_n237 )  ;
assign n23755 = state_in[31:24] ;
assign n23756 =  ( n23755 ) == ( bv_8_73_n275 )  ;
assign n23757 = state_in[31:24] ;
assign n23758 =  ( n23757 ) == ( bv_8_72_n330 )  ;
assign n23759 = state_in[31:24] ;
assign n23760 =  ( n23759 ) == ( bv_8_71_n252 )  ;
assign n23761 = state_in[31:24] ;
assign n23762 =  ( n23761 ) == ( bv_8_70_n609 )  ;
assign n23763 = state_in[31:24] ;
assign n23764 =  ( n23763 ) == ( bv_8_69_n612 )  ;
assign n23765 = state_in[31:24] ;
assign n23766 =  ( n23765 ) == ( bv_8_68_n390 )  ;
assign n23767 = state_in[31:24] ;
assign n23768 =  ( n23767 ) == ( bv_8_67_n318 )  ;
assign n23769 = state_in[31:24] ;
assign n23770 =  ( n23769 ) == ( bv_8_66_n466 )  ;
assign n23771 = state_in[31:24] ;
assign n23772 =  ( n23771 ) == ( bv_8_65_n623 )  ;
assign n23773 = state_in[31:24] ;
assign n23774 =  ( n23773 ) == ( bv_8_64_n573 )  ;
assign n23775 = state_in[31:24] ;
assign n23776 =  ( n23775 ) == ( bv_8_63_n489 )  ;
assign n23777 = state_in[31:24] ;
assign n23778 =  ( n23777 ) == ( bv_8_62_n205 )  ;
assign n23779 = state_in[31:24] ;
assign n23780 =  ( n23779 ) == ( bv_8_61_n634 )  ;
assign n23781 = state_in[31:24] ;
assign n23782 =  ( n23781 ) == ( bv_8_60_n93 )  ;
assign n23783 = state_in[31:24] ;
assign n23784 =  ( n23783 ) == ( bv_8_59_n382 )  ;
assign n23785 = state_in[31:24] ;
assign n23786 =  ( n23785 ) == ( bv_8_58_n136 )  ;
assign n23787 = state_in[31:24] ;
assign n23788 =  ( n23787 ) == ( bv_8_57_n312 )  ;
assign n23789 = state_in[31:24] ;
assign n23790 =  ( n23789 ) == ( bv_8_56_n230 )  ;
assign n23791 = state_in[31:24] ;
assign n23792 =  ( n23791 ) == ( bv_8_55_n650 )  ;
assign n23793 = state_in[31:24] ;
assign n23794 =  ( n23793 ) == ( bv_8_54_n616 )  ;
assign n23795 = state_in[31:24] ;
assign n23796 =  ( n23795 ) == ( bv_8_53_n436 )  ;
assign n23797 = state_in[31:24] ;
assign n23798 =  ( n23797 ) == ( bv_8_52_n619 )  ;
assign n23799 = state_in[31:24] ;
assign n23800 =  ( n23799 ) == ( bv_8_51_n101 )  ;
assign n23801 = state_in[31:24] ;
assign n23802 =  ( n23801 ) == ( bv_8_50_n408 )  ;
assign n23803 = state_in[31:24] ;
assign n23804 =  ( n23803 ) == ( bv_8_49_n309 )  ;
assign n23805 = state_in[31:24] ;
assign n23806 =  ( n23805 ) == ( bv_8_48_n660 )  ;
assign n23807 = state_in[31:24] ;
assign n23808 =  ( n23807 ) == ( bv_8_47_n652 )  ;
assign n23809 = state_in[31:24] ;
assign n23810 =  ( n23809 ) == ( bv_8_46_n429 )  ;
assign n23811 = state_in[31:24] ;
assign n23812 =  ( n23811 ) == ( bv_8_45_n97 )  ;
assign n23813 = state_in[31:24] ;
assign n23814 =  ( n23813 ) == ( bv_8_44_n5 )  ;
assign n23815 = state_in[31:24] ;
assign n23816 =  ( n23815 ) == ( bv_8_43_n121 )  ;
assign n23817 = state_in[31:24] ;
assign n23818 =  ( n23817 ) == ( bv_8_42_n672 )  ;
assign n23819 = state_in[31:24] ;
assign n23820 =  ( n23819 ) == ( bv_8_41_n29 )  ;
assign n23821 = state_in[31:24] ;
assign n23822 =  ( n23821 ) == ( bv_8_40_n366 )  ;
assign n23823 = state_in[31:24] ;
assign n23824 =  ( n23823 ) == ( bv_8_39_n132 )  ;
assign n23825 = state_in[31:24] ;
assign n23826 =  ( n23825 ) == ( bv_8_38_n444 )  ;
assign n23827 = state_in[31:24] ;
assign n23828 =  ( n23827 ) == ( bv_8_37_n506 )  ;
assign n23829 = state_in[31:24] ;
assign n23830 =  ( n23829 ) == ( bv_8_36_n645 )  ;
assign n23831 = state_in[31:24] ;
assign n23832 =  ( n23831 ) == ( bv_8_35_n696 )  ;
assign n23833 = state_in[31:24] ;
assign n23834 =  ( n23833 ) == ( bv_8_34_n117 )  ;
assign n23835 = state_in[31:24] ;
assign n23836 =  ( n23835 ) == ( bv_8_33_n486 )  ;
assign n23837 = state_in[31:24] ;
assign n23838 =  ( n23837 ) == ( bv_8_32_n463 )  ;
assign n23839 = state_in[31:24] ;
assign n23840 =  ( n23839 ) == ( bv_8_31_n705 )  ;
assign n23841 = state_in[31:24] ;
assign n23842 =  ( n23841 ) == ( bv_8_30_n21 )  ;
assign n23843 = state_in[31:24] ;
assign n23844 =  ( n23843 ) == ( bv_8_29_n625 )  ;
assign n23845 = state_in[31:24] ;
assign n23846 =  ( n23845 ) == ( bv_8_28_n162 )  ;
assign n23847 = state_in[31:24] ;
assign n23848 =  ( n23847 ) == ( bv_8_27_n642 )  ;
assign n23849 = state_in[31:24] ;
assign n23850 =  ( n23849 ) == ( bv_8_26_n53 )  ;
assign n23851 = state_in[31:24] ;
assign n23852 =  ( n23851 ) == ( bv_8_25_n399 )  ;
assign n23853 = state_in[31:24] ;
assign n23854 =  ( n23853 ) == ( bv_8_24_n448 )  ;
assign n23855 = state_in[31:24] ;
assign n23856 =  ( n23855 ) == ( bv_8_23_n144 )  ;
assign n23857 = state_in[31:24] ;
assign n23858 =  ( n23857 ) == ( bv_8_22_n357 )  ;
assign n23859 = state_in[31:24] ;
assign n23860 =  ( n23859 ) == ( bv_8_21_n89 )  ;
assign n23861 = state_in[31:24] ;
assign n23862 =  ( n23861 ) == ( bv_8_20_n341 )  ;
assign n23863 = state_in[31:24] ;
assign n23864 =  ( n23863 ) == ( bv_8_19_n588 )  ;
assign n23865 = state_in[31:24] ;
assign n23866 =  ( n23865 ) == ( bv_8_18_n628 )  ;
assign n23867 = state_in[31:24] ;
assign n23868 =  ( n23867 ) == ( bv_8_17_n525 )  ;
assign n23869 = state_in[31:24] ;
assign n23870 =  ( n23869 ) == ( bv_8_16_n248 )  ;
assign n23871 = state_in[31:24] ;
assign n23872 =  ( n23871 ) == ( bv_8_15_n190 )  ;
assign n23873 = state_in[31:24] ;
assign n23874 =  ( n23873 ) == ( bv_8_14_n648 )  ;
assign n23875 = state_in[31:24] ;
assign n23876 =  ( n23875 ) == ( bv_8_13_n194 )  ;
assign n23877 = state_in[31:24] ;
assign n23878 =  ( n23877 ) == ( bv_8_12_n333 )  ;
assign n23879 = state_in[31:24] ;
assign n23880 =  ( n23879 ) == ( bv_8_11_n379 )  ;
assign n23881 = state_in[31:24] ;
assign n23882 =  ( n23881 ) == ( bv_8_10_n655 )  ;
assign n23883 = state_in[31:24] ;
assign n23884 =  ( n23883 ) == ( bv_8_9_n57 )  ;
assign n23885 = state_in[31:24] ;
assign n23886 =  ( n23885 ) == ( bv_8_8_n669 )  ;
assign n23887 = state_in[31:24] ;
assign n23888 =  ( n23887 ) == ( bv_8_7_n105 )  ;
assign n23889 = state_in[31:24] ;
assign n23890 =  ( n23889 ) == ( bv_8_6_n169 )  ;
assign n23891 = state_in[31:24] ;
assign n23892 =  ( n23891 ) == ( bv_8_5_n492 )  ;
assign n23893 = state_in[31:24] ;
assign n23894 =  ( n23893 ) == ( bv_8_4_n516 )  ;
assign n23895 = state_in[31:24] ;
assign n23896 =  ( n23895 ) == ( bv_8_3_n65 )  ;
assign n23897 = state_in[31:24] ;
assign n23898 =  ( n23897 ) == ( bv_8_2_n751 )  ;
assign n23899 = state_in[31:24] ;
assign n23900 =  ( n23899 ) == ( bv_8_1_n287 )  ;
assign n23901 = state_in[31:24] ;
assign n23902 =  ( n23901 ) == ( bv_8_0_n580 )  ;
assign n23903 =  ( n23902 ) ? ( bv_8_99_n476 ) : ( bv_8_0_n580 ) ;
assign n23904 =  ( n23900 ) ? ( bv_8_124_n184 ) : ( n23903 ) ;
assign n23905 =  ( n23898 ) ? ( bv_8_119_n472 ) : ( n23904 ) ;
assign n23906 =  ( n23896 ) ? ( bv_8_123_n17 ) : ( n23905 ) ;
assign n23907 =  ( n23894 ) ? ( bv_8_242_n55 ) : ( n23906 ) ;
assign n23908 =  ( n23892 ) ? ( bv_8_107_n370 ) : ( n23907 ) ;
assign n23909 =  ( n23890 ) ? ( bv_8_111_n244 ) : ( n23908 ) ;
assign n23910 =  ( n23888 ) ? ( bv_8_197_n224 ) : ( n23909 ) ;
assign n23911 =  ( n23886 ) ? ( bv_8_48_n660 ) : ( n23910 ) ;
assign n23912 =  ( n23884 ) ? ( bv_8_1_n287 ) : ( n23911 ) ;
assign n23913 =  ( n23882 ) ? ( bv_8_103_n523 ) : ( n23912 ) ;
assign n23914 =  ( n23880 ) ? ( bv_8_43_n121 ) : ( n23913 ) ;
assign n23915 =  ( n23878 ) ? ( bv_8_254_n7 ) : ( n23914 ) ;
assign n23916 =  ( n23876 ) ? ( bv_8_215_n45 ) : ( n23915 ) ;
assign n23917 =  ( n23874 ) ? ( bv_8_171_n314 ) : ( n23916 ) ;
assign n23918 =  ( n23872 ) ? ( bv_8_118_n480 ) : ( n23917 ) ;
assign n23919 =  ( n23870 ) ? ( bv_8_202_n207 ) : ( n23918 ) ;
assign n23920 =  ( n23868 ) ? ( bv_8_130_n33 ) : ( n23919 ) ;
assign n23921 =  ( n23866 ) ? ( bv_8_201_n85 ) : ( n23920 ) ;
assign n23922 =  ( n23864 ) ? ( bv_8_125_n459 ) : ( n23921 ) ;
assign n23923 =  ( n23862 ) ? ( bv_8_250_n23 ) : ( n23922 ) ;
assign n23924 =  ( n23860 ) ? ( bv_8_89_n61 ) : ( n23923 ) ;
assign n23925 =  ( n23858 ) ? ( bv_8_71_n252 ) : ( n23924 ) ;
assign n23926 =  ( n23856 ) ? ( bv_8_240_n63 ) : ( n23925 ) ;
assign n23927 =  ( n23854 ) ? ( bv_8_173_n307 ) : ( n23926 ) ;
assign n23928 =  ( n23852 ) ? ( bv_8_212_n171 ) : ( n23927 ) ;
assign n23929 =  ( n23850 ) ? ( bv_8_162_n343 ) : ( n23928 ) ;
assign n23930 =  ( n23848 ) ? ( bv_8_175_n302 ) : ( n23929 ) ;
assign n23931 =  ( n23846 ) ? ( bv_8_156_n279 ) : ( n23930 ) ;
assign n23932 =  ( n23844 ) ? ( bv_8_164_n335 ) : ( n23931 ) ;
assign n23933 =  ( n23842 ) ? ( bv_8_114_n494 ) : ( n23932 ) ;
assign n23934 =  ( n23840 ) ? ( bv_8_192_n242 ) : ( n23933 ) ;
assign n23935 =  ( n23838 ) ? ( bv_8_183_n273 ) : ( n23934 ) ;
assign n23936 =  ( n23836 ) ? ( bv_8_253_n11 ) : ( n23935 ) ;
assign n23937 =  ( n23834 ) ? ( bv_8_147_n392 ) : ( n23936 ) ;
assign n23938 =  ( n23832 ) ? ( bv_8_38_n444 ) : ( n23937 ) ;
assign n23939 =  ( n23830 ) ? ( bv_8_54_n616 ) : ( n23938 ) ;
assign n23940 =  ( n23828 ) ? ( bv_8_63_n489 ) : ( n23939 ) ;
assign n23941 =  ( n23826 ) ? ( bv_8_247_n35 ) : ( n23940 ) ;
assign n23942 =  ( n23824 ) ? ( bv_8_204_n177 ) : ( n23941 ) ;
assign n23943 =  ( n23822 ) ? ( bv_8_52_n619 ) : ( n23942 ) ;
assign n23944 =  ( n23820 ) ? ( bv_8_165_n69 ) : ( n23943 ) ;
assign n23945 =  ( n23818 ) ? ( bv_8_229_n107 ) : ( n23944 ) ;
assign n23946 =  ( n23816 ) ? ( bv_8_241_n59 ) : ( n23945 ) ;
assign n23947 =  ( n23814 ) ? ( bv_8_113_n180 ) : ( n23946 ) ;
assign n23948 =  ( n23812 ) ? ( bv_8_216_n157 ) : ( n23947 ) ;
assign n23949 =  ( n23810 ) ? ( bv_8_49_n309 ) : ( n23948 ) ;
assign n23950 =  ( n23808 ) ? ( bv_8_21_n89 ) : ( n23949 ) ;
assign n23951 =  ( n23806 ) ? ( bv_8_4_n516 ) : ( n23950 ) ;
assign n23952 =  ( n23804 ) ? ( bv_8_199_n216 ) : ( n23951 ) ;
assign n23953 =  ( n23802 ) ? ( bv_8_35_n696 ) : ( n23952 ) ;
assign n23954 =  ( n23800 ) ? ( bv_8_195_n232 ) : ( n23953 ) ;
assign n23955 =  ( n23798 ) ? ( bv_8_24_n448 ) : ( n23954 ) ;
assign n23956 =  ( n23796 ) ? ( bv_8_150_n201 ) : ( n23955 ) ;
assign n23957 =  ( n23794 ) ? ( bv_8_5_n492 ) : ( n23956 ) ;
assign n23958 =  ( n23792 ) ? ( bv_8_154_n368 ) : ( n23957 ) ;
assign n23959 =  ( n23790 ) ? ( bv_8_7_n105 ) : ( n23958 ) ;
assign n23960 =  ( n23788 ) ? ( bv_8_18_n628 ) : ( n23959 ) ;
assign n23961 =  ( n23786 ) ? ( bv_8_128_n450 ) : ( n23960 ) ;
assign n23962 =  ( n23784 ) ? ( bv_8_226_n119 ) : ( n23961 ) ;
assign n23963 =  ( n23782 ) ? ( bv_8_235_n83 ) : ( n23962 ) ;
assign n23964 =  ( n23780 ) ? ( bv_8_39_n132 ) : ( n23963 ) ;
assign n23965 =  ( n23778 ) ? ( bv_8_178_n292 ) : ( n23964 ) ;
assign n23966 =  ( n23776 ) ? ( bv_8_117_n484 ) : ( n23965 ) ;
assign n23967 =  ( n23774 ) ? ( bv_8_9_n57 ) : ( n23966 ) ;
assign n23968 =  ( n23772 ) ? ( bv_8_131_n440 ) : ( n23967 ) ;
assign n23969 =  ( n23770 ) ? ( bv_8_44_n5 ) : ( n23968 ) ;
assign n23970 =  ( n23768 ) ? ( bv_8_26_n53 ) : ( n23969 ) ;
assign n23971 =  ( n23766 ) ? ( bv_8_27_n642 ) : ( n23970 ) ;
assign n23972 =  ( n23764 ) ? ( bv_8_110_n294 ) : ( n23971 ) ;
assign n23973 =  ( n23762 ) ? ( bv_8_90_n25 ) : ( n23972 ) ;
assign n23974 =  ( n23760 ) ? ( bv_8_160_n350 ) : ( n23973 ) ;
assign n23975 =  ( n23758 ) ? ( bv_8_82_n578 ) : ( n23974 ) ;
assign n23976 =  ( n23756 ) ? ( bv_8_59_n382 ) : ( n23975 ) ;
assign n23977 =  ( n23754 ) ? ( bv_8_214_n164 ) : ( n23976 ) ;
assign n23978 =  ( n23752 ) ? ( bv_8_179_n289 ) : ( n23977 ) ;
assign n23979 =  ( n23750 ) ? ( bv_8_41_n29 ) : ( n23978 ) ;
assign n23980 =  ( n23748 ) ? ( bv_8_227_n115 ) : ( n23979 ) ;
assign n23981 =  ( n23746 ) ? ( bv_8_47_n652 ) : ( n23980 ) ;
assign n23982 =  ( n23744 ) ? ( bv_8_132_n41 ) : ( n23981 ) ;
assign n23983 =  ( n23742 ) ? ( bv_8_83_n575 ) : ( n23982 ) ;
assign n23984 =  ( n23740 ) ? ( bv_8_209_n182 ) : ( n23983 ) ;
assign n23985 =  ( n23738 ) ? ( bv_8_0_n580 ) : ( n23984 ) ;
assign n23986 =  ( n23736 ) ? ( bv_8_237_n75 ) : ( n23985 ) ;
assign n23987 =  ( n23734 ) ? ( bv_8_32_n463 ) : ( n23986 ) ;
assign n23988 =  ( n23732 ) ? ( bv_8_252_n15 ) : ( n23987 ) ;
assign n23989 =  ( n23730 ) ? ( bv_8_177_n283 ) : ( n23988 ) ;
assign n23990 =  ( n23728 ) ? ( bv_8_91_n555 ) : ( n23989 ) ;
assign n23991 =  ( n23726 ) ? ( bv_8_106_n155 ) : ( n23990 ) ;
assign n23992 =  ( n23724 ) ? ( bv_8_203_n203 ) : ( n23991 ) ;
assign n23993 =  ( n23722 ) ? ( bv_8_190_n250 ) : ( n23992 ) ;
assign n23994 =  ( n23720 ) ? ( bv_8_57_n312 ) : ( n23993 ) ;
assign n23995 =  ( n23718 ) ? ( bv_8_74_n237 ) : ( n23994 ) ;
assign n23996 =  ( n23716 ) ? ( bv_8_76_n596 ) : ( n23995 ) ;
assign n23997 =  ( n23714 ) ? ( bv_8_88_n562 ) : ( n23996 ) ;
assign n23998 =  ( n23712 ) ? ( bv_8_207_n188 ) : ( n23997 ) ;
assign n23999 =  ( n23710 ) ? ( bv_8_208_n37 ) : ( n23998 ) ;
assign n24000 =  ( n23708 ) ? ( bv_8_239_n67 ) : ( n23999 ) ;
assign n24001 =  ( n23706 ) ? ( bv_8_170_n77 ) : ( n24000 ) ;
assign n24002 =  ( n23704 ) ? ( bv_8_251_n19 ) : ( n24001 ) ;
assign n24003 =  ( n23702 ) ? ( bv_8_67_n318 ) : ( n24002 ) ;
assign n24004 =  ( n23700 ) ? ( bv_8_77_n593 ) : ( n24003 ) ;
assign n24005 =  ( n23698 ) ? ( bv_8_51_n101 ) : ( n24004 ) ;
assign n24006 =  ( n23696 ) ? ( bv_8_133_n434 ) : ( n24005 ) ;
assign n24007 =  ( n23694 ) ? ( bv_8_69_n612 ) : ( n24006 ) ;
assign n24008 =  ( n23692 ) ? ( bv_8_249_n27 ) : ( n24007 ) ;
assign n24009 =  ( n23690 ) ? ( bv_8_2_n751 ) : ( n24008 ) ;
assign n24010 =  ( n23688 ) ? ( bv_8_127_n453 ) : ( n24009 ) ;
assign n24011 =  ( n23686 ) ? ( bv_8_80_n73 ) : ( n24010 ) ;
assign n24012 =  ( n23684 ) ? ( bv_8_60_n93 ) : ( n24011 ) ;
assign n24013 =  ( n23682 ) ? ( bv_8_159_n323 ) : ( n24012 ) ;
assign n24014 =  ( n23680 ) ? ( bv_8_168_n13 ) : ( n24013 ) ;
assign n24015 =  ( n23678 ) ? ( bv_8_81_n582 ) : ( n24014 ) ;
assign n24016 =  ( n23676 ) ? ( bv_8_163_n339 ) : ( n24015 ) ;
assign n24017 =  ( n23674 ) ? ( bv_8_64_n573 ) : ( n24016 ) ;
assign n24018 =  ( n23672 ) ? ( bv_8_143_n403 ) : ( n24017 ) ;
assign n24019 =  ( n23670 ) ? ( bv_8_146_n337 ) : ( n24018 ) ;
assign n24020 =  ( n23668 ) ? ( bv_8_157_n359 ) : ( n24019 ) ;
assign n24021 =  ( n23666 ) ? ( bv_8_56_n230 ) : ( n24020 ) ;
assign n24022 =  ( n23664 ) ? ( bv_8_245_n43 ) : ( n24021 ) ;
assign n24023 =  ( n23662 ) ? ( bv_8_188_n257 ) : ( n24022 ) ;
assign n24024 =  ( n23660 ) ? ( bv_8_182_n277 ) : ( n24023 ) ;
assign n24025 =  ( n23658 ) ? ( bv_8_218_n150 ) : ( n24024 ) ;
assign n24026 =  ( n23656 ) ? ( bv_8_33_n486 ) : ( n24025 ) ;
assign n24027 =  ( n23654 ) ? ( bv_8_16_n248 ) : ( n24026 ) ;
assign n24028 =  ( n23652 ) ? ( bv_8_255_n3 ) : ( n24027 ) ;
assign n24029 =  ( n23650 ) ? ( bv_8_243_n51 ) : ( n24028 ) ;
assign n24030 =  ( n23648 ) ? ( bv_8_210_n113 ) : ( n24029 ) ;
assign n24031 =  ( n23646 ) ? ( bv_8_205_n196 ) : ( n24030 ) ;
assign n24032 =  ( n23644 ) ? ( bv_8_12_n333 ) : ( n24031 ) ;
assign n24033 =  ( n23642 ) ? ( bv_8_19_n588 ) : ( n24032 ) ;
assign n24034 =  ( n23640 ) ? ( bv_8_236_n79 ) : ( n24033 ) ;
assign n24035 =  ( n23638 ) ? ( bv_8_95_n545 ) : ( n24034 ) ;
assign n24036 =  ( n23636 ) ? ( bv_8_151_n218 ) : ( n24035 ) ;
assign n24037 =  ( n23634 ) ? ( bv_8_68_n390 ) : ( n24036 ) ;
assign n24038 =  ( n23632 ) ? ( bv_8_23_n144 ) : ( n24037 ) ;
assign n24039 =  ( n23630 ) ? ( bv_8_196_n228 ) : ( n24038 ) ;
assign n24040 =  ( n23628 ) ? ( bv_8_167_n325 ) : ( n24039 ) ;
assign n24041 =  ( n23626 ) ? ( bv_8_126_n456 ) : ( n24040 ) ;
assign n24042 =  ( n23624 ) ? ( bv_8_61_n634 ) : ( n24041 ) ;
assign n24043 =  ( n23622 ) ? ( bv_8_100_n348 ) : ( n24042 ) ;
assign n24044 =  ( n23620 ) ? ( bv_8_93_n498 ) : ( n24043 ) ;
assign n24045 =  ( n23618 ) ? ( bv_8_25_n399 ) : ( n24044 ) ;
assign n24046 =  ( n23616 ) ? ( bv_8_115_n222 ) : ( n24045 ) ;
assign n24047 =  ( n23614 ) ? ( bv_8_96_n542 ) : ( n24046 ) ;
assign n24048 =  ( n23612 ) ? ( bv_8_129_n446 ) : ( n24047 ) ;
assign n24049 =  ( n23610 ) ? ( bv_8_79_n538 ) : ( n24048 ) ;
assign n24050 =  ( n23608 ) ? ( bv_8_220_n142 ) : ( n24049 ) ;
assign n24051 =  ( n23606 ) ? ( bv_8_34_n117 ) : ( n24050 ) ;
assign n24052 =  ( n23604 ) ? ( bv_8_42_n672 ) : ( n24051 ) ;
assign n24053 =  ( n23602 ) ? ( bv_8_144_n173 ) : ( n24052 ) ;
assign n24054 =  ( n23600 ) ? ( bv_8_136_n425 ) : ( n24053 ) ;
assign n24055 =  ( n23598 ) ? ( bv_8_70_n609 ) : ( n24054 ) ;
assign n24056 =  ( n23596 ) ? ( bv_8_238_n71 ) : ( n24055 ) ;
assign n24057 =  ( n23594 ) ? ( bv_8_184_n270 ) : ( n24056 ) ;
assign n24058 =  ( n23592 ) ? ( bv_8_20_n341 ) : ( n24057 ) ;
assign n24059 =  ( n23590 ) ? ( bv_8_222_n134 ) : ( n24058 ) ;
assign n24060 =  ( n23588 ) ? ( bv_8_94_n548 ) : ( n24059 ) ;
assign n24061 =  ( n23586 ) ? ( bv_8_11_n379 ) : ( n24060 ) ;
assign n24062 =  ( n23584 ) ? ( bv_8_219_n146 ) : ( n24061 ) ;
assign n24063 =  ( n23582 ) ? ( bv_8_224_n126 ) : ( n24062 ) ;
assign n24064 =  ( n23580 ) ? ( bv_8_50_n408 ) : ( n24063 ) ;
assign n24065 =  ( n23578 ) ? ( bv_8_58_n136 ) : ( n24064 ) ;
assign n24066 =  ( n23576 ) ? ( bv_8_10_n655 ) : ( n24065 ) ;
assign n24067 =  ( n23574 ) ? ( bv_8_73_n275 ) : ( n24066 ) ;
assign n24068 =  ( n23572 ) ? ( bv_8_6_n169 ) : ( n24067 ) ;
assign n24069 =  ( n23570 ) ? ( bv_8_36_n645 ) : ( n24068 ) ;
assign n24070 =  ( n23568 ) ? ( bv_8_92_n234 ) : ( n24069 ) ;
assign n24071 =  ( n23566 ) ? ( bv_8_194_n159 ) : ( n24070 ) ;
assign n24072 =  ( n23564 ) ? ( bv_8_211_n175 ) : ( n24071 ) ;
assign n24073 =  ( n23562 ) ? ( bv_8_172_n268 ) : ( n24072 ) ;
assign n24074 =  ( n23560 ) ? ( bv_8_98_n536 ) : ( n24073 ) ;
assign n24075 =  ( n23558 ) ? ( bv_8_145_n397 ) : ( n24074 ) ;
assign n24076 =  ( n23556 ) ? ( bv_8_149_n384 ) : ( n24075 ) ;
assign n24077 =  ( n23554 ) ? ( bv_8_228_n111 ) : ( n24076 ) ;
assign n24078 =  ( n23552 ) ? ( bv_8_121_n470 ) : ( n24077 ) ;
assign n24079 =  ( n23550 ) ? ( bv_8_231_n99 ) : ( n24078 ) ;
assign n24080 =  ( n23548 ) ? ( bv_8_200_n213 ) : ( n24079 ) ;
assign n24081 =  ( n23546 ) ? ( bv_8_55_n650 ) : ( n24080 ) ;
assign n24082 =  ( n23544 ) ? ( bv_8_109_n9 ) : ( n24081 ) ;
assign n24083 =  ( n23542 ) ? ( bv_8_141_n410 ) : ( n24082 ) ;
assign n24084 =  ( n23540 ) ? ( bv_8_213_n167 ) : ( n24083 ) ;
assign n24085 =  ( n23538 ) ? ( bv_8_78_n590 ) : ( n24084 ) ;
assign n24086 =  ( n23536 ) ? ( bv_8_169_n109 ) : ( n24085 ) ;
assign n24087 =  ( n23534 ) ? ( bv_8_108_n510 ) : ( n24086 ) ;
assign n24088 =  ( n23532 ) ? ( bv_8_86_n567 ) : ( n24087 ) ;
assign n24089 =  ( n23530 ) ? ( bv_8_244_n47 ) : ( n24088 ) ;
assign n24090 =  ( n23528 ) ? ( bv_8_234_n87 ) : ( n24089 ) ;
assign n24091 =  ( n23526 ) ? ( bv_8_101_n49 ) : ( n24090 ) ;
assign n24092 =  ( n23524 ) ? ( bv_8_122_n416 ) : ( n24091 ) ;
assign n24093 =  ( n23522 ) ? ( bv_8_174_n152 ) : ( n24092 ) ;
assign n24094 =  ( n23520 ) ? ( bv_8_8_n669 ) : ( n24093 ) ;
assign n24095 =  ( n23518 ) ? ( bv_8_186_n263 ) : ( n24094 ) ;
assign n24096 =  ( n23516 ) ? ( bv_8_120_n474 ) : ( n24095 ) ;
assign n24097 =  ( n23514 ) ? ( bv_8_37_n506 ) : ( n24096 ) ;
assign n24098 =  ( n23512 ) ? ( bv_8_46_n429 ) : ( n24097 ) ;
assign n24099 =  ( n23510 ) ? ( bv_8_28_n162 ) : ( n24098 ) ;
assign n24100 =  ( n23508 ) ? ( bv_8_166_n328 ) : ( n24099 ) ;
assign n24101 =  ( n23506 ) ? ( bv_8_180_n285 ) : ( n24100 ) ;
assign n24102 =  ( n23504 ) ? ( bv_8_198_n220 ) : ( n24101 ) ;
assign n24103 =  ( n23502 ) ? ( bv_8_232_n95 ) : ( n24102 ) ;
assign n24104 =  ( n23500 ) ? ( bv_8_221_n138 ) : ( n24103 ) ;
assign n24105 =  ( n23498 ) ? ( bv_8_116_n345 ) : ( n24104 ) ;
assign n24106 =  ( n23496 ) ? ( bv_8_31_n705 ) : ( n24105 ) ;
assign n24107 =  ( n23494 ) ? ( bv_8_75_n503 ) : ( n24106 ) ;
assign n24108 =  ( n23492 ) ? ( bv_8_189_n254 ) : ( n24107 ) ;
assign n24109 =  ( n23490 ) ? ( bv_8_139_n297 ) : ( n24108 ) ;
assign n24110 =  ( n23488 ) ? ( bv_8_138_n418 ) : ( n24109 ) ;
assign n24111 =  ( n23486 ) ? ( bv_8_112_n482 ) : ( n24110 ) ;
assign n24112 =  ( n23484 ) ? ( bv_8_62_n205 ) : ( n24111 ) ;
assign n24113 =  ( n23482 ) ? ( bv_8_181_n281 ) : ( n24112 ) ;
assign n24114 =  ( n23480 ) ? ( bv_8_102_n527 ) : ( n24113 ) ;
assign n24115 =  ( n23478 ) ? ( bv_8_72_n330 ) : ( n24114 ) ;
assign n24116 =  ( n23476 ) ? ( bv_8_3_n65 ) : ( n24115 ) ;
assign n24117 =  ( n23474 ) ? ( bv_8_246_n39 ) : ( n24116 ) ;
assign n24118 =  ( n23472 ) ? ( bv_8_14_n648 ) : ( n24117 ) ;
assign n24119 =  ( n23470 ) ? ( bv_8_97_n198 ) : ( n24118 ) ;
assign n24120 =  ( n23468 ) ? ( bv_8_53_n436 ) : ( n24119 ) ;
assign n24121 =  ( n23466 ) ? ( bv_8_87_n226 ) : ( n24120 ) ;
assign n24122 =  ( n23464 ) ? ( bv_8_185_n266 ) : ( n24121 ) ;
assign n24123 =  ( n23462 ) ? ( bv_8_134_n431 ) : ( n24122 ) ;
assign n24124 =  ( n23460 ) ? ( bv_8_193_n239 ) : ( n24123 ) ;
assign n24125 =  ( n23458 ) ? ( bv_8_29_n625 ) : ( n24124 ) ;
assign n24126 =  ( n23456 ) ? ( bv_8_158_n355 ) : ( n24125 ) ;
assign n24127 =  ( n23454 ) ? ( bv_8_225_n123 ) : ( n24126 ) ;
assign n24128 =  ( n23452 ) ? ( bv_8_248_n31 ) : ( n24127 ) ;
assign n24129 =  ( n23450 ) ? ( bv_8_152_n374 ) : ( n24128 ) ;
assign n24130 =  ( n23448 ) ? ( bv_8_17_n525 ) : ( n24129 ) ;
assign n24131 =  ( n23446 ) ? ( bv_8_105_n148 ) : ( n24130 ) ;
assign n24132 =  ( n23444 ) ? ( bv_8_217_n128 ) : ( n24131 ) ;
assign n24133 =  ( n23442 ) ? ( bv_8_142_n406 ) : ( n24132 ) ;
assign n24134 =  ( n23440 ) ? ( bv_8_148_n388 ) : ( n24133 ) ;
assign n24135 =  ( n23438 ) ? ( bv_8_155_n364 ) : ( n24134 ) ;
assign n24136 =  ( n23436 ) ? ( bv_8_30_n21 ) : ( n24135 ) ;
assign n24137 =  ( n23434 ) ? ( bv_8_135_n81 ) : ( n24136 ) ;
assign n24138 =  ( n23432 ) ? ( bv_8_233_n91 ) : ( n24137 ) ;
assign n24139 =  ( n23430 ) ? ( bv_8_206_n192 ) : ( n24138 ) ;
assign n24140 =  ( n23428 ) ? ( bv_8_85_n423 ) : ( n24139 ) ;
assign n24141 =  ( n23426 ) ? ( bv_8_40_n366 ) : ( n24140 ) ;
assign n24142 =  ( n23424 ) ? ( bv_8_223_n130 ) : ( n24141 ) ;
assign n24143 =  ( n23422 ) ? ( bv_8_140_n376 ) : ( n24142 ) ;
assign n24144 =  ( n23420 ) ? ( bv_8_161_n211 ) : ( n24143 ) ;
assign n24145 =  ( n23418 ) ? ( bv_8_137_n421 ) : ( n24144 ) ;
assign n24146 =  ( n23416 ) ? ( bv_8_13_n194 ) : ( n24145 ) ;
assign n24147 =  ( n23414 ) ? ( bv_8_191_n246 ) : ( n24146 ) ;
assign n24148 =  ( n23412 ) ? ( bv_8_230_n103 ) : ( n24147 ) ;
assign n24149 =  ( n23410 ) ? ( bv_8_66_n466 ) : ( n24148 ) ;
assign n24150 =  ( n23408 ) ? ( bv_8_104_n520 ) : ( n24149 ) ;
assign n24151 =  ( n23406 ) ? ( bv_8_65_n623 ) : ( n24150 ) ;
assign n24152 =  ( n23404 ) ? ( bv_8_153_n140 ) : ( n24151 ) ;
assign n24153 =  ( n23402 ) ? ( bv_8_45_n97 ) : ( n24152 ) ;
assign n24154 =  ( n23400 ) ? ( bv_8_15_n190 ) : ( n24153 ) ;
assign n24155 =  ( n23398 ) ? ( bv_8_176_n299 ) : ( n24154 ) ;
assign n24156 =  ( n23396 ) ? ( bv_8_84_n386 ) : ( n24155 ) ;
assign n24157 =  ( n23394 ) ? ( bv_8_187_n260 ) : ( n24156 ) ;
assign n24158 =  ( n23392 ) ? ( bv_8_22_n357 ) : ( n24157 ) ;
assign n24159 =  ( n23390 ) ^ ( n24158 )  ;
assign n24160 = key[23:16] ;
assign n24161 =  ( n24159 ) ^ ( n24160 )  ;
assign n24162 =  { ( n22619 ) , ( n24161 ) }  ;
assign n24163 =  ( n19540 ) ^ ( n23388 )  ;
assign n24164 =  ( n24163 ) ^ ( n21846 )  ;
assign n24165 = state_in[39:32] ;
assign n24166 =  ( n24165 ) == ( bv_8_255_n3 )  ;
assign n24167 = state_in[39:32] ;
assign n24168 =  ( n24167 ) == ( bv_8_254_n7 )  ;
assign n24169 = state_in[39:32] ;
assign n24170 =  ( n24169 ) == ( bv_8_253_n11 )  ;
assign n24171 = state_in[39:32] ;
assign n24172 =  ( n24171 ) == ( bv_8_252_n15 )  ;
assign n24173 = state_in[39:32] ;
assign n24174 =  ( n24173 ) == ( bv_8_251_n19 )  ;
assign n24175 = state_in[39:32] ;
assign n24176 =  ( n24175 ) == ( bv_8_250_n23 )  ;
assign n24177 = state_in[39:32] ;
assign n24178 =  ( n24177 ) == ( bv_8_249_n27 )  ;
assign n24179 = state_in[39:32] ;
assign n24180 =  ( n24179 ) == ( bv_8_248_n31 )  ;
assign n24181 = state_in[39:32] ;
assign n24182 =  ( n24181 ) == ( bv_8_247_n35 )  ;
assign n24183 = state_in[39:32] ;
assign n24184 =  ( n24183 ) == ( bv_8_246_n39 )  ;
assign n24185 = state_in[39:32] ;
assign n24186 =  ( n24185 ) == ( bv_8_245_n43 )  ;
assign n24187 = state_in[39:32] ;
assign n24188 =  ( n24187 ) == ( bv_8_244_n47 )  ;
assign n24189 = state_in[39:32] ;
assign n24190 =  ( n24189 ) == ( bv_8_243_n51 )  ;
assign n24191 = state_in[39:32] ;
assign n24192 =  ( n24191 ) == ( bv_8_242_n55 )  ;
assign n24193 = state_in[39:32] ;
assign n24194 =  ( n24193 ) == ( bv_8_241_n59 )  ;
assign n24195 = state_in[39:32] ;
assign n24196 =  ( n24195 ) == ( bv_8_240_n63 )  ;
assign n24197 = state_in[39:32] ;
assign n24198 =  ( n24197 ) == ( bv_8_239_n67 )  ;
assign n24199 = state_in[39:32] ;
assign n24200 =  ( n24199 ) == ( bv_8_238_n71 )  ;
assign n24201 = state_in[39:32] ;
assign n24202 =  ( n24201 ) == ( bv_8_237_n75 )  ;
assign n24203 = state_in[39:32] ;
assign n24204 =  ( n24203 ) == ( bv_8_236_n79 )  ;
assign n24205 = state_in[39:32] ;
assign n24206 =  ( n24205 ) == ( bv_8_235_n83 )  ;
assign n24207 = state_in[39:32] ;
assign n24208 =  ( n24207 ) == ( bv_8_234_n87 )  ;
assign n24209 = state_in[39:32] ;
assign n24210 =  ( n24209 ) == ( bv_8_233_n91 )  ;
assign n24211 = state_in[39:32] ;
assign n24212 =  ( n24211 ) == ( bv_8_232_n95 )  ;
assign n24213 = state_in[39:32] ;
assign n24214 =  ( n24213 ) == ( bv_8_231_n99 )  ;
assign n24215 = state_in[39:32] ;
assign n24216 =  ( n24215 ) == ( bv_8_230_n103 )  ;
assign n24217 = state_in[39:32] ;
assign n24218 =  ( n24217 ) == ( bv_8_229_n107 )  ;
assign n24219 = state_in[39:32] ;
assign n24220 =  ( n24219 ) == ( bv_8_228_n111 )  ;
assign n24221 = state_in[39:32] ;
assign n24222 =  ( n24221 ) == ( bv_8_227_n115 )  ;
assign n24223 = state_in[39:32] ;
assign n24224 =  ( n24223 ) == ( bv_8_226_n119 )  ;
assign n24225 = state_in[39:32] ;
assign n24226 =  ( n24225 ) == ( bv_8_225_n123 )  ;
assign n24227 = state_in[39:32] ;
assign n24228 =  ( n24227 ) == ( bv_8_224_n126 )  ;
assign n24229 = state_in[39:32] ;
assign n24230 =  ( n24229 ) == ( bv_8_223_n130 )  ;
assign n24231 = state_in[39:32] ;
assign n24232 =  ( n24231 ) == ( bv_8_222_n134 )  ;
assign n24233 = state_in[39:32] ;
assign n24234 =  ( n24233 ) == ( bv_8_221_n138 )  ;
assign n24235 = state_in[39:32] ;
assign n24236 =  ( n24235 ) == ( bv_8_220_n142 )  ;
assign n24237 = state_in[39:32] ;
assign n24238 =  ( n24237 ) == ( bv_8_219_n146 )  ;
assign n24239 = state_in[39:32] ;
assign n24240 =  ( n24239 ) == ( bv_8_218_n150 )  ;
assign n24241 = state_in[39:32] ;
assign n24242 =  ( n24241 ) == ( bv_8_217_n128 )  ;
assign n24243 = state_in[39:32] ;
assign n24244 =  ( n24243 ) == ( bv_8_216_n157 )  ;
assign n24245 = state_in[39:32] ;
assign n24246 =  ( n24245 ) == ( bv_8_215_n45 )  ;
assign n24247 = state_in[39:32] ;
assign n24248 =  ( n24247 ) == ( bv_8_214_n164 )  ;
assign n24249 = state_in[39:32] ;
assign n24250 =  ( n24249 ) == ( bv_8_213_n167 )  ;
assign n24251 = state_in[39:32] ;
assign n24252 =  ( n24251 ) == ( bv_8_212_n171 )  ;
assign n24253 = state_in[39:32] ;
assign n24254 =  ( n24253 ) == ( bv_8_211_n175 )  ;
assign n24255 = state_in[39:32] ;
assign n24256 =  ( n24255 ) == ( bv_8_210_n113 )  ;
assign n24257 = state_in[39:32] ;
assign n24258 =  ( n24257 ) == ( bv_8_209_n182 )  ;
assign n24259 = state_in[39:32] ;
assign n24260 =  ( n24259 ) == ( bv_8_208_n37 )  ;
assign n24261 = state_in[39:32] ;
assign n24262 =  ( n24261 ) == ( bv_8_207_n188 )  ;
assign n24263 = state_in[39:32] ;
assign n24264 =  ( n24263 ) == ( bv_8_206_n192 )  ;
assign n24265 = state_in[39:32] ;
assign n24266 =  ( n24265 ) == ( bv_8_205_n196 )  ;
assign n24267 = state_in[39:32] ;
assign n24268 =  ( n24267 ) == ( bv_8_204_n177 )  ;
assign n24269 = state_in[39:32] ;
assign n24270 =  ( n24269 ) == ( bv_8_203_n203 )  ;
assign n24271 = state_in[39:32] ;
assign n24272 =  ( n24271 ) == ( bv_8_202_n207 )  ;
assign n24273 = state_in[39:32] ;
assign n24274 =  ( n24273 ) == ( bv_8_201_n85 )  ;
assign n24275 = state_in[39:32] ;
assign n24276 =  ( n24275 ) == ( bv_8_200_n213 )  ;
assign n24277 = state_in[39:32] ;
assign n24278 =  ( n24277 ) == ( bv_8_199_n216 )  ;
assign n24279 = state_in[39:32] ;
assign n24280 =  ( n24279 ) == ( bv_8_198_n220 )  ;
assign n24281 = state_in[39:32] ;
assign n24282 =  ( n24281 ) == ( bv_8_197_n224 )  ;
assign n24283 = state_in[39:32] ;
assign n24284 =  ( n24283 ) == ( bv_8_196_n228 )  ;
assign n24285 = state_in[39:32] ;
assign n24286 =  ( n24285 ) == ( bv_8_195_n232 )  ;
assign n24287 = state_in[39:32] ;
assign n24288 =  ( n24287 ) == ( bv_8_194_n159 )  ;
assign n24289 = state_in[39:32] ;
assign n24290 =  ( n24289 ) == ( bv_8_193_n239 )  ;
assign n24291 = state_in[39:32] ;
assign n24292 =  ( n24291 ) == ( bv_8_192_n242 )  ;
assign n24293 = state_in[39:32] ;
assign n24294 =  ( n24293 ) == ( bv_8_191_n246 )  ;
assign n24295 = state_in[39:32] ;
assign n24296 =  ( n24295 ) == ( bv_8_190_n250 )  ;
assign n24297 = state_in[39:32] ;
assign n24298 =  ( n24297 ) == ( bv_8_189_n254 )  ;
assign n24299 = state_in[39:32] ;
assign n24300 =  ( n24299 ) == ( bv_8_188_n257 )  ;
assign n24301 = state_in[39:32] ;
assign n24302 =  ( n24301 ) == ( bv_8_187_n260 )  ;
assign n24303 = state_in[39:32] ;
assign n24304 =  ( n24303 ) == ( bv_8_186_n263 )  ;
assign n24305 = state_in[39:32] ;
assign n24306 =  ( n24305 ) == ( bv_8_185_n266 )  ;
assign n24307 = state_in[39:32] ;
assign n24308 =  ( n24307 ) == ( bv_8_184_n270 )  ;
assign n24309 = state_in[39:32] ;
assign n24310 =  ( n24309 ) == ( bv_8_183_n273 )  ;
assign n24311 = state_in[39:32] ;
assign n24312 =  ( n24311 ) == ( bv_8_182_n277 )  ;
assign n24313 = state_in[39:32] ;
assign n24314 =  ( n24313 ) == ( bv_8_181_n281 )  ;
assign n24315 = state_in[39:32] ;
assign n24316 =  ( n24315 ) == ( bv_8_180_n285 )  ;
assign n24317 = state_in[39:32] ;
assign n24318 =  ( n24317 ) == ( bv_8_179_n289 )  ;
assign n24319 = state_in[39:32] ;
assign n24320 =  ( n24319 ) == ( bv_8_178_n292 )  ;
assign n24321 = state_in[39:32] ;
assign n24322 =  ( n24321 ) == ( bv_8_177_n283 )  ;
assign n24323 = state_in[39:32] ;
assign n24324 =  ( n24323 ) == ( bv_8_176_n299 )  ;
assign n24325 = state_in[39:32] ;
assign n24326 =  ( n24325 ) == ( bv_8_175_n302 )  ;
assign n24327 = state_in[39:32] ;
assign n24328 =  ( n24327 ) == ( bv_8_174_n152 )  ;
assign n24329 = state_in[39:32] ;
assign n24330 =  ( n24329 ) == ( bv_8_173_n307 )  ;
assign n24331 = state_in[39:32] ;
assign n24332 =  ( n24331 ) == ( bv_8_172_n268 )  ;
assign n24333 = state_in[39:32] ;
assign n24334 =  ( n24333 ) == ( bv_8_171_n314 )  ;
assign n24335 = state_in[39:32] ;
assign n24336 =  ( n24335 ) == ( bv_8_170_n77 )  ;
assign n24337 = state_in[39:32] ;
assign n24338 =  ( n24337 ) == ( bv_8_169_n109 )  ;
assign n24339 = state_in[39:32] ;
assign n24340 =  ( n24339 ) == ( bv_8_168_n13 )  ;
assign n24341 = state_in[39:32] ;
assign n24342 =  ( n24341 ) == ( bv_8_167_n325 )  ;
assign n24343 = state_in[39:32] ;
assign n24344 =  ( n24343 ) == ( bv_8_166_n328 )  ;
assign n24345 = state_in[39:32] ;
assign n24346 =  ( n24345 ) == ( bv_8_165_n69 )  ;
assign n24347 = state_in[39:32] ;
assign n24348 =  ( n24347 ) == ( bv_8_164_n335 )  ;
assign n24349 = state_in[39:32] ;
assign n24350 =  ( n24349 ) == ( bv_8_163_n339 )  ;
assign n24351 = state_in[39:32] ;
assign n24352 =  ( n24351 ) == ( bv_8_162_n343 )  ;
assign n24353 = state_in[39:32] ;
assign n24354 =  ( n24353 ) == ( bv_8_161_n211 )  ;
assign n24355 = state_in[39:32] ;
assign n24356 =  ( n24355 ) == ( bv_8_160_n350 )  ;
assign n24357 = state_in[39:32] ;
assign n24358 =  ( n24357 ) == ( bv_8_159_n323 )  ;
assign n24359 = state_in[39:32] ;
assign n24360 =  ( n24359 ) == ( bv_8_158_n355 )  ;
assign n24361 = state_in[39:32] ;
assign n24362 =  ( n24361 ) == ( bv_8_157_n359 )  ;
assign n24363 = state_in[39:32] ;
assign n24364 =  ( n24363 ) == ( bv_8_156_n279 )  ;
assign n24365 = state_in[39:32] ;
assign n24366 =  ( n24365 ) == ( bv_8_155_n364 )  ;
assign n24367 = state_in[39:32] ;
assign n24368 =  ( n24367 ) == ( bv_8_154_n368 )  ;
assign n24369 = state_in[39:32] ;
assign n24370 =  ( n24369 ) == ( bv_8_153_n140 )  ;
assign n24371 = state_in[39:32] ;
assign n24372 =  ( n24371 ) == ( bv_8_152_n374 )  ;
assign n24373 = state_in[39:32] ;
assign n24374 =  ( n24373 ) == ( bv_8_151_n218 )  ;
assign n24375 = state_in[39:32] ;
assign n24376 =  ( n24375 ) == ( bv_8_150_n201 )  ;
assign n24377 = state_in[39:32] ;
assign n24378 =  ( n24377 ) == ( bv_8_149_n384 )  ;
assign n24379 = state_in[39:32] ;
assign n24380 =  ( n24379 ) == ( bv_8_148_n388 )  ;
assign n24381 = state_in[39:32] ;
assign n24382 =  ( n24381 ) == ( bv_8_147_n392 )  ;
assign n24383 = state_in[39:32] ;
assign n24384 =  ( n24383 ) == ( bv_8_146_n337 )  ;
assign n24385 = state_in[39:32] ;
assign n24386 =  ( n24385 ) == ( bv_8_145_n397 )  ;
assign n24387 = state_in[39:32] ;
assign n24388 =  ( n24387 ) == ( bv_8_144_n173 )  ;
assign n24389 = state_in[39:32] ;
assign n24390 =  ( n24389 ) == ( bv_8_143_n403 )  ;
assign n24391 = state_in[39:32] ;
assign n24392 =  ( n24391 ) == ( bv_8_142_n406 )  ;
assign n24393 = state_in[39:32] ;
assign n24394 =  ( n24393 ) == ( bv_8_141_n410 )  ;
assign n24395 = state_in[39:32] ;
assign n24396 =  ( n24395 ) == ( bv_8_140_n376 )  ;
assign n24397 = state_in[39:32] ;
assign n24398 =  ( n24397 ) == ( bv_8_139_n297 )  ;
assign n24399 = state_in[39:32] ;
assign n24400 =  ( n24399 ) == ( bv_8_138_n418 )  ;
assign n24401 = state_in[39:32] ;
assign n24402 =  ( n24401 ) == ( bv_8_137_n421 )  ;
assign n24403 = state_in[39:32] ;
assign n24404 =  ( n24403 ) == ( bv_8_136_n425 )  ;
assign n24405 = state_in[39:32] ;
assign n24406 =  ( n24405 ) == ( bv_8_135_n81 )  ;
assign n24407 = state_in[39:32] ;
assign n24408 =  ( n24407 ) == ( bv_8_134_n431 )  ;
assign n24409 = state_in[39:32] ;
assign n24410 =  ( n24409 ) == ( bv_8_133_n434 )  ;
assign n24411 = state_in[39:32] ;
assign n24412 =  ( n24411 ) == ( bv_8_132_n41 )  ;
assign n24413 = state_in[39:32] ;
assign n24414 =  ( n24413 ) == ( bv_8_131_n440 )  ;
assign n24415 = state_in[39:32] ;
assign n24416 =  ( n24415 ) == ( bv_8_130_n33 )  ;
assign n24417 = state_in[39:32] ;
assign n24418 =  ( n24417 ) == ( bv_8_129_n446 )  ;
assign n24419 = state_in[39:32] ;
assign n24420 =  ( n24419 ) == ( bv_8_128_n450 )  ;
assign n24421 = state_in[39:32] ;
assign n24422 =  ( n24421 ) == ( bv_8_127_n453 )  ;
assign n24423 = state_in[39:32] ;
assign n24424 =  ( n24423 ) == ( bv_8_126_n456 )  ;
assign n24425 = state_in[39:32] ;
assign n24426 =  ( n24425 ) == ( bv_8_125_n459 )  ;
assign n24427 = state_in[39:32] ;
assign n24428 =  ( n24427 ) == ( bv_8_124_n184 )  ;
assign n24429 = state_in[39:32] ;
assign n24430 =  ( n24429 ) == ( bv_8_123_n17 )  ;
assign n24431 = state_in[39:32] ;
assign n24432 =  ( n24431 ) == ( bv_8_122_n416 )  ;
assign n24433 = state_in[39:32] ;
assign n24434 =  ( n24433 ) == ( bv_8_121_n470 )  ;
assign n24435 = state_in[39:32] ;
assign n24436 =  ( n24435 ) == ( bv_8_120_n474 )  ;
assign n24437 = state_in[39:32] ;
assign n24438 =  ( n24437 ) == ( bv_8_119_n472 )  ;
assign n24439 = state_in[39:32] ;
assign n24440 =  ( n24439 ) == ( bv_8_118_n480 )  ;
assign n24441 = state_in[39:32] ;
assign n24442 =  ( n24441 ) == ( bv_8_117_n484 )  ;
assign n24443 = state_in[39:32] ;
assign n24444 =  ( n24443 ) == ( bv_8_116_n345 )  ;
assign n24445 = state_in[39:32] ;
assign n24446 =  ( n24445 ) == ( bv_8_115_n222 )  ;
assign n24447 = state_in[39:32] ;
assign n24448 =  ( n24447 ) == ( bv_8_114_n494 )  ;
assign n24449 = state_in[39:32] ;
assign n24450 =  ( n24449 ) == ( bv_8_113_n180 )  ;
assign n24451 = state_in[39:32] ;
assign n24452 =  ( n24451 ) == ( bv_8_112_n482 )  ;
assign n24453 = state_in[39:32] ;
assign n24454 =  ( n24453 ) == ( bv_8_111_n244 )  ;
assign n24455 = state_in[39:32] ;
assign n24456 =  ( n24455 ) == ( bv_8_110_n294 )  ;
assign n24457 = state_in[39:32] ;
assign n24458 =  ( n24457 ) == ( bv_8_109_n9 )  ;
assign n24459 = state_in[39:32] ;
assign n24460 =  ( n24459 ) == ( bv_8_108_n510 )  ;
assign n24461 = state_in[39:32] ;
assign n24462 =  ( n24461 ) == ( bv_8_107_n370 )  ;
assign n24463 = state_in[39:32] ;
assign n24464 =  ( n24463 ) == ( bv_8_106_n155 )  ;
assign n24465 = state_in[39:32] ;
assign n24466 =  ( n24465 ) == ( bv_8_105_n148 )  ;
assign n24467 = state_in[39:32] ;
assign n24468 =  ( n24467 ) == ( bv_8_104_n520 )  ;
assign n24469 = state_in[39:32] ;
assign n24470 =  ( n24469 ) == ( bv_8_103_n523 )  ;
assign n24471 = state_in[39:32] ;
assign n24472 =  ( n24471 ) == ( bv_8_102_n527 )  ;
assign n24473 = state_in[39:32] ;
assign n24474 =  ( n24473 ) == ( bv_8_101_n49 )  ;
assign n24475 = state_in[39:32] ;
assign n24476 =  ( n24475 ) == ( bv_8_100_n348 )  ;
assign n24477 = state_in[39:32] ;
assign n24478 =  ( n24477 ) == ( bv_8_99_n476 )  ;
assign n24479 = state_in[39:32] ;
assign n24480 =  ( n24479 ) == ( bv_8_98_n536 )  ;
assign n24481 = state_in[39:32] ;
assign n24482 =  ( n24481 ) == ( bv_8_97_n198 )  ;
assign n24483 = state_in[39:32] ;
assign n24484 =  ( n24483 ) == ( bv_8_96_n542 )  ;
assign n24485 = state_in[39:32] ;
assign n24486 =  ( n24485 ) == ( bv_8_95_n545 )  ;
assign n24487 = state_in[39:32] ;
assign n24488 =  ( n24487 ) == ( bv_8_94_n548 )  ;
assign n24489 = state_in[39:32] ;
assign n24490 =  ( n24489 ) == ( bv_8_93_n498 )  ;
assign n24491 = state_in[39:32] ;
assign n24492 =  ( n24491 ) == ( bv_8_92_n234 )  ;
assign n24493 = state_in[39:32] ;
assign n24494 =  ( n24493 ) == ( bv_8_91_n555 )  ;
assign n24495 = state_in[39:32] ;
assign n24496 =  ( n24495 ) == ( bv_8_90_n25 )  ;
assign n24497 = state_in[39:32] ;
assign n24498 =  ( n24497 ) == ( bv_8_89_n61 )  ;
assign n24499 = state_in[39:32] ;
assign n24500 =  ( n24499 ) == ( bv_8_88_n562 )  ;
assign n24501 = state_in[39:32] ;
assign n24502 =  ( n24501 ) == ( bv_8_87_n226 )  ;
assign n24503 = state_in[39:32] ;
assign n24504 =  ( n24503 ) == ( bv_8_86_n567 )  ;
assign n24505 = state_in[39:32] ;
assign n24506 =  ( n24505 ) == ( bv_8_85_n423 )  ;
assign n24507 = state_in[39:32] ;
assign n24508 =  ( n24507 ) == ( bv_8_84_n386 )  ;
assign n24509 = state_in[39:32] ;
assign n24510 =  ( n24509 ) == ( bv_8_83_n575 )  ;
assign n24511 = state_in[39:32] ;
assign n24512 =  ( n24511 ) == ( bv_8_82_n578 )  ;
assign n24513 = state_in[39:32] ;
assign n24514 =  ( n24513 ) == ( bv_8_81_n582 )  ;
assign n24515 = state_in[39:32] ;
assign n24516 =  ( n24515 ) == ( bv_8_80_n73 )  ;
assign n24517 = state_in[39:32] ;
assign n24518 =  ( n24517 ) == ( bv_8_79_n538 )  ;
assign n24519 = state_in[39:32] ;
assign n24520 =  ( n24519 ) == ( bv_8_78_n590 )  ;
assign n24521 = state_in[39:32] ;
assign n24522 =  ( n24521 ) == ( bv_8_77_n593 )  ;
assign n24523 = state_in[39:32] ;
assign n24524 =  ( n24523 ) == ( bv_8_76_n596 )  ;
assign n24525 = state_in[39:32] ;
assign n24526 =  ( n24525 ) == ( bv_8_75_n503 )  ;
assign n24527 = state_in[39:32] ;
assign n24528 =  ( n24527 ) == ( bv_8_74_n237 )  ;
assign n24529 = state_in[39:32] ;
assign n24530 =  ( n24529 ) == ( bv_8_73_n275 )  ;
assign n24531 = state_in[39:32] ;
assign n24532 =  ( n24531 ) == ( bv_8_72_n330 )  ;
assign n24533 = state_in[39:32] ;
assign n24534 =  ( n24533 ) == ( bv_8_71_n252 )  ;
assign n24535 = state_in[39:32] ;
assign n24536 =  ( n24535 ) == ( bv_8_70_n609 )  ;
assign n24537 = state_in[39:32] ;
assign n24538 =  ( n24537 ) == ( bv_8_69_n612 )  ;
assign n24539 = state_in[39:32] ;
assign n24540 =  ( n24539 ) == ( bv_8_68_n390 )  ;
assign n24541 = state_in[39:32] ;
assign n24542 =  ( n24541 ) == ( bv_8_67_n318 )  ;
assign n24543 = state_in[39:32] ;
assign n24544 =  ( n24543 ) == ( bv_8_66_n466 )  ;
assign n24545 = state_in[39:32] ;
assign n24546 =  ( n24545 ) == ( bv_8_65_n623 )  ;
assign n24547 = state_in[39:32] ;
assign n24548 =  ( n24547 ) == ( bv_8_64_n573 )  ;
assign n24549 = state_in[39:32] ;
assign n24550 =  ( n24549 ) == ( bv_8_63_n489 )  ;
assign n24551 = state_in[39:32] ;
assign n24552 =  ( n24551 ) == ( bv_8_62_n205 )  ;
assign n24553 = state_in[39:32] ;
assign n24554 =  ( n24553 ) == ( bv_8_61_n634 )  ;
assign n24555 = state_in[39:32] ;
assign n24556 =  ( n24555 ) == ( bv_8_60_n93 )  ;
assign n24557 = state_in[39:32] ;
assign n24558 =  ( n24557 ) == ( bv_8_59_n382 )  ;
assign n24559 = state_in[39:32] ;
assign n24560 =  ( n24559 ) == ( bv_8_58_n136 )  ;
assign n24561 = state_in[39:32] ;
assign n24562 =  ( n24561 ) == ( bv_8_57_n312 )  ;
assign n24563 = state_in[39:32] ;
assign n24564 =  ( n24563 ) == ( bv_8_56_n230 )  ;
assign n24565 = state_in[39:32] ;
assign n24566 =  ( n24565 ) == ( bv_8_55_n650 )  ;
assign n24567 = state_in[39:32] ;
assign n24568 =  ( n24567 ) == ( bv_8_54_n616 )  ;
assign n24569 = state_in[39:32] ;
assign n24570 =  ( n24569 ) == ( bv_8_53_n436 )  ;
assign n24571 = state_in[39:32] ;
assign n24572 =  ( n24571 ) == ( bv_8_52_n619 )  ;
assign n24573 = state_in[39:32] ;
assign n24574 =  ( n24573 ) == ( bv_8_51_n101 )  ;
assign n24575 = state_in[39:32] ;
assign n24576 =  ( n24575 ) == ( bv_8_50_n408 )  ;
assign n24577 = state_in[39:32] ;
assign n24578 =  ( n24577 ) == ( bv_8_49_n309 )  ;
assign n24579 = state_in[39:32] ;
assign n24580 =  ( n24579 ) == ( bv_8_48_n660 )  ;
assign n24581 = state_in[39:32] ;
assign n24582 =  ( n24581 ) == ( bv_8_47_n652 )  ;
assign n24583 = state_in[39:32] ;
assign n24584 =  ( n24583 ) == ( bv_8_46_n429 )  ;
assign n24585 = state_in[39:32] ;
assign n24586 =  ( n24585 ) == ( bv_8_45_n97 )  ;
assign n24587 = state_in[39:32] ;
assign n24588 =  ( n24587 ) == ( bv_8_44_n5 )  ;
assign n24589 = state_in[39:32] ;
assign n24590 =  ( n24589 ) == ( bv_8_43_n121 )  ;
assign n24591 = state_in[39:32] ;
assign n24592 =  ( n24591 ) == ( bv_8_42_n672 )  ;
assign n24593 = state_in[39:32] ;
assign n24594 =  ( n24593 ) == ( bv_8_41_n29 )  ;
assign n24595 = state_in[39:32] ;
assign n24596 =  ( n24595 ) == ( bv_8_40_n366 )  ;
assign n24597 = state_in[39:32] ;
assign n24598 =  ( n24597 ) == ( bv_8_39_n132 )  ;
assign n24599 = state_in[39:32] ;
assign n24600 =  ( n24599 ) == ( bv_8_38_n444 )  ;
assign n24601 = state_in[39:32] ;
assign n24602 =  ( n24601 ) == ( bv_8_37_n506 )  ;
assign n24603 = state_in[39:32] ;
assign n24604 =  ( n24603 ) == ( bv_8_36_n645 )  ;
assign n24605 = state_in[39:32] ;
assign n24606 =  ( n24605 ) == ( bv_8_35_n696 )  ;
assign n24607 = state_in[39:32] ;
assign n24608 =  ( n24607 ) == ( bv_8_34_n117 )  ;
assign n24609 = state_in[39:32] ;
assign n24610 =  ( n24609 ) == ( bv_8_33_n486 )  ;
assign n24611 = state_in[39:32] ;
assign n24612 =  ( n24611 ) == ( bv_8_32_n463 )  ;
assign n24613 = state_in[39:32] ;
assign n24614 =  ( n24613 ) == ( bv_8_31_n705 )  ;
assign n24615 = state_in[39:32] ;
assign n24616 =  ( n24615 ) == ( bv_8_30_n21 )  ;
assign n24617 = state_in[39:32] ;
assign n24618 =  ( n24617 ) == ( bv_8_29_n625 )  ;
assign n24619 = state_in[39:32] ;
assign n24620 =  ( n24619 ) == ( bv_8_28_n162 )  ;
assign n24621 = state_in[39:32] ;
assign n24622 =  ( n24621 ) == ( bv_8_27_n642 )  ;
assign n24623 = state_in[39:32] ;
assign n24624 =  ( n24623 ) == ( bv_8_26_n53 )  ;
assign n24625 = state_in[39:32] ;
assign n24626 =  ( n24625 ) == ( bv_8_25_n399 )  ;
assign n24627 = state_in[39:32] ;
assign n24628 =  ( n24627 ) == ( bv_8_24_n448 )  ;
assign n24629 = state_in[39:32] ;
assign n24630 =  ( n24629 ) == ( bv_8_23_n144 )  ;
assign n24631 = state_in[39:32] ;
assign n24632 =  ( n24631 ) == ( bv_8_22_n357 )  ;
assign n24633 = state_in[39:32] ;
assign n24634 =  ( n24633 ) == ( bv_8_21_n89 )  ;
assign n24635 = state_in[39:32] ;
assign n24636 =  ( n24635 ) == ( bv_8_20_n341 )  ;
assign n24637 = state_in[39:32] ;
assign n24638 =  ( n24637 ) == ( bv_8_19_n588 )  ;
assign n24639 = state_in[39:32] ;
assign n24640 =  ( n24639 ) == ( bv_8_18_n628 )  ;
assign n24641 = state_in[39:32] ;
assign n24642 =  ( n24641 ) == ( bv_8_17_n525 )  ;
assign n24643 = state_in[39:32] ;
assign n24644 =  ( n24643 ) == ( bv_8_16_n248 )  ;
assign n24645 = state_in[39:32] ;
assign n24646 =  ( n24645 ) == ( bv_8_15_n190 )  ;
assign n24647 = state_in[39:32] ;
assign n24648 =  ( n24647 ) == ( bv_8_14_n648 )  ;
assign n24649 = state_in[39:32] ;
assign n24650 =  ( n24649 ) == ( bv_8_13_n194 )  ;
assign n24651 = state_in[39:32] ;
assign n24652 =  ( n24651 ) == ( bv_8_12_n333 )  ;
assign n24653 = state_in[39:32] ;
assign n24654 =  ( n24653 ) == ( bv_8_11_n379 )  ;
assign n24655 = state_in[39:32] ;
assign n24656 =  ( n24655 ) == ( bv_8_10_n655 )  ;
assign n24657 = state_in[39:32] ;
assign n24658 =  ( n24657 ) == ( bv_8_9_n57 )  ;
assign n24659 = state_in[39:32] ;
assign n24660 =  ( n24659 ) == ( bv_8_8_n669 )  ;
assign n24661 = state_in[39:32] ;
assign n24662 =  ( n24661 ) == ( bv_8_7_n105 )  ;
assign n24663 = state_in[39:32] ;
assign n24664 =  ( n24663 ) == ( bv_8_6_n169 )  ;
assign n24665 = state_in[39:32] ;
assign n24666 =  ( n24665 ) == ( bv_8_5_n492 )  ;
assign n24667 = state_in[39:32] ;
assign n24668 =  ( n24667 ) == ( bv_8_4_n516 )  ;
assign n24669 = state_in[39:32] ;
assign n24670 =  ( n24669 ) == ( bv_8_3_n65 )  ;
assign n24671 = state_in[39:32] ;
assign n24672 =  ( n24671 ) == ( bv_8_2_n751 )  ;
assign n24673 = state_in[39:32] ;
assign n24674 =  ( n24673 ) == ( bv_8_1_n287 )  ;
assign n24675 = state_in[39:32] ;
assign n24676 =  ( n24675 ) == ( bv_8_0_n580 )  ;
assign n24677 =  ( n24676 ) ? ( bv_8_198_n220 ) : ( bv_8_0_n580 ) ;
assign n24678 =  ( n24674 ) ? ( bv_8_248_n31 ) : ( n24677 ) ;
assign n24679 =  ( n24672 ) ? ( bv_8_238_n71 ) : ( n24678 ) ;
assign n24680 =  ( n24670 ) ? ( bv_8_246_n39 ) : ( n24679 ) ;
assign n24681 =  ( n24668 ) ? ( bv_8_255_n3 ) : ( n24680 ) ;
assign n24682 =  ( n24666 ) ? ( bv_8_214_n164 ) : ( n24681 ) ;
assign n24683 =  ( n24664 ) ? ( bv_8_222_n134 ) : ( n24682 ) ;
assign n24684 =  ( n24662 ) ? ( bv_8_145_n397 ) : ( n24683 ) ;
assign n24685 =  ( n24660 ) ? ( bv_8_96_n542 ) : ( n24684 ) ;
assign n24686 =  ( n24658 ) ? ( bv_8_2_n751 ) : ( n24685 ) ;
assign n24687 =  ( n24656 ) ? ( bv_8_206_n192 ) : ( n24686 ) ;
assign n24688 =  ( n24654 ) ? ( bv_8_86_n567 ) : ( n24687 ) ;
assign n24689 =  ( n24652 ) ? ( bv_8_231_n99 ) : ( n24688 ) ;
assign n24690 =  ( n24650 ) ? ( bv_8_181_n281 ) : ( n24689 ) ;
assign n24691 =  ( n24648 ) ? ( bv_8_77_n593 ) : ( n24690 ) ;
assign n24692 =  ( n24646 ) ? ( bv_8_236_n79 ) : ( n24691 ) ;
assign n24693 =  ( n24644 ) ? ( bv_8_143_n403 ) : ( n24692 ) ;
assign n24694 =  ( n24642 ) ? ( bv_8_31_n705 ) : ( n24693 ) ;
assign n24695 =  ( n24640 ) ? ( bv_8_137_n421 ) : ( n24694 ) ;
assign n24696 =  ( n24638 ) ? ( bv_8_250_n23 ) : ( n24695 ) ;
assign n24697 =  ( n24636 ) ? ( bv_8_239_n67 ) : ( n24696 ) ;
assign n24698 =  ( n24634 ) ? ( bv_8_178_n292 ) : ( n24697 ) ;
assign n24699 =  ( n24632 ) ? ( bv_8_142_n406 ) : ( n24698 ) ;
assign n24700 =  ( n24630 ) ? ( bv_8_251_n19 ) : ( n24699 ) ;
assign n24701 =  ( n24628 ) ? ( bv_8_65_n623 ) : ( n24700 ) ;
assign n24702 =  ( n24626 ) ? ( bv_8_179_n289 ) : ( n24701 ) ;
assign n24703 =  ( n24624 ) ? ( bv_8_95_n545 ) : ( n24702 ) ;
assign n24704 =  ( n24622 ) ? ( bv_8_69_n612 ) : ( n24703 ) ;
assign n24705 =  ( n24620 ) ? ( bv_8_35_n696 ) : ( n24704 ) ;
assign n24706 =  ( n24618 ) ? ( bv_8_83_n575 ) : ( n24705 ) ;
assign n24707 =  ( n24616 ) ? ( bv_8_228_n111 ) : ( n24706 ) ;
assign n24708 =  ( n24614 ) ? ( bv_8_155_n364 ) : ( n24707 ) ;
assign n24709 =  ( n24612 ) ? ( bv_8_117_n484 ) : ( n24708 ) ;
assign n24710 =  ( n24610 ) ? ( bv_8_225_n123 ) : ( n24709 ) ;
assign n24711 =  ( n24608 ) ? ( bv_8_61_n634 ) : ( n24710 ) ;
assign n24712 =  ( n24606 ) ? ( bv_8_76_n596 ) : ( n24711 ) ;
assign n24713 =  ( n24604 ) ? ( bv_8_108_n510 ) : ( n24712 ) ;
assign n24714 =  ( n24602 ) ? ( bv_8_126_n456 ) : ( n24713 ) ;
assign n24715 =  ( n24600 ) ? ( bv_8_245_n43 ) : ( n24714 ) ;
assign n24716 =  ( n24598 ) ? ( bv_8_131_n440 ) : ( n24715 ) ;
assign n24717 =  ( n24596 ) ? ( bv_8_104_n520 ) : ( n24716 ) ;
assign n24718 =  ( n24594 ) ? ( bv_8_81_n582 ) : ( n24717 ) ;
assign n24719 =  ( n24592 ) ? ( bv_8_209_n182 ) : ( n24718 ) ;
assign n24720 =  ( n24590 ) ? ( bv_8_249_n27 ) : ( n24719 ) ;
assign n24721 =  ( n24588 ) ? ( bv_8_226_n119 ) : ( n24720 ) ;
assign n24722 =  ( n24586 ) ? ( bv_8_171_n314 ) : ( n24721 ) ;
assign n24723 =  ( n24584 ) ? ( bv_8_98_n536 ) : ( n24722 ) ;
assign n24724 =  ( n24582 ) ? ( bv_8_42_n672 ) : ( n24723 ) ;
assign n24725 =  ( n24580 ) ? ( bv_8_8_n669 ) : ( n24724 ) ;
assign n24726 =  ( n24578 ) ? ( bv_8_149_n384 ) : ( n24725 ) ;
assign n24727 =  ( n24576 ) ? ( bv_8_70_n609 ) : ( n24726 ) ;
assign n24728 =  ( n24574 ) ? ( bv_8_157_n359 ) : ( n24727 ) ;
assign n24729 =  ( n24572 ) ? ( bv_8_48_n660 ) : ( n24728 ) ;
assign n24730 =  ( n24570 ) ? ( bv_8_55_n650 ) : ( n24729 ) ;
assign n24731 =  ( n24568 ) ? ( bv_8_10_n655 ) : ( n24730 ) ;
assign n24732 =  ( n24566 ) ? ( bv_8_47_n652 ) : ( n24731 ) ;
assign n24733 =  ( n24564 ) ? ( bv_8_14_n648 ) : ( n24732 ) ;
assign n24734 =  ( n24562 ) ? ( bv_8_36_n645 ) : ( n24733 ) ;
assign n24735 =  ( n24560 ) ? ( bv_8_27_n642 ) : ( n24734 ) ;
assign n24736 =  ( n24558 ) ? ( bv_8_223_n130 ) : ( n24735 ) ;
assign n24737 =  ( n24556 ) ? ( bv_8_205_n196 ) : ( n24736 ) ;
assign n24738 =  ( n24554 ) ? ( bv_8_78_n590 ) : ( n24737 ) ;
assign n24739 =  ( n24552 ) ? ( bv_8_127_n453 ) : ( n24738 ) ;
assign n24740 =  ( n24550 ) ? ( bv_8_234_n87 ) : ( n24739 ) ;
assign n24741 =  ( n24548 ) ? ( bv_8_18_n628 ) : ( n24740 ) ;
assign n24742 =  ( n24546 ) ? ( bv_8_29_n625 ) : ( n24741 ) ;
assign n24743 =  ( n24544 ) ? ( bv_8_88_n562 ) : ( n24742 ) ;
assign n24744 =  ( n24542 ) ? ( bv_8_52_n619 ) : ( n24743 ) ;
assign n24745 =  ( n24540 ) ? ( bv_8_54_n616 ) : ( n24744 ) ;
assign n24746 =  ( n24538 ) ? ( bv_8_220_n142 ) : ( n24745 ) ;
assign n24747 =  ( n24536 ) ? ( bv_8_180_n285 ) : ( n24746 ) ;
assign n24748 =  ( n24534 ) ? ( bv_8_91_n555 ) : ( n24747 ) ;
assign n24749 =  ( n24532 ) ? ( bv_8_164_n335 ) : ( n24748 ) ;
assign n24750 =  ( n24530 ) ? ( bv_8_118_n480 ) : ( n24749 ) ;
assign n24751 =  ( n24528 ) ? ( bv_8_183_n273 ) : ( n24750 ) ;
assign n24752 =  ( n24526 ) ? ( bv_8_125_n459 ) : ( n24751 ) ;
assign n24753 =  ( n24524 ) ? ( bv_8_82_n578 ) : ( n24752 ) ;
assign n24754 =  ( n24522 ) ? ( bv_8_221_n138 ) : ( n24753 ) ;
assign n24755 =  ( n24520 ) ? ( bv_8_94_n548 ) : ( n24754 ) ;
assign n24756 =  ( n24518 ) ? ( bv_8_19_n588 ) : ( n24755 ) ;
assign n24757 =  ( n24516 ) ? ( bv_8_166_n328 ) : ( n24756 ) ;
assign n24758 =  ( n24514 ) ? ( bv_8_185_n266 ) : ( n24757 ) ;
assign n24759 =  ( n24512 ) ? ( bv_8_0_n580 ) : ( n24758 ) ;
assign n24760 =  ( n24510 ) ? ( bv_8_193_n239 ) : ( n24759 ) ;
assign n24761 =  ( n24508 ) ? ( bv_8_64_n573 ) : ( n24760 ) ;
assign n24762 =  ( n24506 ) ? ( bv_8_227_n115 ) : ( n24761 ) ;
assign n24763 =  ( n24504 ) ? ( bv_8_121_n470 ) : ( n24762 ) ;
assign n24764 =  ( n24502 ) ? ( bv_8_182_n277 ) : ( n24763 ) ;
assign n24765 =  ( n24500 ) ? ( bv_8_212_n171 ) : ( n24764 ) ;
assign n24766 =  ( n24498 ) ? ( bv_8_141_n410 ) : ( n24765 ) ;
assign n24767 =  ( n24496 ) ? ( bv_8_103_n523 ) : ( n24766 ) ;
assign n24768 =  ( n24494 ) ? ( bv_8_114_n494 ) : ( n24767 ) ;
assign n24769 =  ( n24492 ) ? ( bv_8_148_n388 ) : ( n24768 ) ;
assign n24770 =  ( n24490 ) ? ( bv_8_152_n374 ) : ( n24769 ) ;
assign n24771 =  ( n24488 ) ? ( bv_8_176_n299 ) : ( n24770 ) ;
assign n24772 =  ( n24486 ) ? ( bv_8_133_n434 ) : ( n24771 ) ;
assign n24773 =  ( n24484 ) ? ( bv_8_187_n260 ) : ( n24772 ) ;
assign n24774 =  ( n24482 ) ? ( bv_8_197_n224 ) : ( n24773 ) ;
assign n24775 =  ( n24480 ) ? ( bv_8_79_n538 ) : ( n24774 ) ;
assign n24776 =  ( n24478 ) ? ( bv_8_237_n75 ) : ( n24775 ) ;
assign n24777 =  ( n24476 ) ? ( bv_8_134_n431 ) : ( n24776 ) ;
assign n24778 =  ( n24474 ) ? ( bv_8_154_n368 ) : ( n24777 ) ;
assign n24779 =  ( n24472 ) ? ( bv_8_102_n527 ) : ( n24778 ) ;
assign n24780 =  ( n24470 ) ? ( bv_8_17_n525 ) : ( n24779 ) ;
assign n24781 =  ( n24468 ) ? ( bv_8_138_n418 ) : ( n24780 ) ;
assign n24782 =  ( n24466 ) ? ( bv_8_233_n91 ) : ( n24781 ) ;
assign n24783 =  ( n24464 ) ? ( bv_8_4_n516 ) : ( n24782 ) ;
assign n24784 =  ( n24462 ) ? ( bv_8_254_n7 ) : ( n24783 ) ;
assign n24785 =  ( n24460 ) ? ( bv_8_160_n350 ) : ( n24784 ) ;
assign n24786 =  ( n24458 ) ? ( bv_8_120_n474 ) : ( n24785 ) ;
assign n24787 =  ( n24456 ) ? ( bv_8_37_n506 ) : ( n24786 ) ;
assign n24788 =  ( n24454 ) ? ( bv_8_75_n503 ) : ( n24787 ) ;
assign n24789 =  ( n24452 ) ? ( bv_8_162_n343 ) : ( n24788 ) ;
assign n24790 =  ( n24450 ) ? ( bv_8_93_n498 ) : ( n24789 ) ;
assign n24791 =  ( n24448 ) ? ( bv_8_128_n450 ) : ( n24790 ) ;
assign n24792 =  ( n24446 ) ? ( bv_8_5_n492 ) : ( n24791 ) ;
assign n24793 =  ( n24444 ) ? ( bv_8_63_n489 ) : ( n24792 ) ;
assign n24794 =  ( n24442 ) ? ( bv_8_33_n486 ) : ( n24793 ) ;
assign n24795 =  ( n24440 ) ? ( bv_8_112_n482 ) : ( n24794 ) ;
assign n24796 =  ( n24438 ) ? ( bv_8_241_n59 ) : ( n24795 ) ;
assign n24797 =  ( n24436 ) ? ( bv_8_99_n476 ) : ( n24796 ) ;
assign n24798 =  ( n24434 ) ? ( bv_8_119_n472 ) : ( n24797 ) ;
assign n24799 =  ( n24432 ) ? ( bv_8_175_n302 ) : ( n24798 ) ;
assign n24800 =  ( n24430 ) ? ( bv_8_66_n466 ) : ( n24799 ) ;
assign n24801 =  ( n24428 ) ? ( bv_8_32_n463 ) : ( n24800 ) ;
assign n24802 =  ( n24426 ) ? ( bv_8_229_n107 ) : ( n24801 ) ;
assign n24803 =  ( n24424 ) ? ( bv_8_253_n11 ) : ( n24802 ) ;
assign n24804 =  ( n24422 ) ? ( bv_8_191_n246 ) : ( n24803 ) ;
assign n24805 =  ( n24420 ) ? ( bv_8_129_n446 ) : ( n24804 ) ;
assign n24806 =  ( n24418 ) ? ( bv_8_24_n448 ) : ( n24805 ) ;
assign n24807 =  ( n24416 ) ? ( bv_8_38_n444 ) : ( n24806 ) ;
assign n24808 =  ( n24414 ) ? ( bv_8_195_n232 ) : ( n24807 ) ;
assign n24809 =  ( n24412 ) ? ( bv_8_190_n250 ) : ( n24808 ) ;
assign n24810 =  ( n24410 ) ? ( bv_8_53_n436 ) : ( n24809 ) ;
assign n24811 =  ( n24408 ) ? ( bv_8_136_n425 ) : ( n24810 ) ;
assign n24812 =  ( n24406 ) ? ( bv_8_46_n429 ) : ( n24811 ) ;
assign n24813 =  ( n24404 ) ? ( bv_8_147_n392 ) : ( n24812 ) ;
assign n24814 =  ( n24402 ) ? ( bv_8_85_n423 ) : ( n24813 ) ;
assign n24815 =  ( n24400 ) ? ( bv_8_252_n15 ) : ( n24814 ) ;
assign n24816 =  ( n24398 ) ? ( bv_8_122_n416 ) : ( n24815 ) ;
assign n24817 =  ( n24396 ) ? ( bv_8_200_n213 ) : ( n24816 ) ;
assign n24818 =  ( n24394 ) ? ( bv_8_186_n263 ) : ( n24817 ) ;
assign n24819 =  ( n24392 ) ? ( bv_8_50_n408 ) : ( n24818 ) ;
assign n24820 =  ( n24390 ) ? ( bv_8_230_n103 ) : ( n24819 ) ;
assign n24821 =  ( n24388 ) ? ( bv_8_192_n242 ) : ( n24820 ) ;
assign n24822 =  ( n24386 ) ? ( bv_8_25_n399 ) : ( n24821 ) ;
assign n24823 =  ( n24384 ) ? ( bv_8_158_n355 ) : ( n24822 ) ;
assign n24824 =  ( n24382 ) ? ( bv_8_163_n339 ) : ( n24823 ) ;
assign n24825 =  ( n24380 ) ? ( bv_8_68_n390 ) : ( n24824 ) ;
assign n24826 =  ( n24378 ) ? ( bv_8_84_n386 ) : ( n24825 ) ;
assign n24827 =  ( n24376 ) ? ( bv_8_59_n382 ) : ( n24826 ) ;
assign n24828 =  ( n24374 ) ? ( bv_8_11_n379 ) : ( n24827 ) ;
assign n24829 =  ( n24372 ) ? ( bv_8_140_n376 ) : ( n24828 ) ;
assign n24830 =  ( n24370 ) ? ( bv_8_199_n216 ) : ( n24829 ) ;
assign n24831 =  ( n24368 ) ? ( bv_8_107_n370 ) : ( n24830 ) ;
assign n24832 =  ( n24366 ) ? ( bv_8_40_n366 ) : ( n24831 ) ;
assign n24833 =  ( n24364 ) ? ( bv_8_167_n325 ) : ( n24832 ) ;
assign n24834 =  ( n24362 ) ? ( bv_8_188_n257 ) : ( n24833 ) ;
assign n24835 =  ( n24360 ) ? ( bv_8_22_n357 ) : ( n24834 ) ;
assign n24836 =  ( n24358 ) ? ( bv_8_173_n307 ) : ( n24835 ) ;
assign n24837 =  ( n24356 ) ? ( bv_8_219_n146 ) : ( n24836 ) ;
assign n24838 =  ( n24354 ) ? ( bv_8_100_n348 ) : ( n24837 ) ;
assign n24839 =  ( n24352 ) ? ( bv_8_116_n345 ) : ( n24838 ) ;
assign n24840 =  ( n24350 ) ? ( bv_8_20_n341 ) : ( n24839 ) ;
assign n24841 =  ( n24348 ) ? ( bv_8_146_n337 ) : ( n24840 ) ;
assign n24842 =  ( n24346 ) ? ( bv_8_12_n333 ) : ( n24841 ) ;
assign n24843 =  ( n24344 ) ? ( bv_8_72_n330 ) : ( n24842 ) ;
assign n24844 =  ( n24342 ) ? ( bv_8_184_n270 ) : ( n24843 ) ;
assign n24845 =  ( n24340 ) ? ( bv_8_159_n323 ) : ( n24844 ) ;
assign n24846 =  ( n24338 ) ? ( bv_8_189_n254 ) : ( n24845 ) ;
assign n24847 =  ( n24336 ) ? ( bv_8_67_n318 ) : ( n24846 ) ;
assign n24848 =  ( n24334 ) ? ( bv_8_196_n228 ) : ( n24847 ) ;
assign n24849 =  ( n24332 ) ? ( bv_8_57_n312 ) : ( n24848 ) ;
assign n24850 =  ( n24330 ) ? ( bv_8_49_n309 ) : ( n24849 ) ;
assign n24851 =  ( n24328 ) ? ( bv_8_211_n175 ) : ( n24850 ) ;
assign n24852 =  ( n24326 ) ? ( bv_8_242_n55 ) : ( n24851 ) ;
assign n24853 =  ( n24324 ) ? ( bv_8_213_n167 ) : ( n24852 ) ;
assign n24854 =  ( n24322 ) ? ( bv_8_139_n297 ) : ( n24853 ) ;
assign n24855 =  ( n24320 ) ? ( bv_8_110_n294 ) : ( n24854 ) ;
assign n24856 =  ( n24318 ) ? ( bv_8_218_n150 ) : ( n24855 ) ;
assign n24857 =  ( n24316 ) ? ( bv_8_1_n287 ) : ( n24856 ) ;
assign n24858 =  ( n24314 ) ? ( bv_8_177_n283 ) : ( n24857 ) ;
assign n24859 =  ( n24312 ) ? ( bv_8_156_n279 ) : ( n24858 ) ;
assign n24860 =  ( n24310 ) ? ( bv_8_73_n275 ) : ( n24859 ) ;
assign n24861 =  ( n24308 ) ? ( bv_8_216_n157 ) : ( n24860 ) ;
assign n24862 =  ( n24306 ) ? ( bv_8_172_n268 ) : ( n24861 ) ;
assign n24863 =  ( n24304 ) ? ( bv_8_243_n51 ) : ( n24862 ) ;
assign n24864 =  ( n24302 ) ? ( bv_8_207_n188 ) : ( n24863 ) ;
assign n24865 =  ( n24300 ) ? ( bv_8_202_n207 ) : ( n24864 ) ;
assign n24866 =  ( n24298 ) ? ( bv_8_244_n47 ) : ( n24865 ) ;
assign n24867 =  ( n24296 ) ? ( bv_8_71_n252 ) : ( n24866 ) ;
assign n24868 =  ( n24294 ) ? ( bv_8_16_n248 ) : ( n24867 ) ;
assign n24869 =  ( n24292 ) ? ( bv_8_111_n244 ) : ( n24868 ) ;
assign n24870 =  ( n24290 ) ? ( bv_8_240_n63 ) : ( n24869 ) ;
assign n24871 =  ( n24288 ) ? ( bv_8_74_n237 ) : ( n24870 ) ;
assign n24872 =  ( n24286 ) ? ( bv_8_92_n234 ) : ( n24871 ) ;
assign n24873 =  ( n24284 ) ? ( bv_8_56_n230 ) : ( n24872 ) ;
assign n24874 =  ( n24282 ) ? ( bv_8_87_n226 ) : ( n24873 ) ;
assign n24875 =  ( n24280 ) ? ( bv_8_115_n222 ) : ( n24874 ) ;
assign n24876 =  ( n24278 ) ? ( bv_8_151_n218 ) : ( n24875 ) ;
assign n24877 =  ( n24276 ) ? ( bv_8_203_n203 ) : ( n24876 ) ;
assign n24878 =  ( n24274 ) ? ( bv_8_161_n211 ) : ( n24877 ) ;
assign n24879 =  ( n24272 ) ? ( bv_8_232_n95 ) : ( n24878 ) ;
assign n24880 =  ( n24270 ) ? ( bv_8_62_n205 ) : ( n24879 ) ;
assign n24881 =  ( n24268 ) ? ( bv_8_150_n201 ) : ( n24880 ) ;
assign n24882 =  ( n24266 ) ? ( bv_8_97_n198 ) : ( n24881 ) ;
assign n24883 =  ( n24264 ) ? ( bv_8_13_n194 ) : ( n24882 ) ;
assign n24884 =  ( n24262 ) ? ( bv_8_15_n190 ) : ( n24883 ) ;
assign n24885 =  ( n24260 ) ? ( bv_8_224_n126 ) : ( n24884 ) ;
assign n24886 =  ( n24258 ) ? ( bv_8_124_n184 ) : ( n24885 ) ;
assign n24887 =  ( n24256 ) ? ( bv_8_113_n180 ) : ( n24886 ) ;
assign n24888 =  ( n24254 ) ? ( bv_8_204_n177 ) : ( n24887 ) ;
assign n24889 =  ( n24252 ) ? ( bv_8_144_n173 ) : ( n24888 ) ;
assign n24890 =  ( n24250 ) ? ( bv_8_6_n169 ) : ( n24889 ) ;
assign n24891 =  ( n24248 ) ? ( bv_8_247_n35 ) : ( n24890 ) ;
assign n24892 =  ( n24246 ) ? ( bv_8_28_n162 ) : ( n24891 ) ;
assign n24893 =  ( n24244 ) ? ( bv_8_194_n159 ) : ( n24892 ) ;
assign n24894 =  ( n24242 ) ? ( bv_8_106_n155 ) : ( n24893 ) ;
assign n24895 =  ( n24240 ) ? ( bv_8_174_n152 ) : ( n24894 ) ;
assign n24896 =  ( n24238 ) ? ( bv_8_105_n148 ) : ( n24895 ) ;
assign n24897 =  ( n24236 ) ? ( bv_8_23_n144 ) : ( n24896 ) ;
assign n24898 =  ( n24234 ) ? ( bv_8_153_n140 ) : ( n24897 ) ;
assign n24899 =  ( n24232 ) ? ( bv_8_58_n136 ) : ( n24898 ) ;
assign n24900 =  ( n24230 ) ? ( bv_8_39_n132 ) : ( n24899 ) ;
assign n24901 =  ( n24228 ) ? ( bv_8_217_n128 ) : ( n24900 ) ;
assign n24902 =  ( n24226 ) ? ( bv_8_235_n83 ) : ( n24901 ) ;
assign n24903 =  ( n24224 ) ? ( bv_8_43_n121 ) : ( n24902 ) ;
assign n24904 =  ( n24222 ) ? ( bv_8_34_n117 ) : ( n24903 ) ;
assign n24905 =  ( n24220 ) ? ( bv_8_210_n113 ) : ( n24904 ) ;
assign n24906 =  ( n24218 ) ? ( bv_8_169_n109 ) : ( n24905 ) ;
assign n24907 =  ( n24216 ) ? ( bv_8_7_n105 ) : ( n24906 ) ;
assign n24908 =  ( n24214 ) ? ( bv_8_51_n101 ) : ( n24907 ) ;
assign n24909 =  ( n24212 ) ? ( bv_8_45_n97 ) : ( n24908 ) ;
assign n24910 =  ( n24210 ) ? ( bv_8_60_n93 ) : ( n24909 ) ;
assign n24911 =  ( n24208 ) ? ( bv_8_21_n89 ) : ( n24910 ) ;
assign n24912 =  ( n24206 ) ? ( bv_8_201_n85 ) : ( n24911 ) ;
assign n24913 =  ( n24204 ) ? ( bv_8_135_n81 ) : ( n24912 ) ;
assign n24914 =  ( n24202 ) ? ( bv_8_170_n77 ) : ( n24913 ) ;
assign n24915 =  ( n24200 ) ? ( bv_8_80_n73 ) : ( n24914 ) ;
assign n24916 =  ( n24198 ) ? ( bv_8_165_n69 ) : ( n24915 ) ;
assign n24917 =  ( n24196 ) ? ( bv_8_3_n65 ) : ( n24916 ) ;
assign n24918 =  ( n24194 ) ? ( bv_8_89_n61 ) : ( n24917 ) ;
assign n24919 =  ( n24192 ) ? ( bv_8_9_n57 ) : ( n24918 ) ;
assign n24920 =  ( n24190 ) ? ( bv_8_26_n53 ) : ( n24919 ) ;
assign n24921 =  ( n24188 ) ? ( bv_8_101_n49 ) : ( n24920 ) ;
assign n24922 =  ( n24186 ) ? ( bv_8_215_n45 ) : ( n24921 ) ;
assign n24923 =  ( n24184 ) ? ( bv_8_132_n41 ) : ( n24922 ) ;
assign n24924 =  ( n24182 ) ? ( bv_8_208_n37 ) : ( n24923 ) ;
assign n24925 =  ( n24180 ) ? ( bv_8_130_n33 ) : ( n24924 ) ;
assign n24926 =  ( n24178 ) ? ( bv_8_41_n29 ) : ( n24925 ) ;
assign n24927 =  ( n24176 ) ? ( bv_8_90_n25 ) : ( n24926 ) ;
assign n24928 =  ( n24174 ) ? ( bv_8_30_n21 ) : ( n24927 ) ;
assign n24929 =  ( n24172 ) ? ( bv_8_123_n17 ) : ( n24928 ) ;
assign n24930 =  ( n24170 ) ? ( bv_8_168_n13 ) : ( n24929 ) ;
assign n24931 =  ( n24168 ) ? ( bv_8_109_n9 ) : ( n24930 ) ;
assign n24932 =  ( n24166 ) ? ( bv_8_44_n5 ) : ( n24931 ) ;
assign n24933 =  ( n24164 ) ^ ( n24932 )  ;
assign n24934 =  ( n24933 ) ^ ( n24158 )  ;
assign n24935 = key[15:8] ;
assign n24936 =  ( n24934 ) ^ ( n24935 )  ;
assign n24937 =  { ( n24162 ) , ( n24936 ) }  ;
assign n24938 =  ( n19540 ) ^ ( n21077 )  ;
assign n24939 =  ( n24938 ) ^ ( n24932 )  ;
assign n24940 =  ( n24939 ) ^ ( n24158 )  ;
assign n24941 =  ( n24940 ) ^ ( n22615 )  ;
assign n24942 = key[7:0] ;
assign n24943 =  ( n24941 ) ^ ( n24942 )  ;
assign n24944 =  { ( n24937 ) , ( n24943 ) }  ;
assign n24945 =  ( bv_128_0_n1 ) + ( n24944 )  ;
always @(posedge clk) begin
   if(rst) begin
       key <= key_randinit ;
       state_in <= state_in_randinit ;
       state_out <= state_out_randinit ;
       __COUNTER_start__n0 <= 0;
   end
   else if(__START__ && __ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           key <= key ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           state_in <= state_in ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           state_out <= n24945 ;
       end
   end
end
endmodule
