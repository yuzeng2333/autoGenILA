module NV_NVDLA_CDP_RDMA_cq_flopram_rwsa_32x7(clk, pwrbus_ram_pd, di, we, wa, ra, dout);
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _000_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _001_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _002_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _003_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _004_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _005_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _006_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _007_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _008_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _009_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _010_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _011_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _012_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _013_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _014_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _015_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _016_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _017_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _018_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _019_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _020_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _021_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _022_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _023_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _024_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _025_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _026_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _027_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _028_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _029_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _030_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:457" *)
  wire [6:0] _031_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:458" *)
  wire _032_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:461" *)
  wire _033_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:464" *)
  wire _034_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:467" *)
  wire _035_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:470" *)
  wire _036_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:473" *)
  wire _037_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:476" *)
  wire _038_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:479" *)
  wire _039_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:482" *)
  wire _040_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:485" *)
  wire _041_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:488" *)
  wire _042_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:491" *)
  wire _043_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:494" *)
  wire _044_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:497" *)
  wire _045_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:500" *)
  wire _046_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:503" *)
  wire _047_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:506" *)
  wire _048_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:509" *)
  wire _049_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:512" *)
  wire _050_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:515" *)
  wire _051_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:518" *)
  wire _052_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:521" *)
  wire _053_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:524" *)
  wire _054_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:527" *)
  wire _055_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:530" *)
  wire _056_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:533" *)
  wire _057_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:536" *)
  wire _058_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:539" *)
  wire _059_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:542" *)
  wire _060_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:545" *)
  wire _061_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:548" *)
  wire _062_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:551" *)
  wire _063_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:458" *)
  wire _064_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:461" *)
  wire _065_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:464" *)
  wire _066_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:467" *)
  wire _067_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:470" *)
  wire _068_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:473" *)
  wire _069_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:476" *)
  wire _070_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:479" *)
  wire _071_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:482" *)
  wire _072_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:485" *)
  wire _073_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:488" *)
  wire _074_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:491" *)
  wire _075_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:494" *)
  wire _076_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:497" *)
  wire _077_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:500" *)
  wire _078_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:503" *)
  wire _079_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:506" *)
  wire _080_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:509" *)
  wire _081_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:512" *)
  wire _082_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:515" *)
  wire _083_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:518" *)
  wire _084_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:521" *)
  wire _085_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:524" *)
  wire _086_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:527" *)
  wire _087_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:530" *)
  wire _088_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:533" *)
  wire _089_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:536" *)
  wire _090_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:539" *)
  wire _091_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:542" *)
  wire _092_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:545" *)
  wire _093_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:548" *)
  wire _094_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:551" *)
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:366" *)
  input clk;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:368" *)
  input [6:0] di;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:372" *)
  output [6:0] dout;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:367" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:371" *)
  input [4:0] ra;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:425" *)
  reg [6:0] ram_ff0;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:426" *)
  reg [6:0] ram_ff1;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:435" *)
  reg [6:0] ram_ff10;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:436" *)
  reg [6:0] ram_ff11;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:437" *)
  reg [6:0] ram_ff12;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:438" *)
  reg [6:0] ram_ff13;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:439" *)
  reg [6:0] ram_ff14;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:440" *)
  reg [6:0] ram_ff15;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:441" *)
  reg [6:0] ram_ff16;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:442" *)
  reg [6:0] ram_ff17;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:443" *)
  reg [6:0] ram_ff18;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:444" *)
  reg [6:0] ram_ff19;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:427" *)
  reg [6:0] ram_ff2;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:445" *)
  reg [6:0] ram_ff20;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:446" *)
  reg [6:0] ram_ff21;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:447" *)
  reg [6:0] ram_ff22;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:448" *)
  reg [6:0] ram_ff23;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:449" *)
  reg [6:0] ram_ff24;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:450" *)
  reg [6:0] ram_ff25;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:451" *)
  reg [6:0] ram_ff26;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:452" *)
  reg [6:0] ram_ff27;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:453" *)
  reg [6:0] ram_ff28;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:454" *)
  reg [6:0] ram_ff29;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:428" *)
  reg [6:0] ram_ff3;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:455" *)
  reg [6:0] ram_ff30;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:456" *)
  reg [6:0] ram_ff31;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:429" *)
  reg [6:0] ram_ff4;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:430" *)
  reg [6:0] ram_ff5;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:431" *)
  reg [6:0] ram_ff6;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:432" *)
  reg [6:0] ram_ff7;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:433" *)
  reg [6:0] ram_ff8;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:434" *)
  reg [6:0] ram_ff9;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:370" *)
  input [4:0] wa;
  (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:369" *)
  input we;
  assign _032_ = ! (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:458" *) wa;
  assign _033_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:461" *) 1'b1;
  assign _034_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:464" *) 2'b10;
  assign _035_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:467" *) 2'b11;
  assign _036_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:470" *) 3'b100;
  assign _037_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:473" *) 3'b101;
  assign _038_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:476" *) 3'b110;
  assign _039_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:479" *) 3'b111;
  assign _040_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:482" *) 4'b1000;
  assign _041_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:485" *) 4'b1001;
  assign _042_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:488" *) 4'b1010;
  assign _043_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:491" *) 4'b1011;
  assign _044_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:494" *) 4'b1100;
  assign _045_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:497" *) 4'b1101;
  assign _046_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:500" *) 4'b1110;
  assign _047_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:503" *) 4'b1111;
  assign _048_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:506" *) 5'b10000;
  assign _049_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:509" *) 5'b10001;
  assign _050_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:512" *) 5'b10010;
  assign _051_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:515" *) 5'b10011;
  assign _052_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:518" *) 5'b10100;
  assign _053_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:521" *) 5'b10101;
  assign _054_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:524" *) 5'b10110;
  assign _055_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:527" *) 5'b10111;
  assign _056_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:530" *) 5'b11000;
  assign _057_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:533" *) 5'b11001;
  assign _058_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:536" *) 5'b11010;
  assign _059_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:539" *) 5'b11011;
  assign _060_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:542" *) 5'b11100;
  assign _061_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:545" *) 5'b11101;
  assign _062_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:548" *) 5'b11110;
  assign _063_ = wa == (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:551" *) 5'b11111;
  assign _064_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:458" *) _032_;
  assign _065_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:461" *) _033_;
  assign _066_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:464" *) _034_;
  assign _067_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:467" *) _035_;
  assign _068_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:470" *) _036_;
  assign _069_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:473" *) _037_;
  assign _070_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:476" *) _038_;
  assign _071_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:479" *) _039_;
  assign _072_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:482" *) _040_;
  assign _073_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:485" *) _041_;
  assign _074_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:488" *) _042_;
  assign _075_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:491" *) _043_;
  assign _076_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:494" *) _044_;
  assign _077_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:497" *) _045_;
  assign _078_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:500" *) _046_;
  assign _079_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:503" *) _047_;
  assign _080_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:506" *) _048_;
  assign _081_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:509" *) _049_;
  assign _082_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:512" *) _050_;
  assign _083_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:515" *) _051_;
  assign _084_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:518" *) _052_;
  assign _085_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:521" *) _053_;
  assign _086_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:524" *) _054_;
  assign _087_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:527" *) _055_;
  assign _088_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:530" *) _056_;
  assign _089_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:533" *) _057_;
  assign _090_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:536" *) _058_;
  assign _091_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:539" *) _059_;
  assign _092_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:542" *) _060_;
  assign _093_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:545" *) _061_;
  assign _094_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:548" *) _062_;
  assign _095_ = we && (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:551" *) _063_;
  always @(posedge clk)
      ram_ff0 <= _000_;
  always @(posedge clk)
      ram_ff1 <= _011_;
  always @(posedge clk)
      ram_ff2 <= _022_;
  always @(posedge clk)
      ram_ff3 <= _025_;
  always @(posedge clk)
      ram_ff4 <= _026_;
  always @(posedge clk)
      ram_ff5 <= _027_;
  always @(posedge clk)
      ram_ff6 <= _028_;
  always @(posedge clk)
      ram_ff7 <= _029_;
  always @(posedge clk)
      ram_ff8 <= _030_;
  always @(posedge clk)
      ram_ff9 <= _031_;
  always @(posedge clk)
      ram_ff10 <= _001_;
  always @(posedge clk)
      ram_ff11 <= _002_;
  always @(posedge clk)
      ram_ff12 <= _003_;
  always @(posedge clk)
      ram_ff13 <= _004_;
  always @(posedge clk)
      ram_ff14 <= _005_;
  always @(posedge clk)
      ram_ff15 <= _006_;
  always @(posedge clk)
      ram_ff16 <= _007_;
  always @(posedge clk)
      ram_ff17 <= _008_;
  always @(posedge clk)
      ram_ff18 <= _009_;
  always @(posedge clk)
      ram_ff19 <= _010_;
  always @(posedge clk)
      ram_ff20 <= _012_;
  always @(posedge clk)
      ram_ff21 <= _013_;
  always @(posedge clk)
      ram_ff22 <= _014_;
  always @(posedge clk)
      ram_ff23 <= _015_;
  always @(posedge clk)
      ram_ff24 <= _016_;
  always @(posedge clk)
      ram_ff25 <= _017_;
  always @(posedge clk)
      ram_ff26 <= _018_;
  always @(posedge clk)
      ram_ff27 <= _019_;
  always @(posedge clk)
      ram_ff28 <= _020_;
  always @(posedge clk)
      ram_ff29 <= _021_;
  always @(posedge clk)
      ram_ff30 <= _023_;
  always @(posedge clk)
      ram_ff31 <= _024_;
  function [6:0] _223_;
    input [6:0] a;
    input [216:0] b;
    input [30:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:589|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *)
    (* parallel_case *)
    casez (s)
      31'b??????????????????????????????1:
        _223_ = b[6:0];
      31'b?????????????????????????????1?:
        _223_ = b[13:7];
      31'b????????????????????????????1??:
        _223_ = b[20:14];
      31'b???????????????????????????1???:
        _223_ = b[27:21];
      31'b??????????????????????????1????:
        _223_ = b[34:28];
      31'b?????????????????????????1?????:
        _223_ = b[41:35];
      31'b????????????????????????1??????:
        _223_ = b[48:42];
      31'b???????????????????????1???????:
        _223_ = b[55:49];
      31'b??????????????????????1????????:
        _223_ = b[62:56];
      31'b?????????????????????1?????????:
        _223_ = b[69:63];
      31'b????????????????????1??????????:
        _223_ = b[76:70];
      31'b???????????????????1???????????:
        _223_ = b[83:77];
      31'b??????????????????1????????????:
        _223_ = b[90:84];
      31'b?????????????????1?????????????:
        _223_ = b[97:91];
      31'b????????????????1??????????????:
        _223_ = b[104:98];
      31'b???????????????1???????????????:
        _223_ = b[111:105];
      31'b??????????????1????????????????:
        _223_ = b[118:112];
      31'b?????????????1?????????????????:
        _223_ = b[125:119];
      31'b????????????1??????????????????:
        _223_ = b[132:126];
      31'b???????????1???????????????????:
        _223_ = b[139:133];
      31'b??????????1????????????????????:
        _223_ = b[146:140];
      31'b?????????1?????????????????????:
        _223_ = b[153:147];
      31'b????????1??????????????????????:
        _223_ = b[160:154];
      31'b???????1???????????????????????:
        _223_ = b[167:161];
      31'b??????1????????????????????????:
        _223_ = b[174:168];
      31'b?????1?????????????????????????:
        _223_ = b[181:175];
      31'b????1??????????????????????????:
        _223_ = b[188:182];
      31'b???1???????????????????????????:
        _223_ = b[195:189];
      31'b??1????????????????????????????:
        _223_ = b[202:196];
      31'b?1?????????????????????????????:
        _223_ = b[209:203];
      31'b1??????????????????????????????:
        _223_ = b[216:210];
      default:
        _223_ = a;
    endcase
  endfunction
  assign dout = _223_(ram_ff0, { ram_ff1, ram_ff2, ram_ff3, ram_ff4, ram_ff5, ram_ff6, ram_ff7, ram_ff8, ram_ff9, ram_ff10, ram_ff11, ram_ff12, ram_ff13, ram_ff14, ram_ff15, ram_ff16, ram_ff17, ram_ff18, ram_ff19, ram_ff20, ram_ff21, ram_ff22, ram_ff23, ram_ff24, ram_ff25, ram_ff26, ram_ff27, ram_ff28, ram_ff29, ram_ff30, ram_ff31 }, { _126_, _125_, _124_, _123_, _122_, _121_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _110_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_, _099_, _098_, _097_, _096_ });
  assign _096_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:589|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11111;
  assign _097_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:588|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11110;
  assign _098_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:587|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11101;
  assign _099_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:586|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11100;
  assign _100_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:585|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11011;
  assign _101_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:584|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11010;
  assign _102_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:583|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11001;
  assign _103_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:582|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b11000;
  assign _104_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:581|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10111;
  assign _105_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:580|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10110;
  assign _106_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:579|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10101;
  assign _107_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:578|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10100;
  assign _108_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:577|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10011;
  assign _109_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:576|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10010;
  assign _110_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:575|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10001;
  assign _111_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:574|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 5'b10000;
  assign _112_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:573|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1111;
  assign _113_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:572|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1110;
  assign _114_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:571|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1101;
  assign _115_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:570|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1100;
  assign _116_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:569|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1011;
  assign _117_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:568|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1010;
  assign _118_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:567|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1001;
  assign _119_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:566|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 4'b1000;
  assign _120_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:565|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 3'b111;
  assign _121_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:564|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 3'b110;
  assign _122_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:563|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 3'b101;
  assign _123_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:562|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 3'b100;
  assign _124_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:561|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 2'b11;
  assign _125_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:560|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 2'b10;
  assign _126_ = ra == (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:559|./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:557" *) 1'b1;
  assign _024_ = _095_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:551" *) di : ram_ff31;
  assign _023_ = _094_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:548" *) di : ram_ff30;
  assign _021_ = _093_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:545" *) di : ram_ff29;
  assign _020_ = _092_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:542" *) di : ram_ff28;
  assign _019_ = _091_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:539" *) di : ram_ff27;
  assign _018_ = _090_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:536" *) di : ram_ff26;
  assign _017_ = _089_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:533" *) di : ram_ff25;
  assign _016_ = _088_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:530" *) di : ram_ff24;
  assign _015_ = _087_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:527" *) di : ram_ff23;
  assign _014_ = _086_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:524" *) di : ram_ff22;
  assign _013_ = _085_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:521" *) di : ram_ff21;
  assign _012_ = _084_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:518" *) di : ram_ff20;
  assign _010_ = _083_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:515" *) di : ram_ff19;
  assign _009_ = _082_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:512" *) di : ram_ff18;
  assign _008_ = _081_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:509" *) di : ram_ff17;
  assign _007_ = _080_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:506" *) di : ram_ff16;
  assign _006_ = _079_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:503" *) di : ram_ff15;
  assign _005_ = _078_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:500" *) di : ram_ff14;
  assign _004_ = _077_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:497" *) di : ram_ff13;
  assign _003_ = _076_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:494" *) di : ram_ff12;
  assign _002_ = _075_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:491" *) di : ram_ff11;
  assign _001_ = _074_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:488" *) di : ram_ff10;
  assign _031_ = _073_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:485" *) di : ram_ff9;
  assign _030_ = _072_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:482" *) di : ram_ff8;
  assign _029_ = _071_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:479" *) di : ram_ff7;
  assign _028_ = _070_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:476" *) di : ram_ff6;
  assign _027_ = _069_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:473" *) di : ram_ff5;
  assign _026_ = _068_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:470" *) di : ram_ff4;
  assign _025_ = _067_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:467" *) di : ram_ff3;
  assign _022_ = _066_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:464" *) di : ram_ff2;
  assign _011_ = _065_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:461" *) di : ram_ff1;
  assign _000_ = _064_ ? (* src = "./vmod/nvdla/cdp/NV_NVDLA_CDP_RDMA_cq.v:458" *) di : ram_ff0;
endmodule
