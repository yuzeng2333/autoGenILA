module \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=5\width=8 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:78" *)
  output [7:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:79" *)
  input [7:0] z;
  assign d = z;
endmodule
