module NV_NVDLA_SDP_MRDMA_EG_dout(nvdla_core_clk, nvdla_core_rstn, cmd2dat_dma_pd, cmd2dat_dma_pvld, op_load, pfifo0_rd_pd, pfifo0_rd_pvld, pfifo1_rd_pd, pfifo1_rd_pvld, pfifo2_rd_pd, pfifo2_rd_pvld, pfifo3_rd_pd, pfifo3_rd_pvld, reg2dp_height, reg2dp_in_precision, reg2dp_perf_nan_inf_count_en, reg2dp_proc_precision, reg2dp_width, sdp_mrdma2cmux_ready, sfifo0_rd_pd, sfifo0_rd_pvld, sfifo1_rd_pd, sfifo1_rd_pvld, cmd2dat_dma_prdy, dp2reg_status_inf_input_num, dp2reg_status_nan_input_num, eg_done, pfifo0_rd_prdy, pfifo1_rd_prdy, pfifo2_rd_prdy, pfifo3_rd_prdy, sdp_mrdma2cmux_pd, sdp_mrdma2cmux_valid, sfifo0_rd_prdy, sfifo1_rd_prdy);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0102_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0103_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0104_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0105_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0106_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0107_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0108_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0109_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0110_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0111_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0112_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0113_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire _0127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:587" *)
  wire [13:0] _0128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1181" *)
  wire _0129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:639" *)
  wire [31:0] _0130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:693" *)
  wire [31:0] _0131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [7:0] _0322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1417" *)
  wire [22:0] _0323_;
  wire [4:0] _0324_;
  wire [4:0] _0325_;
  wire [4:0] _0326_;
  wire [4:0] _0327_;
  wire [4:0] _0328_;
  wire [4:0] _0329_;
  wire [4:0] _0330_;
  wire [4:0] _0331_;
  wire [4:0] _0332_;
  wire [4:0] _0333_;
  wire [4:0] _0334_;
  wire [4:0] _0335_;
  wire [4:0] _0336_;
  wire [4:0] _0337_;
  wire [4:0] _0338_;
  wire [4:0] _0339_;
  wire [4:0] _0340_;
  wire [4:0] _0341_;
  wire [4:0] _0342_;
  wire [4:0] _0343_;
  wire [4:0] _0344_;
  wire [4:0] _0345_;
  wire [4:0] _0346_;
  wire [4:0] _0347_;
  wire [4:0] _0348_;
  wire [4:0] _0349_;
  wire [4:0] _0350_;
  wire [4:0] _0351_;
  wire [4:0] _0352_;
  wire [4:0] _0353_;
  wire [4:0] _0354_;
  wire [4:0] _0355_;
  wire [7:0] _0356_;
  wire [7:0] _0357_;
  wire [7:0] _0358_;
  wire [7:0] _0359_;
  wire [7:0] _0360_;
  wire [7:0] _0361_;
  wire [7:0] _0362_;
  wire [7:0] _0363_;
  wire [7:0] _0364_;
  wire [7:0] _0365_;
  wire [7:0] _0366_;
  wire [7:0] _0367_;
  wire [7:0] _0368_;
  wire [7:0] _0369_;
  wire [7:0] _0370_;
  wire [7:0] _0371_;
  wire [7:0] _0372_;
  wire [7:0] _0373_;
  wire [7:0] _0374_;
  wire [7:0] _0375_;
  wire [7:0] _0376_;
  wire [7:0] _0377_;
  wire [7:0] _0378_;
  wire [7:0] _0379_;
  wire [7:0] _0380_;
  wire [7:0] _0381_;
  wire [7:0] _0382_;
  wire [7:0] _0383_;
  wire [7:0] _0384_;
  wire [7:0] _0385_;
  wire [7:0] _0386_;
  wire [7:0] _0387_;
  wire [1:0] _0388_;
  wire [1:0] _0389_;
  wire [1:0] _0390_;
  wire [1:0] _0391_;
  wire [1:0] _0392_;
  wire [1:0] _0393_;
  wire [1:0] _0394_;
  wire [1:0] _0395_;
  wire [1:0] _0396_;
  wire [1:0] _0397_;
  wire [1:0] _0398_;
  wire [1:0] _0399_;
  wire [1:0] _0400_;
  wire [1:0] _0401_;
  wire [1:0] _0402_;
  wire [1:0] _0403_;
  wire [1:0] _0404_;
  wire [1:0] _0405_;
  wire [1:0] _0406_;
  wire [1:0] _0407_;
  wire [1:0] _0408_;
  wire [1:0] _0409_;
  wire [1:0] _0410_;
  wire [1:0] _0411_;
  wire [1:0] _0412_;
  wire [1:0] _0413_;
  wire [1:0] _0414_;
  wire [1:0] _0415_;
  wire [1:0] _0416_;
  wire [1:0] _0417_;
  wire [1:0] _0418_;
  wire [1:0] _0419_;
  wire [2:0] _0420_;
  wire [2:0] _0421_;
  wire [2:0] _0422_;
  wire [2:0] _0423_;
  wire [2:0] _0424_;
  wire [2:0] _0425_;
  wire [2:0] _0426_;
  wire [2:0] _0427_;
  wire [2:0] _0428_;
  wire [2:0] _0429_;
  wire [2:0] _0430_;
  wire [2:0] _0431_;
  wire [2:0] _0432_;
  wire [2:0] _0433_;
  wire [2:0] _0434_;
  wire [2:0] _0435_;
  wire [2:0] _0436_;
  wire [2:0] _0437_;
  wire [2:0] _0438_;
  wire [2:0] _0439_;
  wire [2:0] _0440_;
  wire [2:0] _0441_;
  wire [2:0] _0442_;
  wire [2:0] _0443_;
  wire [2:0] _0444_;
  wire [2:0] _0445_;
  wire [2:0] _0446_;
  wire [2:0] _0447_;
  wire [2:0] _0448_;
  wire [2:0] _0449_;
  wire [2:0] _0450_;
  wire [2:0] _0451_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0452_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0453_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0454_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0455_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0456_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0457_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0458_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0459_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0460_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0461_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0462_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0463_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0464_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0465_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0466_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0467_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0468_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0469_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0470_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0471_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0472_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0473_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0474_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0475_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0476_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0477_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0478_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0479_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0480_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0481_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0482_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *)
  wire [3:0] _0483_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0484_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0485_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0486_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0487_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0488_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0489_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0490_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0491_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0492_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0493_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0494_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0495_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0496_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0497_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0498_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0499_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0500_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0501_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0502_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0503_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0504_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0505_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0506_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0507_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0508_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0509_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0510_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0511_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0512_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0513_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0514_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *)
  wire [3:0] _0515_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0516_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0517_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0518_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0519_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0520_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0521_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0522_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0523_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0524_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0525_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0526_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0527_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0528_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0529_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0530_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0531_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0532_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0533_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0534_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0535_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0536_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0537_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0538_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0539_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0540_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0541_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0542_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0543_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0544_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0545_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0546_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *)
  wire [3:0] _0547_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0548_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0549_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0550_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0551_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0552_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0553_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0554_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0555_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0556_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0557_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0558_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0559_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0560_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0561_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0562_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0563_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0564_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0565_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0566_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0567_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0568_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0569_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0570_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0571_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0572_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0573_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0574_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0575_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0576_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0577_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0578_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *)
  wire [3:0] _0579_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0580_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0581_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0582_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0583_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0584_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0585_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0586_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0587_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0588_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0589_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0590_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0591_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0592_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0593_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0594_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0595_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0596_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0597_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0598_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0599_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0600_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0601_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0602_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0603_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0604_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0605_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0606_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0607_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0608_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0609_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0610_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *)
  wire [3:0] _0611_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0612_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0613_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0614_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0615_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0616_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0617_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0618_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0619_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0620_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0621_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0622_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0623_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0624_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0625_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0626_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0627_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0628_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0629_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0630_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0631_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0632_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0633_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0634_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0635_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0636_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0637_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0638_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0639_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0640_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0641_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0642_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *)
  wire [3:0] _0643_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0644_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0645_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0646_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0647_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0648_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0649_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0650_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0651_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0652_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0653_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0654_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0655_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0656_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0657_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0658_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0659_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0660_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0661_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0662_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0663_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0664_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0665_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0666_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0667_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0668_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0669_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0670_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0671_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0672_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0673_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0674_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *)
  wire [3:0] _0675_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0676_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0677_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0678_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0679_;
  wire _0680_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0681_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0682_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0683_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0684_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0685_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0686_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0687_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0688_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0689_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0690_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0691_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0692_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0693_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0694_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0695_;
  wire _0696_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0697_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0698_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0699_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0700_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0701_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0702_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0703_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0704_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0705_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0706_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0707_;
  wire [13:0] _0708_;
  wire [1:0] _0709_;
  wire [2:0] _0710_;
  wire [3:0] _0711_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0712_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0713_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0714_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0715_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0716_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0717_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0718_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0719_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0720_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0721_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *)
  wire [4:0] _0722_;
  wire [1:0] _0723_;
  wire [2:0] _0724_;
  wire [3:0] _0725_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0726_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0727_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0728_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0729_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0730_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0731_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0732_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0733_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0734_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0735_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *)
  wire [4:0] _0736_;
  wire [1:0] _0737_;
  wire [2:0] _0738_;
  wire [3:0] _0739_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0740_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0741_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0742_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0743_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0744_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0745_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0746_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0747_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0748_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0749_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *)
  wire [4:0] _0750_;
  wire [1:0] _0751_;
  wire [2:0] _0752_;
  wire [3:0] _0753_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0754_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0755_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0756_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0757_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0758_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0759_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0760_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0761_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0762_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0763_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *)
  wire [4:0] _0764_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1185" *)
  wire _0765_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:580" *)
  wire _0766_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:580" *)
  wire _0767_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *)
  wire _0768_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *)
  wire _0769_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *)
  wire _0770_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *)
  wire _0771_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:738" *)
  wire _0772_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:738" *)
  wire _0773_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:742" *)
  wire _0774_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:743" *)
  wire _0775_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:744" *)
  wire _0776_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:745" *)
  wire _0777_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:746" *)
  wire _0778_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:747" *)
  wire _0779_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0780_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *)
  wire [3:0] _0781_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0782_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0783_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0784_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0785_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0786_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0787_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0788_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0789_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0790_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0791_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0792_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0793_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0794_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0795_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0796_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0797_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0798_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0799_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0800_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0801_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0802_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0803_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0804_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0805_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0806_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0807_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0808_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0809_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0810_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0811_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0812_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *)
  wire [10:0] _0813_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0814_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0815_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0816_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0817_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0818_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0819_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0820_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0821_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0822_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0823_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0824_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0825_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0826_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0827_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0828_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0829_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0830_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0831_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0832_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0833_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0834_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0835_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0836_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0837_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0838_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0839_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0840_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0841_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0842_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _0843_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0844_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0845_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0846_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0847_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0848_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0849_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0850_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0851_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0852_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0853_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0854_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0855_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0856_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0857_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0858_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0859_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0860_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0861_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0862_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0863_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0864_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0865_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0866_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _0867_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0868_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0869_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0870_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0871_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0872_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0873_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0874_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0875_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0876_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0877_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0878_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0879_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0880_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0881_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0882_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0883_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0884_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0885_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0886_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0887_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0888_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0889_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0890_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0891_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0892_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0893_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0894_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0895_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0896_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0897_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0898_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0899_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0900_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0901_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0902_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0903_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0904_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0905_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0906_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0907_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0908_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0909_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0910_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0911_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0912_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0913_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0914_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0915_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0916_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0917_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0918_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0919_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0920_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0921_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0922_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0923_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0924_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0925_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0926_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0927_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0928_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0929_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0930_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _0931_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0932_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0933_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0934_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0935_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0936_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0937_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0938_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0939_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0940_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0941_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0942_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0943_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0944_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0945_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0946_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0947_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0948_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0949_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0950_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0951_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0952_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0953_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0954_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0955_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0956_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0957_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0958_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0959_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0960_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0961_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0962_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *)
  wire _0963_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0964_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0965_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0966_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0967_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0968_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0969_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0970_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0971_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0972_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0973_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0974_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0975_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0976_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0977_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0978_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0979_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0980_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0981_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0982_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0983_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0984_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0985_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0986_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0987_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0988_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0989_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0990_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0991_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0992_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0993_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0994_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *)
  wire _0995_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:578" *)
  wire _0996_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:578" *)
  wire _0997_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:603" *)
  wire _0998_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:603" *)
  wire _0999_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:604" *)
  wire _1000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:604" *)
  wire _1001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:605" *)
  wire _1002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:605" *)
  wire _1003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:606" *)
  wire _1004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:606" *)
  wire _1005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:607" *)
  wire _1006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:607" *)
  wire _1007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:608" *)
  wire _1008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:608" *)
  wire _1009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:609" *)
  wire _1010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:609" *)
  wire _1011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:610" *)
  wire _1012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:610" *)
  wire _1013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:611" *)
  wire _1014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:611" *)
  wire _1015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:612" *)
  wire _1016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:612" *)
  wire _1017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:613" *)
  wire _1018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:613" *)
  wire _1019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:614" *)
  wire _1020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:614" *)
  wire _1021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:615" *)
  wire _1022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:615" *)
  wire _1023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:616" *)
  wire _1024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:616" *)
  wire _1025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:617" *)
  wire _1026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:617" *)
  wire _1027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:618" *)
  wire _1028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:618" *)
  wire _1029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:619" *)
  wire _1030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:619" *)
  wire _1031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:620" *)
  wire _1032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:620" *)
  wire _1033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:621" *)
  wire _1034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:621" *)
  wire _1035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:622" *)
  wire _1036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:622" *)
  wire _1037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:623" *)
  wire _1038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:623" *)
  wire _1039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:624" *)
  wire _1040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:624" *)
  wire _1041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:625" *)
  wire _1042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:625" *)
  wire _1043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:626" *)
  wire _1044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:626" *)
  wire _1045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:627" *)
  wire _1046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:627" *)
  wire _1047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:628" *)
  wire _1048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:628" *)
  wire _1049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:629" *)
  wire _1050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:629" *)
  wire _1051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:630" *)
  wire _1052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:630" *)
  wire _1053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:631" *)
  wire _1054_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:631" *)
  wire _1055_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:632" *)
  wire _1056_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:632" *)
  wire _1057_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:633" *)
  wire _1058_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:633" *)
  wire _1059_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:634" *)
  wire _1060_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:634" *)
  wire _1061_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:643" *)
  wire _1062_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:730" *)
  wire _1063_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:730" *)
  wire _1064_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:647" *)
  wire _1065_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:701" *)
  wire _1066_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:657" *)
  wire _1067_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:658" *)
  wire _1068_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:659" *)
  wire _1069_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:660" *)
  wire _1070_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:661" *)
  wire _1071_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:662" *)
  wire _1072_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:663" *)
  wire _1073_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:664" *)
  wire _1074_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:665" *)
  wire _1075_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:666" *)
  wire _1076_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:667" *)
  wire _1077_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:668" *)
  wire _1078_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:669" *)
  wire _1079_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:670" *)
  wire _1080_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:671" *)
  wire _1081_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:672" *)
  wire _1082_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:673" *)
  wire _1083_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:674" *)
  wire _1084_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:675" *)
  wire _1085_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:676" *)
  wire _1086_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:677" *)
  wire _1087_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:678" *)
  wire _1088_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:679" *)
  wire _1089_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:680" *)
  wire _1090_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:681" *)
  wire _1091_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:682" *)
  wire _1092_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:683" *)
  wire _1093_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:684" *)
  wire _1094_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:685" *)
  wire _1095_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:686" *)
  wire _1096_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:687" *)
  wire _1097_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:688" *)
  wire _1098_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1156" *)
  wire _1099_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1156" *)
  wire _1100_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *)
  wire _1101_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *)
  wire _1102_;
  wire [511:0] _1103_;
  wire [511:0] _1104_;
  wire [511:0] _1105_;
  wire [511:0] _1106_;
  wire [511:0] _1107_;
  wire [31:0] _1108_;
  wire [31:0] _1109_;
  wire [31:0] _1110_;
  wire [31:0] _1111_;
  wire [31:0] _1112_;
  wire [31:0] _1113_;
  wire [13:0] _1114_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:647" *)
  wire _1115_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:701" *)
  wire _1116_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1117_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1118_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1119_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1120_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1121_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1122_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1123_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1124_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1125_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1126_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1127_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1128_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1129_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1130_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1131_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1132_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1133_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1134_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1135_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1136_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1137_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1138_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1139_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1140_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1141_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1142_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1143_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1144_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1145_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1146_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1147_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *)
  wire _1148_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1149_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1150_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1151_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1152_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1153_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1154_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1155_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1156_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1157_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1158_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1159_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1160_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1161_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1162_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1163_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1164_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1165_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1166_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1167_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1168_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1169_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1170_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1171_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1172_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1173_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1174_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1175_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1176_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1177_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1178_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1179_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *)
  wire _1180_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1181_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1182_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1183_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1184_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1185_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1186_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1187_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1188_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1189_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1190_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1191_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1192_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1193_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1194_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1195_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1196_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1197_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1198_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1199_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1200_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1201_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1202_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1203_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1204_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1205_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1206_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1207_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1208_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1209_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1210_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1211_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *)
  wire _1212_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1213_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1214_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1215_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1216_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1217_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1218_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1219_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1220_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1221_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1222_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1223_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1224_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1225_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1226_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1227_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1228_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1229_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1230_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1231_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1232_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1233_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1234_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1235_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1236_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1237_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1238_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1239_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1240_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1241_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1242_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1243_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *)
  wire _1244_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1245_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1246_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1247_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1248_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1249_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1250_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1251_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1252_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1253_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1254_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1255_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1256_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1257_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1258_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1259_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1260_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1261_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1262_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1263_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1264_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1265_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1266_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1267_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1268_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1269_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1270_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1271_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1272_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1273_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1274_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1275_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *)
  wire _1276_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1277_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1278_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1279_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1280_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1281_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1282_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1283_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1284_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1285_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1286_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1287_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1288_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1289_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1290_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1291_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1292_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1293_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1294_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1295_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1296_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1297_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1298_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1299_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1300_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1301_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1302_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1303_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1304_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1305_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1306_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1307_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *)
  wire _1308_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1309_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1310_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1311_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1312_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1313_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1314_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1315_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1316_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1317_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1318_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1319_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1320_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1321_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1322_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1323_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1324_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1325_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1326_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1327_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1328_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1329_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1330_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1331_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1332_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1333_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1334_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1335_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1336_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1337_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1338_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1339_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *)
  wire _1340_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1341_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1342_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1343_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1344_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1345_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1346_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1347_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1348_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1349_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1350_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1351_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1352_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1353_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1354_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1355_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1356_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1357_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1358_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1359_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1360_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1361_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1362_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1363_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1364_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1365_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1366_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1367_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1368_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1369_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1370_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1371_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *)
  wire _1372_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1373_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1374_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1375_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1376_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1377_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1378_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1379_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1380_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1381_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1382_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1383_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1384_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1385_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1386_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1387_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1388_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1389_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1390_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1391_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1392_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1393_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1394_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1395_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1396_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1397_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1398_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1399_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1400_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1401_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1402_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1403_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *)
  wire _1404_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _1405_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *)
  (* unused_bits = "23" *)
  wire [23:0] _1406_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1407_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1408_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1409_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1410_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1411_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1412_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1413_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *)
  (* unused_bits = "8 9 10 11 12 13 14 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31" *)
  wire [31:0] _1414_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1158" *)
  wire [511:0] _1415_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:86" *)
  reg [13:0] beat_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:93" *)
  wire cfg_di_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:94" *)
  wire cfg_di_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:95" *)
  wire cfg_di_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:96" *)
  wire cfg_di_int8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:97" *)
  wire cfg_do_int8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:98" *)
  wire cfg_mode_16to8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:99" *)
  wire cfg_mode_1x1_pack;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:100" *)
  wire cfg_perf_nan_inf_count_en;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:101" *)
  wire cmd2dat_dma_cube_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:54" *)
  input [14:0] cmd2dat_dma_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:53" *)
  output cmd2dat_dma_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:52" *)
  input cmd2dat_dma_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:102" *)
  wire [13:0] cmd2dat_dma_size;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:103" *)
  wire cmd_cube_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:104" *)
  wire dat_accept;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:105" *)
  wire dat_batch_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:106" *)
  wire [511:0] dat_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:107" *)
  wire dat_layer_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:108" *)
  wire [513:0] dat_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:109" *)
  wire dat_rdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:110" *)
  wire dat_vld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:83" *)
  output [31:0] dp2reg_status_inf_input_num;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:84" *)
  output [31:0] dp2reg_status_nan_input_num;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:77" *)
  output eg_done;
  reg eg_done;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:111" *)
  wire fifo_vld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:88" *)
  reg [31:0] inf_input_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:112" *)
  wire [31:0] inf_input_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:113" *)
  wire inf_input_cnt_nxt_c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:114" *)
  wire is_last_beat;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:115" *)
  wire mode_16to8_pfifo0_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:116" *)
  wire mode_16to8_pfifo1_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:117" *)
  wire mode_16to8_pfifo2_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:118" *)
  wire mode_16to8_pfifo3_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:119" *)
  wire mode_16to8_sfifo0_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:120" *)
  wire mode_16to8_sfifo1_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:121" *)
  wire mode_norm_pfifo0_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:122" *)
  wire mode_norm_pfifo0_sel_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:123" *)
  wire mode_norm_pfifo0_sel_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:124" *)
  wire mode_norm_pfifo1_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:125" *)
  wire mode_norm_pfifo1_sel_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:126" *)
  wire mode_norm_pfifo1_sel_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:127" *)
  wire mode_norm_pfifo2_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:128" *)
  wire mode_norm_pfifo2_sel_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:129" *)
  wire mode_norm_pfifo2_sel_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:130" *)
  wire mode_norm_pfifo3_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:131" *)
  wire mode_norm_pfifo3_sel_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:132" *)
  wire mode_norm_pfifo3_sel_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:89" *)
  reg [31:0] nan_input_cnt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:133" *)
  wire [31:0] nan_input_cnt_nxt;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:134" *)
  wire nan_input_cnt_nxt_c;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:50" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:51" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:76" *)
  input op_load;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:135" *)
  wire [255:0] pfifo0_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:136" *)
  wire [15:0] pfifo0_data_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:137" *)
  wire [7:0] pfifo0_data_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:138" *)
  wire pfifo0_data_byte0_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:139" *)
  wire pfifo0_data_byte0_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:140" *)
  wire [7:0] pfifo0_data_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:141" *)
  wire [7:0] pfifo0_data_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:142" *)
  wire [7:0] pfifo0_data_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:143" *)
  wire [7:0] pfifo0_data_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:144" *)
  wire [7:0] pfifo0_data_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:145" *)
  wire [7:0] pfifo0_data_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:146" *)
  wire [15:0] pfifo0_data_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:147" *)
  wire [7:0] pfifo0_data_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:148" *)
  wire pfifo0_data_byte1_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:149" *)
  wire pfifo0_data_byte1_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:150" *)
  wire [15:0] pfifo0_data_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:151" *)
  wire [7:0] pfifo0_data_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:152" *)
  wire pfifo0_data_byte2_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:153" *)
  wire pfifo0_data_byte2_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:154" *)
  wire [15:0] pfifo0_data_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:155" *)
  wire [7:0] pfifo0_data_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:156" *)
  wire pfifo0_data_byte3_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:157" *)
  wire pfifo0_data_byte3_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:158" *)
  wire [15:0] pfifo0_data_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:159" *)
  wire [7:0] pfifo0_data_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:160" *)
  wire pfifo0_data_byte4_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:161" *)
  wire pfifo0_data_byte4_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:162" *)
  wire [15:0] pfifo0_data_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:163" *)
  wire [7:0] pfifo0_data_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:164" *)
  wire pfifo0_data_byte5_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:165" *)
  wire pfifo0_data_byte5_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:166" *)
  wire [15:0] pfifo0_data_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:167" *)
  wire [7:0] pfifo0_data_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:168" *)
  wire pfifo0_data_byte6_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:169" *)
  wire pfifo0_data_byte6_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:170" *)
  wire [15:0] pfifo0_data_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:171" *)
  wire [7:0] pfifo0_data_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:172" *)
  wire pfifo0_data_byte7_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:173" *)
  wire pfifo0_data_byte7_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:174" *)
  wire [7:0] pfifo0_data_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:175" *)
  wire [7:0] pfifo0_data_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:176" *)
  wire [31:0] pfifo0_data_ext_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:177" *)
  wire [31:0] pfifo0_data_ext_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:178" *)
  wire [31:0] pfifo0_data_ext_byte0_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:179" *)
  wire [31:0] pfifo0_data_ext_byte0_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:180" *)
  wire [31:0] pfifo0_data_ext_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:181" *)
  wire [31:0] pfifo0_data_ext_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:182" *)
  wire [31:0] pfifo0_data_ext_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:183" *)
  wire [31:0] pfifo0_data_ext_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:184" *)
  wire [31:0] pfifo0_data_ext_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:185" *)
  wire [31:0] pfifo0_data_ext_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:186" *)
  wire [31:0] pfifo0_data_ext_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:187" *)
  wire [31:0] pfifo0_data_ext_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:188" *)
  wire [31:0] pfifo0_data_ext_byte1_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:189" *)
  wire [31:0] pfifo0_data_ext_byte1_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:190" *)
  wire [31:0] pfifo0_data_ext_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:191" *)
  wire [31:0] pfifo0_data_ext_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:192" *)
  wire [31:0] pfifo0_data_ext_byte2_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:193" *)
  wire [31:0] pfifo0_data_ext_byte2_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:194" *)
  wire [31:0] pfifo0_data_ext_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:195" *)
  wire [31:0] pfifo0_data_ext_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:196" *)
  wire [31:0] pfifo0_data_ext_byte3_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:197" *)
  wire [31:0] pfifo0_data_ext_byte3_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:198" *)
  wire [31:0] pfifo0_data_ext_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:199" *)
  wire [31:0] pfifo0_data_ext_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:200" *)
  wire [31:0] pfifo0_data_ext_byte4_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:201" *)
  wire [31:0] pfifo0_data_ext_byte4_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:202" *)
  wire [31:0] pfifo0_data_ext_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:203" *)
  wire [31:0] pfifo0_data_ext_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:204" *)
  wire [31:0] pfifo0_data_ext_byte5_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:205" *)
  wire [31:0] pfifo0_data_ext_byte5_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:206" *)
  wire [31:0] pfifo0_data_ext_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:207" *)
  wire [31:0] pfifo0_data_ext_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:208" *)
  wire [31:0] pfifo0_data_ext_byte6_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:209" *)
  wire [31:0] pfifo0_data_ext_byte6_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:210" *)
  wire [31:0] pfifo0_data_ext_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:211" *)
  wire [31:0] pfifo0_data_ext_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:212" *)
  wire [31:0] pfifo0_data_ext_byte7_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:213" *)
  wire [31:0] pfifo0_data_ext_byte7_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:214" *)
  wire [31:0] pfifo0_data_ext_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:215" *)
  wire [31:0] pfifo0_data_ext_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:216" *)
  wire [127:0] pfifo0_rd_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:57" *)
  input [127:0] pfifo0_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:56" *)
  output pfifo0_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:55" *)
  input pfifo0_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:217" *)
  wire pfifo0_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:218" *)
  wire [255:0] pfifo1_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:219" *)
  wire [15:0] pfifo1_data_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:220" *)
  wire [7:0] pfifo1_data_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:221" *)
  wire pfifo1_data_byte0_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:222" *)
  wire pfifo1_data_byte0_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:223" *)
  wire [7:0] pfifo1_data_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:224" *)
  wire [7:0] pfifo1_data_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:225" *)
  wire [7:0] pfifo1_data_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:226" *)
  wire [7:0] pfifo1_data_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:227" *)
  wire [7:0] pfifo1_data_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:228" *)
  wire [7:0] pfifo1_data_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:229" *)
  wire [15:0] pfifo1_data_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:230" *)
  wire [7:0] pfifo1_data_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:231" *)
  wire pfifo1_data_byte1_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:232" *)
  wire pfifo1_data_byte1_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:233" *)
  wire [15:0] pfifo1_data_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:234" *)
  wire [7:0] pfifo1_data_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:235" *)
  wire pfifo1_data_byte2_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:236" *)
  wire pfifo1_data_byte2_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:237" *)
  wire [15:0] pfifo1_data_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:238" *)
  wire [7:0] pfifo1_data_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:239" *)
  wire pfifo1_data_byte3_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:240" *)
  wire pfifo1_data_byte3_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:241" *)
  wire [15:0] pfifo1_data_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:242" *)
  wire [7:0] pfifo1_data_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:243" *)
  wire pfifo1_data_byte4_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:244" *)
  wire pfifo1_data_byte4_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:245" *)
  wire [15:0] pfifo1_data_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:246" *)
  wire [7:0] pfifo1_data_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:247" *)
  wire pfifo1_data_byte5_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:248" *)
  wire pfifo1_data_byte5_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:249" *)
  wire [15:0] pfifo1_data_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:250" *)
  wire [7:0] pfifo1_data_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:251" *)
  wire pfifo1_data_byte6_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:252" *)
  wire pfifo1_data_byte6_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:253" *)
  wire [15:0] pfifo1_data_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:254" *)
  wire [7:0] pfifo1_data_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:255" *)
  wire pfifo1_data_byte7_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:256" *)
  wire pfifo1_data_byte7_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:257" *)
  wire [7:0] pfifo1_data_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:258" *)
  wire [7:0] pfifo1_data_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:259" *)
  wire [31:0] pfifo1_data_ext_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:260" *)
  wire [31:0] pfifo1_data_ext_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:261" *)
  wire [31:0] pfifo1_data_ext_byte0_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:262" *)
  wire [31:0] pfifo1_data_ext_byte0_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:263" *)
  wire [31:0] pfifo1_data_ext_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:264" *)
  wire [31:0] pfifo1_data_ext_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:265" *)
  wire [31:0] pfifo1_data_ext_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:266" *)
  wire [31:0] pfifo1_data_ext_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:267" *)
  wire [31:0] pfifo1_data_ext_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:268" *)
  wire [31:0] pfifo1_data_ext_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:269" *)
  wire [31:0] pfifo1_data_ext_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:270" *)
  wire [31:0] pfifo1_data_ext_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:271" *)
  wire [31:0] pfifo1_data_ext_byte1_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:272" *)
  wire [31:0] pfifo1_data_ext_byte1_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:273" *)
  wire [31:0] pfifo1_data_ext_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:274" *)
  wire [31:0] pfifo1_data_ext_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:275" *)
  wire [31:0] pfifo1_data_ext_byte2_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:276" *)
  wire [31:0] pfifo1_data_ext_byte2_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:277" *)
  wire [31:0] pfifo1_data_ext_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:278" *)
  wire [31:0] pfifo1_data_ext_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:279" *)
  wire [31:0] pfifo1_data_ext_byte3_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:280" *)
  wire [31:0] pfifo1_data_ext_byte3_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:281" *)
  wire [31:0] pfifo1_data_ext_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:282" *)
  wire [31:0] pfifo1_data_ext_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:283" *)
  wire [31:0] pfifo1_data_ext_byte4_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:284" *)
  wire [31:0] pfifo1_data_ext_byte4_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:285" *)
  wire [31:0] pfifo1_data_ext_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:286" *)
  wire [31:0] pfifo1_data_ext_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:287" *)
  wire [31:0] pfifo1_data_ext_byte5_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:288" *)
  wire [31:0] pfifo1_data_ext_byte5_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:289" *)
  wire [31:0] pfifo1_data_ext_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:290" *)
  wire [31:0] pfifo1_data_ext_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:291" *)
  wire [31:0] pfifo1_data_ext_byte6_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:292" *)
  wire [31:0] pfifo1_data_ext_byte6_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:293" *)
  wire [31:0] pfifo1_data_ext_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:294" *)
  wire [31:0] pfifo1_data_ext_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:295" *)
  wire [31:0] pfifo1_data_ext_byte7_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:296" *)
  wire [31:0] pfifo1_data_ext_byte7_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:297" *)
  wire [31:0] pfifo1_data_ext_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:298" *)
  wire [31:0] pfifo1_data_ext_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:299" *)
  wire [127:0] pfifo1_rd_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:60" *)
  input [127:0] pfifo1_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:59" *)
  output pfifo1_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:58" *)
  input pfifo1_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:300" *)
  wire pfifo1_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:301" *)
  wire [255:0] pfifo2_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:302" *)
  wire [15:0] pfifo2_data_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:303" *)
  wire [7:0] pfifo2_data_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:304" *)
  wire pfifo2_data_byte0_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:305" *)
  wire pfifo2_data_byte0_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:306" *)
  wire [7:0] pfifo2_data_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:307" *)
  wire [7:0] pfifo2_data_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:308" *)
  wire [7:0] pfifo2_data_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:309" *)
  wire [7:0] pfifo2_data_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:310" *)
  wire [7:0] pfifo2_data_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:311" *)
  wire [7:0] pfifo2_data_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:312" *)
  wire [15:0] pfifo2_data_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:313" *)
  wire [7:0] pfifo2_data_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:314" *)
  wire pfifo2_data_byte1_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:315" *)
  wire pfifo2_data_byte1_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:316" *)
  wire [15:0] pfifo2_data_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:317" *)
  wire [7:0] pfifo2_data_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:318" *)
  wire pfifo2_data_byte2_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:319" *)
  wire pfifo2_data_byte2_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:320" *)
  wire [15:0] pfifo2_data_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:321" *)
  wire [7:0] pfifo2_data_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:322" *)
  wire pfifo2_data_byte3_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:323" *)
  wire pfifo2_data_byte3_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:324" *)
  wire [15:0] pfifo2_data_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:325" *)
  wire [7:0] pfifo2_data_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:326" *)
  wire pfifo2_data_byte4_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:327" *)
  wire pfifo2_data_byte4_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:328" *)
  wire [15:0] pfifo2_data_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:329" *)
  wire [7:0] pfifo2_data_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:330" *)
  wire pfifo2_data_byte5_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:331" *)
  wire pfifo2_data_byte5_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:332" *)
  wire [15:0] pfifo2_data_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:333" *)
  wire [7:0] pfifo2_data_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:334" *)
  wire pfifo2_data_byte6_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:335" *)
  wire pfifo2_data_byte6_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:336" *)
  wire [15:0] pfifo2_data_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:337" *)
  wire [7:0] pfifo2_data_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:338" *)
  wire pfifo2_data_byte7_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:339" *)
  wire pfifo2_data_byte7_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:340" *)
  wire [7:0] pfifo2_data_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:341" *)
  wire [7:0] pfifo2_data_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:342" *)
  wire [31:0] pfifo2_data_ext_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:343" *)
  wire [31:0] pfifo2_data_ext_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:344" *)
  wire [31:0] pfifo2_data_ext_byte0_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:345" *)
  wire [31:0] pfifo2_data_ext_byte0_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:346" *)
  wire [31:0] pfifo2_data_ext_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:347" *)
  wire [31:0] pfifo2_data_ext_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:348" *)
  wire [31:0] pfifo2_data_ext_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:349" *)
  wire [31:0] pfifo2_data_ext_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:350" *)
  wire [31:0] pfifo2_data_ext_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:351" *)
  wire [31:0] pfifo2_data_ext_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:352" *)
  wire [31:0] pfifo2_data_ext_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:353" *)
  wire [31:0] pfifo2_data_ext_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:354" *)
  wire [31:0] pfifo2_data_ext_byte1_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:355" *)
  wire [31:0] pfifo2_data_ext_byte1_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:356" *)
  wire [31:0] pfifo2_data_ext_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:357" *)
  wire [31:0] pfifo2_data_ext_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:358" *)
  wire [31:0] pfifo2_data_ext_byte2_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:359" *)
  wire [31:0] pfifo2_data_ext_byte2_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:360" *)
  wire [31:0] pfifo2_data_ext_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:361" *)
  wire [31:0] pfifo2_data_ext_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:362" *)
  wire [31:0] pfifo2_data_ext_byte3_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:363" *)
  wire [31:0] pfifo2_data_ext_byte3_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:364" *)
  wire [31:0] pfifo2_data_ext_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:365" *)
  wire [31:0] pfifo2_data_ext_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:366" *)
  wire [31:0] pfifo2_data_ext_byte4_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:367" *)
  wire [31:0] pfifo2_data_ext_byte4_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:368" *)
  wire [31:0] pfifo2_data_ext_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:369" *)
  wire [31:0] pfifo2_data_ext_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:370" *)
  wire [31:0] pfifo2_data_ext_byte5_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:371" *)
  wire [31:0] pfifo2_data_ext_byte5_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:372" *)
  wire [31:0] pfifo2_data_ext_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:373" *)
  wire [31:0] pfifo2_data_ext_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:374" *)
  wire [31:0] pfifo2_data_ext_byte6_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:375" *)
  wire [31:0] pfifo2_data_ext_byte6_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:376" *)
  wire [31:0] pfifo2_data_ext_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:377" *)
  wire [31:0] pfifo2_data_ext_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:378" *)
  wire [31:0] pfifo2_data_ext_byte7_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:379" *)
  wire [31:0] pfifo2_data_ext_byte7_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:380" *)
  wire [31:0] pfifo2_data_ext_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:381" *)
  wire [31:0] pfifo2_data_ext_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:382" *)
  wire [127:0] pfifo2_rd_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:63" *)
  input [127:0] pfifo2_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:62" *)
  output pfifo2_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:61" *)
  input pfifo2_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:383" *)
  wire pfifo2_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:384" *)
  wire [255:0] pfifo3_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:385" *)
  wire [15:0] pfifo3_data_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:386" *)
  wire [7:0] pfifo3_data_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:387" *)
  wire pfifo3_data_byte0_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:388" *)
  wire pfifo3_data_byte0_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:389" *)
  wire [7:0] pfifo3_data_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:390" *)
  wire [7:0] pfifo3_data_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:391" *)
  wire [7:0] pfifo3_data_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:392" *)
  wire [7:0] pfifo3_data_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:393" *)
  wire [7:0] pfifo3_data_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:394" *)
  wire [7:0] pfifo3_data_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:395" *)
  wire [15:0] pfifo3_data_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:396" *)
  wire [7:0] pfifo3_data_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:397" *)
  wire pfifo3_data_byte1_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:398" *)
  wire pfifo3_data_byte1_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:399" *)
  wire [15:0] pfifo3_data_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:400" *)
  wire [7:0] pfifo3_data_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:401" *)
  wire pfifo3_data_byte2_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:402" *)
  wire pfifo3_data_byte2_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:403" *)
  wire [15:0] pfifo3_data_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:404" *)
  wire [7:0] pfifo3_data_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:405" *)
  wire pfifo3_data_byte3_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:406" *)
  wire pfifo3_data_byte3_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:407" *)
  wire [15:0] pfifo3_data_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:408" *)
  wire [7:0] pfifo3_data_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:409" *)
  wire pfifo3_data_byte4_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:410" *)
  wire pfifo3_data_byte4_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:411" *)
  wire [15:0] pfifo3_data_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:412" *)
  wire [7:0] pfifo3_data_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:413" *)
  wire pfifo3_data_byte5_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:414" *)
  wire pfifo3_data_byte5_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:415" *)
  wire [15:0] pfifo3_data_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:416" *)
  wire [7:0] pfifo3_data_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:417" *)
  wire pfifo3_data_byte6_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:418" *)
  wire pfifo3_data_byte6_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:419" *)
  wire [15:0] pfifo3_data_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:420" *)
  wire [7:0] pfifo3_data_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:421" *)
  wire pfifo3_data_byte7_is_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:422" *)
  wire pfifo3_data_byte7_is_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:423" *)
  wire [7:0] pfifo3_data_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:424" *)
  wire [7:0] pfifo3_data_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:425" *)
  wire [31:0] pfifo3_data_ext_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:426" *)
  wire [31:0] pfifo3_data_ext_byte0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:427" *)
  wire [31:0] pfifo3_data_ext_byte0_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:428" *)
  wire [31:0] pfifo3_data_ext_byte0_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:429" *)
  wire [31:0] pfifo3_data_ext_byte10_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:430" *)
  wire [31:0] pfifo3_data_ext_byte11_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:431" *)
  wire [31:0] pfifo3_data_ext_byte12_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:432" *)
  wire [31:0] pfifo3_data_ext_byte13_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:433" *)
  wire [31:0] pfifo3_data_ext_byte14_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:434" *)
  wire [31:0] pfifo3_data_ext_byte15_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:435" *)
  wire [31:0] pfifo3_data_ext_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:436" *)
  wire [31:0] pfifo3_data_ext_byte1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:437" *)
  wire [31:0] pfifo3_data_ext_byte1_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:438" *)
  wire [31:0] pfifo3_data_ext_byte1_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:439" *)
  wire [31:0] pfifo3_data_ext_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:440" *)
  wire [31:0] pfifo3_data_ext_byte2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:441" *)
  wire [31:0] pfifo3_data_ext_byte2_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:442" *)
  wire [31:0] pfifo3_data_ext_byte2_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:443" *)
  wire [31:0] pfifo3_data_ext_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:444" *)
  wire [31:0] pfifo3_data_ext_byte3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:445" *)
  wire [31:0] pfifo3_data_ext_byte3_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:446" *)
  wire [31:0] pfifo3_data_ext_byte3_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:447" *)
  wire [31:0] pfifo3_data_ext_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:448" *)
  wire [31:0] pfifo3_data_ext_byte4_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:449" *)
  wire [31:0] pfifo3_data_ext_byte4_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:450" *)
  wire [31:0] pfifo3_data_ext_byte4_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:451" *)
  wire [31:0] pfifo3_data_ext_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:452" *)
  wire [31:0] pfifo3_data_ext_byte5_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:453" *)
  wire [31:0] pfifo3_data_ext_byte5_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:454" *)
  wire [31:0] pfifo3_data_ext_byte5_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:455" *)
  wire [31:0] pfifo3_data_ext_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:456" *)
  wire [31:0] pfifo3_data_ext_byte6_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:457" *)
  wire [31:0] pfifo3_data_ext_byte6_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:458" *)
  wire [31:0] pfifo3_data_ext_byte6_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:459" *)
  wire [31:0] pfifo3_data_ext_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:460" *)
  wire [31:0] pfifo3_data_ext_byte7_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:461" *)
  wire [31:0] pfifo3_data_ext_byte7_fp16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:462" *)
  wire [31:0] pfifo3_data_ext_byte7_int16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:463" *)
  wire [31:0] pfifo3_data_ext_byte8_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:464" *)
  wire [31:0] pfifo3_data_ext_byte9_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:465" *)
  wire [127:0] pfifo3_rd_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:66" *)
  input [127:0] pfifo3_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:65" *)
  output pfifo3_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:64" *)
  input pfifo3_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:466" *)
  wire pfifo3_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:467" *)
  wire [511:0] pfifo_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:468" *)
  wire [511:0] pfifo_data0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:469" *)
  wire [511:0] pfifo_data0_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:470" *)
  wire [511:0] pfifo_data1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:471" *)
  wire [511:0] pfifo_data1_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:472" *)
  wire [511:0] pfifo_data2_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:473" *)
  wire [511:0] pfifo_data3_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:90" *)
  wire [511:0] pfifo_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:91" *)
  wire [511:0] pfifo_data_8;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:474" *)
  wire pfifo_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:475" *)
  wire pfifo_vld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:78" *)
  input [12:0] reg2dp_height;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:79" *)
  input [1:0] reg2dp_in_precision;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:80" *)
  input reg2dp_perf_nan_inf_count_en;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:81" *)
  input [1:0] reg2dp_proc_precision;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:82" *)
  input [12:0] reg2dp_width;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:476" *)
  wire sdp_mrdma2cmux_layer_end;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:75" *)
  output [513:0] sdp_mrdma2cmux_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:74" *)
  input sdp_mrdma2cmux_ready;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:73" *)
  output sdp_mrdma2cmux_valid;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:477" *)
  wire [511:0] sfifo0_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:478" *)
  wire [15:0] sfifo0_data_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:479" *)
  wire [15:0] sfifo0_data_byte10_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:480" *)
  wire [15:0] sfifo0_data_byte11_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:481" *)
  wire [15:0] sfifo0_data_byte12_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:482" *)
  wire [15:0] sfifo0_data_byte13_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:483" *)
  wire [15:0] sfifo0_data_byte14_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:484" *)
  wire [15:0] sfifo0_data_byte15_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:485" *)
  wire [15:0] sfifo0_data_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:486" *)
  wire [15:0] sfifo0_data_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:487" *)
  wire [15:0] sfifo0_data_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:488" *)
  wire [15:0] sfifo0_data_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:489" *)
  wire [15:0] sfifo0_data_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:490" *)
  wire [15:0] sfifo0_data_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:491" *)
  wire [15:0] sfifo0_data_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:492" *)
  wire [15:0] sfifo0_data_byte8_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:493" *)
  wire [15:0] sfifo0_data_byte9_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:494" *)
  wire [31:0] sfifo0_data_ext_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:495" *)
  wire [31:0] sfifo0_data_ext_byte10_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:496" *)
  wire [31:0] sfifo0_data_ext_byte11_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:497" *)
  wire [31:0] sfifo0_data_ext_byte12_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:498" *)
  wire [31:0] sfifo0_data_ext_byte13_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:499" *)
  wire [31:0] sfifo0_data_ext_byte14_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:500" *)
  wire [31:0] sfifo0_data_ext_byte15_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:501" *)
  wire [31:0] sfifo0_data_ext_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:502" *)
  wire [31:0] sfifo0_data_ext_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:503" *)
  wire [31:0] sfifo0_data_ext_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:504" *)
  wire [31:0] sfifo0_data_ext_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:505" *)
  wire [31:0] sfifo0_data_ext_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:506" *)
  wire [31:0] sfifo0_data_ext_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:507" *)
  wire [31:0] sfifo0_data_ext_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:508" *)
  wire [31:0] sfifo0_data_ext_byte8_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:509" *)
  wire [31:0] sfifo0_data_ext_byte9_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:510" *)
  wire [255:0] sfifo0_rd_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:69" *)
  input [255:0] sfifo0_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:68" *)
  output sfifo0_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:67" *)
  input sfifo0_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:511" *)
  wire sfifo0_sel;
  wire [351:0] sfifo1_data_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:513" *)
  wire [15:0] sfifo1_data_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:514" *)
  wire [15:0] sfifo1_data_byte10_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:515" *)
  wire [15:0] sfifo1_data_byte11_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:516" *)
  wire [15:0] sfifo1_data_byte12_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:517" *)
  wire [15:0] sfifo1_data_byte13_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:518" *)
  wire [15:0] sfifo1_data_byte14_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:519" *)
  wire [15:0] sfifo1_data_byte15_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:520" *)
  wire [15:0] sfifo1_data_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:521" *)
  wire [15:0] sfifo1_data_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:522" *)
  wire [15:0] sfifo1_data_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:523" *)
  wire [15:0] sfifo1_data_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:524" *)
  wire [15:0] sfifo1_data_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:525" *)
  wire [15:0] sfifo1_data_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:526" *)
  wire [15:0] sfifo1_data_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:527" *)
  wire [15:0] sfifo1_data_byte8_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:528" *)
  wire [15:0] sfifo1_data_byte9_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:529" *)
  wire [31:0] sfifo1_data_ext_byte0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:530" *)
  wire [31:0] sfifo1_data_ext_byte10_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:531" *)
  wire [31:0] sfifo1_data_ext_byte11_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:532" *)
  wire [31:0] sfifo1_data_ext_byte12_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:533" *)
  wire [31:0] sfifo1_data_ext_byte13_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:534" *)
  wire [31:0] sfifo1_data_ext_byte14_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:535" *)
  wire [31:0] sfifo1_data_ext_byte15_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:536" *)
  wire [31:0] sfifo1_data_ext_byte1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:537" *)
  wire [31:0] sfifo1_data_ext_byte2_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:538" *)
  wire [31:0] sfifo1_data_ext_byte3_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:539" *)
  wire [31:0] sfifo1_data_ext_byte4_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:540" *)
  wire [31:0] sfifo1_data_ext_byte5_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:541" *)
  wire [31:0] sfifo1_data_ext_byte6_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:542" *)
  wire [31:0] sfifo1_data_ext_byte7_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:543" *)
  wire [31:0] sfifo1_data_ext_byte8_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:544" *)
  wire [31:0] sfifo1_data_ext_byte9_16;
  wire [175:0] sfifo1_rd_data;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:72" *)
  input [255:0] sfifo1_rd_pd;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:71" *)
  output sfifo1_rd_prdy;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:70" *)
  input sfifo1_rd_pvld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:546" *)
  wire sfifo1_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:92" *)
  wire [511:0] sfifo_data;
  wire [352:0] sfifo_data0_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:548" *)
  wire [511:0] sfifo_data1_16;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:549" *)
  wire sfifo_sel;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:550" *)
  wire sfifo_vld;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:551" *)
  wire [13:0] size_of_beat;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:552" *)
  wire [4:0] sum0_of_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:553" *)
  wire [4:0] sum0_of_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:554" *)
  wire [4:0] sum1_of_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:555" *)
  wire [4:0] sum1_of_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:556" *)
  wire [4:0] sum_of_inf;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:557" *)
  wire [4:0] sum_of_nan;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:558" *)
  wire sum_of_sel;
  assign _0324_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0676_;
  assign _0325_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0677_;
  assign _0326_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0678_;
  assign _0327_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0679_;
  assign _0328_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) { _0780_[3:1], _0680_ };
  assign _0329_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0681_;
  assign _0330_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0682_;
  assign _0331_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0683_;
  assign _0332_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0684_;
  assign _0333_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0685_;
  assign _0334_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0686_;
  assign _0335_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0687_;
  assign _0336_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0688_;
  assign _0337_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0689_;
  assign _0338_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0690_;
  assign _0339_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0691_;
  assign _0340_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0692_;
  assign _0341_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0693_;
  assign _0342_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0694_;
  assign _0343_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0695_;
  assign _0344_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) { _0781_[3:1], _0696_ };
  assign _0345_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0697_;
  assign _0346_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0698_;
  assign _0347_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0699_;
  assign _0348_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0700_;
  assign _0349_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0701_;
  assign _0350_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0702_;
  assign _0351_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0703_;
  assign _0352_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0704_;
  assign _0353_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0705_;
  assign _0354_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0706_;
  assign _0355_ = 4'b1101 + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0707_;
  assign _0356_ = pfifo0_rd_data[14:10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0357_ = pfifo0_rd_data[30:26] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0358_ = pfifo0_rd_data[46:42] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0359_ = pfifo0_rd_data[62:58] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0360_ = pfifo0_rd_data[78:74] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0361_ = pfifo0_rd_data[94:90] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0362_ = pfifo0_rd_data[110:106] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0363_ = pfifo0_rd_data[126:122] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0364_ = pfifo1_rd_data[14:10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0365_ = pfifo1_rd_data[30:26] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0366_ = pfifo1_rd_data[46:42] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0367_ = pfifo1_rd_data[62:58] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0368_ = pfifo1_rd_data[78:74] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0369_ = pfifo1_rd_data[94:90] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0370_ = pfifo1_rd_data[110:106] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0371_ = pfifo1_rd_data[126:122] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0372_ = pfifo2_rd_data[14:10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0373_ = pfifo2_rd_data[30:26] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0374_ = pfifo2_rd_data[46:42] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0375_ = pfifo2_rd_data[62:58] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0376_ = pfifo2_rd_data[78:74] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0377_ = pfifo2_rd_data[94:90] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0378_ = pfifo2_rd_data[110:106] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0379_ = pfifo2_rd_data[126:122] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0380_ = pfifo3_rd_data[14:10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0381_ = pfifo3_rd_data[30:26] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0382_ = pfifo3_rd_data[46:42] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0383_ = pfifo3_rd_data[62:58] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0384_ = pfifo3_rd_data[78:74] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0385_ = pfifo3_rd_data[94:90] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0386_ = pfifo3_rd_data[110:106] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0387_ = pfifo3_rd_data[126:122] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1459" *) 7'b1110000;
  assign _0388_ = _0782_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0782_[9];
  assign _0389_ = _0783_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0783_[9];
  assign _0390_ = _0784_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0784_[9];
  assign _0391_ = _0785_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0785_[9];
  assign _0392_ = _0786_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0786_[9];
  assign _0393_ = _0787_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0787_[9];
  assign _0394_ = _0788_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0788_[9];
  assign _0395_ = _0789_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0789_[9];
  assign _0396_ = _0790_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0790_[9];
  assign _0397_ = _0791_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0791_[9];
  assign _0398_ = _0792_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0792_[9];
  assign _0399_ = _0793_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0793_[9];
  assign _0400_ = _0794_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0794_[9];
  assign _0401_ = _0795_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0795_[9];
  assign _0402_ = _0796_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0796_[9];
  assign _0403_ = _0797_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0797_[9];
  assign _0404_ = _0798_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0798_[9];
  assign _0405_ = _0799_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0799_[9];
  assign _0406_ = _0800_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0800_[9];
  assign _0407_ = _0801_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0801_[9];
  assign _0408_ = _0802_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0802_[9];
  assign _0409_ = _0803_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0803_[9];
  assign _0410_ = _0804_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0804_[9];
  assign _0411_ = _0805_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0805_[9];
  assign _0412_ = _0806_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0806_[9];
  assign _0413_ = _0807_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0807_[9];
  assign _0414_ = _0808_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0808_[9];
  assign _0415_ = _0809_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0809_[9];
  assign _0416_ = _0810_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0810_[9];
  assign _0417_ = _0811_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0811_[9];
  assign _0418_ = _0812_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0812_[9];
  assign _0419_ = _0813_[10] + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1487" *) _0813_[9];
  assign _0420_ = _0388_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0782_[8];
  assign _0421_ = _0389_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0783_[8];
  assign _0422_ = _0390_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0784_[8];
  assign _0423_ = _0391_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0785_[8];
  assign _0424_ = _0392_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0786_[8];
  assign _0425_ = _0393_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0787_[8];
  assign _0426_ = _0394_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0788_[8];
  assign _0427_ = _0395_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0789_[8];
  assign _0428_ = _0396_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0790_[8];
  assign _0429_ = _0397_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0791_[8];
  assign _0430_ = _0398_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0792_[8];
  assign _0431_ = _0399_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0793_[8];
  assign _0432_ = _0400_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0794_[8];
  assign _0433_ = _0401_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0795_[8];
  assign _0434_ = _0402_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0796_[8];
  assign _0435_ = _0403_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0797_[8];
  assign _0436_ = _0404_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0798_[8];
  assign _0437_ = _0405_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0799_[8];
  assign _0438_ = _0406_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0800_[8];
  assign _0439_ = _0407_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0801_[8];
  assign _0440_ = _0408_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0802_[8];
  assign _0441_ = _0409_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0803_[8];
  assign _0442_ = _0410_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0804_[8];
  assign _0443_ = _0411_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0805_[8];
  assign _0444_ = _0412_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0806_[8];
  assign _0445_ = _0413_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0807_[8];
  assign _0446_ = _0414_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0808_[8];
  assign _0447_ = _0415_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0809_[8];
  assign _0448_ = _0416_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0810_[8];
  assign _0449_ = _0417_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0811_[8];
  assign _0450_ = _0418_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0812_[8];
  assign _0451_ = _0419_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1488" *) _0813_[8];
  assign _0452_ = _0420_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0782_[7];
  assign _0453_ = _0421_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0783_[7];
  assign _0454_ = _0422_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0784_[7];
  assign _0455_ = _0423_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0785_[7];
  assign _0456_ = _0424_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0786_[7];
  assign _0457_ = _0425_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0787_[7];
  assign _0458_ = _0426_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0788_[7];
  assign _0459_ = _0427_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0789_[7];
  assign _0460_ = _0428_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0790_[7];
  assign _0461_ = _0429_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0791_[7];
  assign _0462_ = _0430_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0792_[7];
  assign _0463_ = _0431_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0793_[7];
  assign _0464_ = _0432_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0794_[7];
  assign _0465_ = _0433_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0795_[7];
  assign _0466_ = _0434_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0796_[7];
  assign _0467_ = _0435_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0797_[7];
  assign _0468_ = _0436_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0798_[7];
  assign _0469_ = _0437_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0799_[7];
  assign _0470_ = _0438_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0800_[7];
  assign _0471_ = _0439_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0801_[7];
  assign _0472_ = _0440_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0802_[7];
  assign _0473_ = _0441_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0803_[7];
  assign _0474_ = _0442_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0804_[7];
  assign _0475_ = _0443_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0805_[7];
  assign _0476_ = _0444_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0806_[7];
  assign _0477_ = _0445_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0807_[7];
  assign _0478_ = _0446_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0808_[7];
  assign _0479_ = _0447_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0809_[7];
  assign _0480_ = _0448_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0810_[7];
  assign _0481_ = _0449_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0811_[7];
  assign _0482_ = _0450_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0812_[7];
  assign _0483_ = _0451_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1489" *) _0813_[7];
  assign _0484_ = _0452_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0782_[6];
  assign _0485_ = _0453_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0783_[6];
  assign _0486_ = _0454_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0784_[6];
  assign _0487_ = _0455_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0785_[6];
  assign _0488_ = _0456_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0786_[6];
  assign _0489_ = _0457_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0787_[6];
  assign _0490_ = _0458_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0788_[6];
  assign _0491_ = _0459_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0789_[6];
  assign _0492_ = _0460_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0790_[6];
  assign _0493_ = _0461_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0791_[6];
  assign _0494_ = _0462_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0792_[6];
  assign _0495_ = _0463_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0793_[6];
  assign _0496_ = _0464_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0794_[6];
  assign _0497_ = _0465_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0795_[6];
  assign _0498_ = _0466_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0796_[6];
  assign _0499_ = _0467_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0797_[6];
  assign _0500_ = _0468_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0798_[6];
  assign _0501_ = _0469_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0799_[6];
  assign _0502_ = _0470_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0800_[6];
  assign _0503_ = _0471_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0801_[6];
  assign _0504_ = _0472_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0802_[6];
  assign _0505_ = _0473_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0803_[6];
  assign _0506_ = _0474_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0804_[6];
  assign _0507_ = _0475_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0805_[6];
  assign _0508_ = _0476_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0806_[6];
  assign _0509_ = _0477_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0807_[6];
  assign _0510_ = _0478_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0808_[6];
  assign _0511_ = _0479_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0809_[6];
  assign _0512_ = _0480_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0810_[6];
  assign _0513_ = _0481_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0811_[6];
  assign _0514_ = _0482_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0812_[6];
  assign _0515_ = _0483_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1490" *) _0813_[6];
  assign _0516_ = _0484_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0782_[5];
  assign _0517_ = _0485_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0783_[5];
  assign _0518_ = _0486_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0784_[5];
  assign _0519_ = _0487_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0785_[5];
  assign _0520_ = _0488_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0786_[5];
  assign _0521_ = _0489_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0787_[5];
  assign _0522_ = _0490_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0788_[5];
  assign _0523_ = _0491_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0789_[5];
  assign _0524_ = _0492_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0790_[5];
  assign _0525_ = _0493_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0791_[5];
  assign _0526_ = _0494_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0792_[5];
  assign _0527_ = _0495_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0793_[5];
  assign _0528_ = _0496_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0794_[5];
  assign _0529_ = _0497_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0795_[5];
  assign _0530_ = _0498_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0796_[5];
  assign _0531_ = _0499_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0797_[5];
  assign _0532_ = _0500_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0798_[5];
  assign _0533_ = _0501_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0799_[5];
  assign _0534_ = _0502_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0800_[5];
  assign _0535_ = _0503_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0801_[5];
  assign _0536_ = _0504_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0802_[5];
  assign _0537_ = _0505_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0803_[5];
  assign _0538_ = _0506_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0804_[5];
  assign _0539_ = _0507_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0805_[5];
  assign _0540_ = _0508_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0806_[5];
  assign _0541_ = _0509_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0807_[5];
  assign _0542_ = _0510_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0808_[5];
  assign _0543_ = _0511_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0809_[5];
  assign _0544_ = _0512_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0810_[5];
  assign _0545_ = _0513_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0811_[5];
  assign _0546_ = _0514_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0812_[5];
  assign _0547_ = _0515_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1491" *) _0813_[5];
  assign _0548_ = _0516_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0782_[4];
  assign _0549_ = _0517_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0783_[4];
  assign _0550_ = _0518_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0784_[4];
  assign _0551_ = _0519_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0785_[4];
  assign _0552_ = _0520_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0786_[4];
  assign _0553_ = _0521_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0787_[4];
  assign _0554_ = _0522_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0788_[4];
  assign _0555_ = _0523_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0789_[4];
  assign _0556_ = _0524_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0790_[4];
  assign _0557_ = _0525_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0791_[4];
  assign _0558_ = _0526_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0792_[4];
  assign _0559_ = _0527_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0793_[4];
  assign _0560_ = _0528_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0794_[4];
  assign _0561_ = _0529_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0795_[4];
  assign _0562_ = _0530_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0796_[4];
  assign _0563_ = _0531_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0797_[4];
  assign _0564_ = _0532_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0798_[4];
  assign _0565_ = _0533_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0799_[4];
  assign _0566_ = _0534_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0800_[4];
  assign _0567_ = _0535_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0801_[4];
  assign _0568_ = _0536_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0802_[4];
  assign _0569_ = _0537_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0803_[4];
  assign _0570_ = _0538_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0804_[4];
  assign _0571_ = _0539_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0805_[4];
  assign _0572_ = _0540_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0806_[4];
  assign _0573_ = _0541_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0807_[4];
  assign _0574_ = _0542_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0808_[4];
  assign _0575_ = _0543_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0809_[4];
  assign _0576_ = _0544_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0810_[4];
  assign _0577_ = _0545_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0811_[4];
  assign _0578_ = _0546_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0812_[4];
  assign _0579_ = _0547_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1492" *) _0813_[4];
  assign _0580_ = _0548_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0782_[3];
  assign _0581_ = _0549_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0783_[3];
  assign _0582_ = _0550_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0784_[3];
  assign _0583_ = _0551_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0785_[3];
  assign _0584_ = _0552_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0786_[3];
  assign _0585_ = _0553_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0787_[3];
  assign _0586_ = _0554_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0788_[3];
  assign _0587_ = _0555_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0789_[3];
  assign _0588_ = _0556_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0790_[3];
  assign _0589_ = _0557_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0791_[3];
  assign _0590_ = _0558_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0792_[3];
  assign _0591_ = _0559_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0793_[3];
  assign _0592_ = _0560_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0794_[3];
  assign _0593_ = _0561_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0795_[3];
  assign _0594_ = _0562_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0796_[3];
  assign _0595_ = _0563_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0797_[3];
  assign _0596_ = _0564_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0798_[3];
  assign _0597_ = _0565_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0799_[3];
  assign _0598_ = _0566_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0800_[3];
  assign _0599_ = _0567_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0801_[3];
  assign _0600_ = _0568_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0802_[3];
  assign _0601_ = _0569_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0803_[3];
  assign _0602_ = _0570_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0804_[3];
  assign _0603_ = _0571_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0805_[3];
  assign _0604_ = _0572_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0806_[3];
  assign _0605_ = _0573_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0807_[3];
  assign _0606_ = _0574_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0808_[3];
  assign _0607_ = _0575_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0809_[3];
  assign _0608_ = _0576_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0810_[3];
  assign _0609_ = _0577_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0811_[3];
  assign _0610_ = _0578_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0812_[3];
  assign _0611_ = _0579_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1493" *) _0813_[3];
  assign _0612_ = _0580_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0782_[2];
  assign _0613_ = _0581_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0783_[2];
  assign _0614_ = _0582_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0784_[2];
  assign _0615_ = _0583_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0785_[2];
  assign _0616_ = _0584_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0786_[2];
  assign _0617_ = _0585_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0787_[2];
  assign _0618_ = _0586_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0788_[2];
  assign _0619_ = _0587_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0789_[2];
  assign _0620_ = _0588_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0790_[2];
  assign _0621_ = _0589_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0791_[2];
  assign _0622_ = _0590_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0792_[2];
  assign _0623_ = _0591_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0793_[2];
  assign _0624_ = _0592_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0794_[2];
  assign _0625_ = _0593_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0795_[2];
  assign _0626_ = _0594_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0796_[2];
  assign _0627_ = _0595_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0797_[2];
  assign _0628_ = _0596_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0798_[2];
  assign _0629_ = _0597_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0799_[2];
  assign _0630_ = _0598_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0800_[2];
  assign _0631_ = _0599_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0801_[2];
  assign _0632_ = _0600_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0802_[2];
  assign _0633_ = _0601_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0803_[2];
  assign _0634_ = _0602_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0804_[2];
  assign _0635_ = _0603_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0805_[2];
  assign _0636_ = _0604_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0806_[2];
  assign _0637_ = _0605_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0807_[2];
  assign _0638_ = _0606_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0808_[2];
  assign _0639_ = _0607_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0809_[2];
  assign _0640_ = _0608_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0810_[2];
  assign _0641_ = _0609_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0811_[2];
  assign _0642_ = _0610_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0812_[2];
  assign _0643_ = _0611_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1494" *) _0813_[2];
  assign _0644_ = _0612_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0782_[1];
  assign _0645_ = _0613_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0783_[1];
  assign _0646_ = _0614_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0784_[1];
  assign _0647_ = _0615_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0785_[1];
  assign _0648_ = _0616_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0786_[1];
  assign _0649_ = _0617_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0787_[1];
  assign _0650_ = _0618_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0788_[1];
  assign _0651_ = _0619_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0789_[1];
  assign _0652_ = _0620_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0790_[1];
  assign _0653_ = _0621_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0791_[1];
  assign _0654_ = _0622_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0792_[1];
  assign _0655_ = _0623_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0793_[1];
  assign _0656_ = _0624_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0794_[1];
  assign _0657_ = _0625_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0795_[1];
  assign _0658_ = _0626_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0796_[1];
  assign _0659_ = _0627_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0797_[1];
  assign _0660_ = _0628_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0798_[1];
  assign _0661_ = _0629_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0799_[1];
  assign _0662_ = _0630_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0800_[1];
  assign _0663_ = _0631_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0801_[1];
  assign _0664_ = _0632_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0802_[1];
  assign _0665_ = _0633_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0803_[1];
  assign _0666_ = _0634_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0804_[1];
  assign _0667_ = _0635_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0805_[1];
  assign _0668_ = _0636_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0806_[1];
  assign _0669_ = _0637_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0807_[1];
  assign _0670_ = _0638_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0808_[1];
  assign _0671_ = _0639_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0809_[1];
  assign _0672_ = _0640_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0810_[1];
  assign _0673_ = _0641_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0811_[1];
  assign _0674_ = _0642_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0812_[1];
  assign _0675_ = _0643_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1495" *) _0813_[1];
  assign _0676_ = _0644_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0782_[0];
  assign _0677_ = _0645_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0783_[0];
  assign _0678_ = _0646_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0784_[0];
  assign _0679_ = _0647_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0785_[0];
  assign { _0780_[3:1], _0680_ } = _0648_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0786_[0];
  assign _0681_ = _0649_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0787_[0];
  assign _0682_ = _0650_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0788_[0];
  assign _0683_ = _0651_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0789_[0];
  assign _0684_ = _0652_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0790_[0];
  assign _0685_ = _0653_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0791_[0];
  assign _0686_ = _0654_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0792_[0];
  assign _0687_ = _0655_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0793_[0];
  assign _0688_ = _0656_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0794_[0];
  assign _0689_ = _0657_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0795_[0];
  assign _0690_ = _0658_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0796_[0];
  assign _0691_ = _0659_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0797_[0];
  assign _0692_ = _0660_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0798_[0];
  assign _0693_ = _0661_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0799_[0];
  assign _0694_ = _0662_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0800_[0];
  assign _0695_ = _0663_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0801_[0];
  assign { _0781_[3:1], _0696_ } = _0664_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0802_[0];
  assign _0697_ = _0665_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0803_[0];
  assign _0698_ = _0666_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0804_[0];
  assign _0699_ = _0667_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0805_[0];
  assign _0700_ = _0668_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0806_[0];
  assign _0701_ = _0669_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0807_[0];
  assign _0702_ = _0670_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0808_[0];
  assign _0703_ = _0671_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0809_[0];
  assign _0704_ = _0672_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0810_[0];
  assign _0705_ = _0673_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0811_[0];
  assign _0706_ = _0674_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0812_[0];
  assign _0707_ = _0675_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1496" *) _0813_[0];
  assign _0708_ = beat_cnt + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:595" *) 1'b1;
  assign _0709_ = pfifo1_data_byte7_is_inf + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte6_is_inf;
  assign _0710_ = _0709_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte5_is_inf;
  assign _0711_ = _0710_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte4_is_inf;
  assign _0712_ = _0711_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte3_is_inf;
  assign _0713_ = _0712_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte2_is_inf;
  assign _0714_ = _0713_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte1_is_inf;
  assign _0715_ = _0714_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo1_data_byte0_is_inf;
  assign _0716_ = _0715_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte7_is_inf;
  assign _0717_ = _0716_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte6_is_inf;
  assign _0718_ = _0717_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte5_is_inf;
  assign _0719_ = _0718_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte4_is_inf;
  assign _0720_ = _0719_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte3_is_inf;
  assign _0721_ = _0720_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte2_is_inf;
  assign _0722_ = _0721_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte1_is_inf;
  assign sum0_of_inf = _0722_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:635" *) pfifo0_data_byte0_is_inf;
  assign _0723_ = pfifo3_data_byte7_is_inf + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte6_is_inf;
  assign _0724_ = _0723_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte5_is_inf;
  assign _0725_ = _0724_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte4_is_inf;
  assign _0726_ = _0725_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte3_is_inf;
  assign _0727_ = _0726_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte2_is_inf;
  assign _0728_ = _0727_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte1_is_inf;
  assign _0729_ = _0728_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo3_data_byte0_is_inf;
  assign _0730_ = _0729_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte7_is_inf;
  assign _0731_ = _0730_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte6_is_inf;
  assign _0732_ = _0731_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte5_is_inf;
  assign _0733_ = _0732_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte4_is_inf;
  assign _0734_ = _0733_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte3_is_inf;
  assign _0735_ = _0734_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte2_is_inf;
  assign _0736_ = _0735_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte1_is_inf;
  assign sum1_of_inf = _0736_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:636" *) pfifo2_data_byte0_is_inf;
  assign { inf_input_cnt_nxt_c, inf_input_cnt_nxt } = inf_input_cnt + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:638" *) sum_of_inf;
  assign _0737_ = pfifo1_data_byte7_is_nan + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte6_is_nan;
  assign _0738_ = _0737_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte5_is_nan;
  assign _0739_ = _0738_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte4_is_nan;
  assign _0740_ = _0739_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte3_is_nan;
  assign _0741_ = _0740_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte2_is_nan;
  assign _0742_ = _0741_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte1_is_nan;
  assign _0743_ = _0742_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo1_data_byte0_is_nan;
  assign _0744_ = _0743_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte7_is_nan;
  assign _0745_ = _0744_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte6_is_nan;
  assign _0746_ = _0745_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte5_is_nan;
  assign _0747_ = _0746_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte4_is_nan;
  assign _0748_ = _0747_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte3_is_nan;
  assign _0749_ = _0748_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte2_is_nan;
  assign _0750_ = _0749_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte1_is_nan;
  assign sum0_of_nan = _0750_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:689" *) pfifo0_data_byte0_is_nan;
  assign _0751_ = pfifo3_data_byte7_is_nan + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte6_is_nan;
  assign _0752_ = _0751_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte5_is_nan;
  assign _0753_ = _0752_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte4_is_nan;
  assign _0754_ = _0753_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte3_is_nan;
  assign _0755_ = _0754_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte2_is_nan;
  assign _0756_ = _0755_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte1_is_nan;
  assign _0757_ = _0756_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo3_data_byte0_is_nan;
  assign _0758_ = _0757_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte7_is_nan;
  assign _0759_ = _0758_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte6_is_nan;
  assign _0760_ = _0759_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte5_is_nan;
  assign _0761_ = _0760_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte4_is_nan;
  assign _0762_ = _0761_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte3_is_nan;
  assign _0763_ = _0762_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte2_is_nan;
  assign _0764_ = _0763_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte1_is_nan;
  assign sum1_of_nan = _0764_ + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:690" *) pfifo2_data_byte0_is_nan;
  assign { nan_input_cnt_nxt_c, nan_input_cnt_nxt } = nan_input_cnt + (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:692" *) sum_of_nan;
  assign sfifo0_rd_data = { sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel, sfifo0_sel } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1027" *) sfifo0_rd_pd;
  assign { sfifo1_data_byte15_16, sfifo1_data_byte14_16, sfifo1_data_byte13_16, sfifo1_data_byte12_16, sfifo1_data_byte11_16, sfifo1_data_16[351], sfifo1_data_16[334:319], sfifo1_data_16[302:287], sfifo1_data_16[270:255], sfifo1_data_16[238:223], sfifo1_data_16[206:191], sfifo1_data_16[174:159], sfifo1_data_16[142:127], sfifo1_data_16[110:95], sfifo1_data_16[78:63], sfifo1_data_16[46:31], sfifo1_data_16[14:0] } = { sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel, sfifo1_sel } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1028" *) sfifo1_rd_pd;
  assign dat_accept = dat_vld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1159" *) dat_rdy;
  assign dat_batch_end = cmd_cube_end & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1160" *) is_last_beat;
  assign _0765_ = sdp_mrdma2cmux_pd[513] & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1185" *) sdp_mrdma2cmux_valid;
  assign _0129_ = _0765_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1185" *) sdp_mrdma2cmux_ready;
  assign _0003_ = _0868_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0869_;
  assign _0007_ = _0870_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0871_;
  assign _0011_ = _0872_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0873_;
  assign _0015_ = _0874_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0875_;
  assign _0019_ = _0876_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0877_;
  assign _0023_ = _0878_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0879_;
  assign _0027_ = _0880_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0881_;
  assign _0031_ = _0882_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0883_;
  assign _0035_ = _0884_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0885_;
  assign _0039_ = _0886_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0887_;
  assign _0043_ = _0888_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0889_;
  assign _0047_ = _0890_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0891_;
  assign _0051_ = _0892_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0893_;
  assign _0055_ = _0894_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0895_;
  assign _0059_ = _0896_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0897_;
  assign _0063_ = _0898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0899_;
  assign _0067_ = _0900_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0901_;
  assign _0071_ = _0902_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0903_;
  assign _0075_ = _0904_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0905_;
  assign _0079_ = _0906_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0907_;
  assign _0083_ = _0908_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0909_;
  assign _0087_ = _0910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0911_;
  assign _0091_ = _0912_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0913_;
  assign _0095_ = _0914_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0915_;
  assign _0099_ = _0916_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0917_;
  assign _0103_ = _0918_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0919_;
  assign _0107_ = _0920_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0921_;
  assign _0111_ = _0922_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0923_;
  assign _0115_ = _0924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0925_;
  assign _0119_ = _0926_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0927_;
  assign _0123_ = _0928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0929_;
  assign _0127_ = _0930_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0931_;
  assign _0000_ = _0868_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0932_;
  assign _0004_ = _0870_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0933_;
  assign _0008_ = _0872_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0934_;
  assign _0012_ = _0874_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0935_;
  assign _0016_ = _0876_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0936_;
  assign _0020_ = _0878_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0937_;
  assign _0024_ = _0880_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0938_;
  assign _0028_ = _0882_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0939_;
  assign _0032_ = _0884_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0940_;
  assign _0036_ = _0886_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0941_;
  assign _0040_ = _0888_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0942_;
  assign _0044_ = _0890_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0943_;
  assign _0048_ = _0892_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0944_;
  assign _0052_ = _0894_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0945_;
  assign _0056_ = _0896_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0946_;
  assign _0060_ = _0898_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0947_;
  assign _0064_ = _0900_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0948_;
  assign _0068_ = _0902_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0949_;
  assign _0072_ = _0904_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0950_;
  assign _0076_ = _0906_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0951_;
  assign _0080_ = _0908_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0952_;
  assign _0084_ = _0910_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0953_;
  assign _0088_ = _0912_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0954_;
  assign _0092_ = _0914_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0955_;
  assign _0096_ = _0916_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0956_;
  assign _0100_ = _0918_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0957_;
  assign _0104_ = _0920_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0958_;
  assign _0108_ = _0922_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0959_;
  assign _0112_ = _0924_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0960_;
  assign _0116_ = _0926_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0961_;
  assign _0120_ = _0928_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0962_;
  assign _0124_ = _0930_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1438" *) _0963_;
  assign _0002_ = _0964_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0932_;
  assign _0006_ = _0965_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0933_;
  assign _0010_ = _0966_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0934_;
  assign _0014_ = _0967_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0935_;
  assign _0018_ = _0968_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0936_;
  assign _0022_ = _0969_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0937_;
  assign _0026_ = _0970_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0938_;
  assign _0030_ = _0971_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0939_;
  assign _0034_ = _0972_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0940_;
  assign _0038_ = _0973_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0941_;
  assign _0042_ = _0974_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0942_;
  assign _0046_ = _0975_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0943_;
  assign _0050_ = _0976_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0944_;
  assign _0054_ = _0977_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0945_;
  assign _0058_ = _0978_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0946_;
  assign _0062_ = _0979_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0947_;
  assign _0066_ = _0980_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0948_;
  assign _0070_ = _0981_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0949_;
  assign _0074_ = _0982_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0950_;
  assign _0078_ = _0983_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0951_;
  assign _0082_ = _0984_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0952_;
  assign _0086_ = _0985_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0953_;
  assign _0090_ = _0986_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0954_;
  assign _0094_ = _0987_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0955_;
  assign _0098_ = _0988_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0956_;
  assign _0102_ = _0989_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0957_;
  assign _0106_ = _0990_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0958_;
  assign _0110_ = _0991_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0959_;
  assign _0114_ = _0992_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0960_;
  assign _0118_ = _0993_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0961_;
  assign _0122_ = _0994_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0962_;
  assign _0126_ = _0995_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) _0963_;
  assign _0001_ = _0964_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0869_;
  assign _0005_ = _0965_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0871_;
  assign _0009_ = _0966_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0873_;
  assign _0013_ = _0967_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0875_;
  assign _0017_ = _0968_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0877_;
  assign _0021_ = _0969_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0879_;
  assign _0025_ = _0970_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0881_;
  assign _0029_ = _0971_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0883_;
  assign _0033_ = _0972_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0885_;
  assign _0037_ = _0973_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0887_;
  assign _0041_ = _0974_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0889_;
  assign _0045_ = _0975_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0891_;
  assign _0049_ = _0976_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0893_;
  assign _0053_ = _0977_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0895_;
  assign _0057_ = _0978_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0897_;
  assign _0061_ = _0979_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0899_;
  assign _0065_ = _0980_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0901_;
  assign _0069_ = _0981_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0903_;
  assign _0073_ = _0982_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0905_;
  assign _0077_ = _0983_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0907_;
  assign _0081_ = _0984_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0909_;
  assign _0085_ = _0985_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0911_;
  assign _0089_ = _0986_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0913_;
  assign _0093_ = _0987_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0915_;
  assign _0097_ = _0988_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0917_;
  assign _0101_ = _0989_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0919_;
  assign _0105_ = _0990_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0921_;
  assign _0109_ = _0991_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0923_;
  assign _0113_ = _0992_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0925_;
  assign _0117_ = _0993_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0927_;
  assign _0121_ = _0994_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0929_;
  assign _0125_ = _0995_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1440" *) _0931_;
  assign cfg_mode_16to8 = cfg_di_int16 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:577" *) cfg_do_int8;
  assign cfg_mode_1x1_pack = _0996_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:578" *) _0997_;
  assign _0766_ = dat_accept & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:580" *) is_last_beat;
  assign _0767_ = _0766_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:580" *) fifo_vld;
  assign cmd2dat_dma_prdy = _0767_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:580" *) dat_rdy;
  assign size_of_beat = { cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld, cmd2dat_dma_pvld } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:585" *) cmd2dat_dma_pd[13:0];
  assign cmd_cube_end = cmd2dat_dma_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:586" *) cmd2dat_dma_pd[14];
  assign _0768_ = pfifo3_rd_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) pfifo3_sel;
  assign _0769_ = pfifo2_rd_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) pfifo2_sel;
  assign _0770_ = pfifo1_rd_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) pfifo1_sel;
  assign _0771_ = pfifo0_rd_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) pfifo0_sel;
  assign _0772_ = sfifo1_rd_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:738" *) sfifo1_sel;
  assign _0773_ = sfifo0_rd_pvld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:738" *) sfifo0_sel;
  assign dat_vld = fifo_vld & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:740" *) cmd2dat_dma_pvld;
  assign _0774_ = dat_rdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:742" *) pfifo0_sel;
  assign pfifo0_rd_prdy = _0774_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:742" *) cmd2dat_dma_pvld;
  assign _0775_ = dat_rdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:743" *) pfifo1_sel;
  assign pfifo1_rd_prdy = _0775_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:743" *) cmd2dat_dma_pvld;
  assign _0776_ = dat_rdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:744" *) pfifo2_sel;
  assign pfifo2_rd_prdy = _0776_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:744" *) cmd2dat_dma_pvld;
  assign _0777_ = dat_rdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:745" *) pfifo3_sel;
  assign pfifo3_rd_prdy = _0777_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:745" *) cmd2dat_dma_pvld;
  assign _0778_ = dat_rdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:746" *) sfifo0_sel;
  assign sfifo0_rd_prdy = _0778_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:746" *) cmd2dat_dma_pvld;
  assign _0779_ = dat_rdy & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:747" *) sfifo1_sel;
  assign sfifo1_rd_prdy = _0779_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:747" *) cmd2dat_dma_pvld;
  assign pfifo0_rd_data = { pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel, pfifo0_sel } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:749" *) pfifo0_rd_pd;
  assign pfifo1_rd_data = { pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel, pfifo1_sel } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:750" *) pfifo1_rd_pd;
  assign pfifo2_rd_data = { pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel, pfifo2_sel } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:751" *) pfifo2_rd_pd;
  assign pfifo3_rd_data = { pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel, pfifo3_sel } & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:752" *) pfifo3_rd_pd;
  assign _0868_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1117_;
  assign _0869_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0932_;
  assign _0870_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1118_;
  assign _0871_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0933_;
  assign _0872_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1119_;
  assign _0873_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0934_;
  assign _0874_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1120_;
  assign _0875_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0935_;
  assign _0876_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1121_;
  assign _0877_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0936_;
  assign _0878_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1122_;
  assign _0879_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0937_;
  assign _0880_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1123_;
  assign _0881_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0938_;
  assign _0882_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1124_;
  assign _0883_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0939_;
  assign _0884_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1125_;
  assign _0885_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0940_;
  assign _0886_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1126_;
  assign _0887_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0941_;
  assign _0888_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1127_;
  assign _0889_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0942_;
  assign _0890_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1128_;
  assign _0891_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0943_;
  assign _0892_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1129_;
  assign _0893_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0944_;
  assign _0894_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1130_;
  assign _0895_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0945_;
  assign _0896_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1131_;
  assign _0897_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0946_;
  assign _0898_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1132_;
  assign _0899_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0947_;
  assign _0900_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1133_;
  assign _0901_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0948_;
  assign _0902_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1134_;
  assign _0903_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0949_;
  assign _0904_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1135_;
  assign _0905_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0950_;
  assign _0906_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1136_;
  assign _0907_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0951_;
  assign _0908_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1137_;
  assign _0909_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0952_;
  assign _0910_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1138_;
  assign _0911_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0953_;
  assign _0912_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1139_;
  assign _0913_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0954_;
  assign _0914_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1140_;
  assign _0915_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0955_;
  assign _0916_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1141_;
  assign _0917_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0956_;
  assign _0918_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1142_;
  assign _0919_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0957_;
  assign _0920_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1143_;
  assign _0921_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0958_;
  assign _0922_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1144_;
  assign _0923_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0959_;
  assign _0924_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1145_;
  assign _0925_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0960_;
  assign _0926_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1146_;
  assign _0927_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0961_;
  assign _0928_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1147_;
  assign _0929_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0962_;
  assign _0930_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _1148_;
  assign _0931_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) _0963_;
  assign cfg_di_int8 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:571" *) reg2dp_in_precision;
  assign cfg_di_int16 = reg2dp_in_precision == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:572" *) 1'b1;
  assign cfg_di_fp16 = reg2dp_in_precision == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:573" *) 2'b10;
  assign cfg_do_int8 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:575" *) reg2dp_proc_precision;
  assign _0996_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:578" *) reg2dp_width;
  assign _0997_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:578" *) reg2dp_height;
  assign is_last_beat = beat_cnt == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:600" *) size_of_beat;
  assign _0998_ = pfifo0_rd_data[14:10] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:603" *) 5'b11111;
  assign _0999_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:603" *) pfifo0_rd_data[9:0];
  assign _1000_ = pfifo0_rd_data[30:26] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:604" *) 5'b11111;
  assign _1001_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:604" *) pfifo0_rd_data[25:16];
  assign _1002_ = pfifo0_rd_data[46:42] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:605" *) 5'b11111;
  assign _1003_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:605" *) pfifo0_rd_data[41:32];
  assign _1004_ = pfifo0_rd_data[62:58] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:606" *) 5'b11111;
  assign _1005_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:606" *) pfifo0_rd_data[57:48];
  assign _1006_ = pfifo0_rd_data[78:74] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:607" *) 5'b11111;
  assign _1007_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:607" *) pfifo0_rd_data[73:64];
  assign _1008_ = pfifo0_rd_data[94:90] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:608" *) 5'b11111;
  assign _1009_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:608" *) pfifo0_rd_data[89:80];
  assign _1010_ = pfifo0_rd_data[110:106] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:609" *) 5'b11111;
  assign _1011_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:609" *) pfifo0_rd_data[105:96];
  assign _1012_ = pfifo0_rd_data[126:122] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:610" *) 5'b11111;
  assign _1013_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:610" *) pfifo0_rd_data[121:112];
  assign _1014_ = pfifo1_rd_data[14:10] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:611" *) 5'b11111;
  assign _1015_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:611" *) pfifo1_rd_data[9:0];
  assign _1016_ = pfifo1_rd_data[30:26] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:612" *) 5'b11111;
  assign _1017_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:612" *) pfifo1_rd_data[25:16];
  assign _1018_ = pfifo1_rd_data[46:42] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:613" *) 5'b11111;
  assign _1019_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:613" *) pfifo1_rd_data[41:32];
  assign _1020_ = pfifo1_rd_data[62:58] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:614" *) 5'b11111;
  assign _1021_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:614" *) pfifo1_rd_data[57:48];
  assign _1022_ = pfifo1_rd_data[78:74] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:615" *) 5'b11111;
  assign _1023_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:615" *) pfifo1_rd_data[73:64];
  assign _1024_ = pfifo1_rd_data[94:90] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:616" *) 5'b11111;
  assign _1025_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:616" *) pfifo1_rd_data[89:80];
  assign _1026_ = pfifo1_rd_data[110:106] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:617" *) 5'b11111;
  assign _1027_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:617" *) pfifo1_rd_data[105:96];
  assign _1028_ = pfifo1_rd_data[126:122] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:618" *) 5'b11111;
  assign _1029_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:618" *) pfifo1_rd_data[121:112];
  assign _1030_ = pfifo2_rd_data[14:10] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:619" *) 5'b11111;
  assign _1031_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:619" *) pfifo2_rd_data[9:0];
  assign _1032_ = pfifo2_rd_data[30:26] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:620" *) 5'b11111;
  assign _1033_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:620" *) pfifo2_rd_data[25:16];
  assign _1034_ = pfifo2_rd_data[46:42] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:621" *) 5'b11111;
  assign _1035_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:621" *) pfifo2_rd_data[41:32];
  assign _1036_ = pfifo2_rd_data[62:58] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:622" *) 5'b11111;
  assign _1037_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:622" *) pfifo2_rd_data[57:48];
  assign _1038_ = pfifo2_rd_data[78:74] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:623" *) 5'b11111;
  assign _1039_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:623" *) pfifo2_rd_data[73:64];
  assign _1040_ = pfifo2_rd_data[94:90] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:624" *) 5'b11111;
  assign _1041_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:624" *) pfifo2_rd_data[89:80];
  assign _1042_ = pfifo2_rd_data[110:106] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:625" *) 5'b11111;
  assign _1043_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:625" *) pfifo2_rd_data[105:96];
  assign _1044_ = pfifo2_rd_data[126:122] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:626" *) 5'b11111;
  assign _1045_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:626" *) pfifo2_rd_data[121:112];
  assign _1046_ = pfifo3_rd_data[14:10] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:627" *) 5'b11111;
  assign _1047_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:627" *) pfifo3_rd_data[9:0];
  assign _1048_ = pfifo3_rd_data[30:26] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:628" *) 5'b11111;
  assign _1049_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:628" *) pfifo3_rd_data[25:16];
  assign _1050_ = pfifo3_rd_data[46:42] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:629" *) 5'b11111;
  assign _1051_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:629" *) pfifo3_rd_data[41:32];
  assign _1052_ = pfifo3_rd_data[62:58] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:630" *) 5'b11111;
  assign _1053_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:630" *) pfifo3_rd_data[57:48];
  assign _1054_ = pfifo3_rd_data[78:74] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:631" *) 5'b11111;
  assign _1055_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:631" *) pfifo3_rd_data[73:64];
  assign _1056_ = pfifo3_rd_data[94:90] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:632" *) 5'b11111;
  assign _1057_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:632" *) pfifo3_rd_data[89:80];
  assign _1058_ = pfifo3_rd_data[110:106] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:633" *) 5'b11111;
  assign _1059_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:633" *) pfifo3_rd_data[105:96];
  assign _1060_ = pfifo3_rd_data[126:122] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:634" *) 5'b11111;
  assign _1061_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:634" *) pfifo3_rd_data[121:112];
  assign mode_norm_pfifo0_sel_16 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:712" *) beat_cnt[0];
  assign mode_norm_pfifo0_sel_8 = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:716" *) beat_cnt[1:0];
  assign mode_norm_pfifo1_sel_8 = beat_cnt[1:0] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:717" *) 1'b1;
  assign mode_norm_pfifo2_sel_8 = beat_cnt[1:0] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:718" *) 2'b10;
  assign mode_norm_pfifo3_sel_8 = beat_cnt[1:0] == (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:719" *) 2'b11;
  assign pfifo0_data_byte0_is_inf = _0998_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:603" *) _0999_;
  assign pfifo0_data_byte1_is_inf = _1000_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:604" *) _1001_;
  assign pfifo0_data_byte2_is_inf = _1002_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:605" *) _1003_;
  assign pfifo0_data_byte3_is_inf = _1004_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:606" *) _1005_;
  assign pfifo0_data_byte4_is_inf = _1006_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:607" *) _1007_;
  assign pfifo0_data_byte5_is_inf = _1008_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:608" *) _1009_;
  assign pfifo0_data_byte6_is_inf = _1010_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:609" *) _1011_;
  assign pfifo0_data_byte7_is_inf = _1012_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:610" *) _1013_;
  assign pfifo1_data_byte0_is_inf = _1014_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:611" *) _1015_;
  assign pfifo1_data_byte1_is_inf = _1016_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:612" *) _1017_;
  assign pfifo1_data_byte2_is_inf = _1018_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:613" *) _1019_;
  assign pfifo1_data_byte3_is_inf = _1020_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:614" *) _1021_;
  assign pfifo1_data_byte4_is_inf = _1022_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:615" *) _1023_;
  assign pfifo1_data_byte5_is_inf = _1024_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:616" *) _1025_;
  assign pfifo1_data_byte6_is_inf = _1026_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:617" *) _1027_;
  assign pfifo1_data_byte7_is_inf = _1028_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:618" *) _1029_;
  assign pfifo2_data_byte0_is_inf = _1030_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:619" *) _1031_;
  assign pfifo2_data_byte1_is_inf = _1032_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:620" *) _1033_;
  assign pfifo2_data_byte2_is_inf = _1034_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:621" *) _1035_;
  assign pfifo2_data_byte3_is_inf = _1036_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:622" *) _1037_;
  assign pfifo2_data_byte4_is_inf = _1038_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:623" *) _1039_;
  assign pfifo2_data_byte5_is_inf = _1040_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:624" *) _1041_;
  assign pfifo2_data_byte6_is_inf = _1042_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:625" *) _1043_;
  assign pfifo2_data_byte7_is_inf = _1044_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:626" *) _1045_;
  assign pfifo3_data_byte0_is_inf = _1046_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:627" *) _1047_;
  assign pfifo3_data_byte1_is_inf = _1048_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:628" *) _1049_;
  assign pfifo3_data_byte2_is_inf = _1050_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:629" *) _1051_;
  assign pfifo3_data_byte3_is_inf = _1052_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:630" *) _1053_;
  assign pfifo3_data_byte4_is_inf = _1054_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:631" *) _1055_;
  assign pfifo3_data_byte5_is_inf = _1056_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:632" *) _1057_;
  assign pfifo3_data_byte6_is_inf = _1058_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:633" *) _1059_;
  assign pfifo3_data_byte7_is_inf = _1060_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:634" *) _1061_;
  assign _1062_ = cfg_di_fp16 && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:643" *) reg2dp_perf_nan_inf_count_en;
  assign pfifo0_data_byte0_is_nan = _0998_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:657" *) _1067_;
  assign pfifo0_data_byte1_is_nan = _1000_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:658" *) _1068_;
  assign pfifo0_data_byte2_is_nan = _1002_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:659" *) _1069_;
  assign pfifo0_data_byte3_is_nan = _1004_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:660" *) _1070_;
  assign pfifo0_data_byte4_is_nan = _1006_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:661" *) _1071_;
  assign pfifo0_data_byte5_is_nan = _1008_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:662" *) _1072_;
  assign pfifo0_data_byte6_is_nan = _1010_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:663" *) _1073_;
  assign pfifo0_data_byte7_is_nan = _1012_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:664" *) _1074_;
  assign pfifo1_data_byte0_is_nan = _1014_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:665" *) _1075_;
  assign pfifo1_data_byte1_is_nan = _1016_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:666" *) _1076_;
  assign pfifo1_data_byte2_is_nan = _1018_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:667" *) _1077_;
  assign pfifo1_data_byte3_is_nan = _1020_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:668" *) _1078_;
  assign pfifo1_data_byte4_is_nan = _1022_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:669" *) _1079_;
  assign pfifo1_data_byte5_is_nan = _1024_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:670" *) _1080_;
  assign pfifo1_data_byte6_is_nan = _1026_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:671" *) _1081_;
  assign pfifo1_data_byte7_is_nan = _1028_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:672" *) _1082_;
  assign pfifo2_data_byte0_is_nan = _1030_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:673" *) _1083_;
  assign pfifo2_data_byte1_is_nan = _1032_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:674" *) _1084_;
  assign pfifo2_data_byte2_is_nan = _1034_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:675" *) _1085_;
  assign pfifo2_data_byte3_is_nan = _1036_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:676" *) _1086_;
  assign pfifo2_data_byte4_is_nan = _1038_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:677" *) _1087_;
  assign pfifo2_data_byte5_is_nan = _1040_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:678" *) _1088_;
  assign pfifo2_data_byte6_is_nan = _1042_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:679" *) _1089_;
  assign pfifo2_data_byte7_is_nan = _1044_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:680" *) _1090_;
  assign pfifo3_data_byte0_is_nan = _1046_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:681" *) _1091_;
  assign pfifo3_data_byte1_is_nan = _1048_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:682" *) _1092_;
  assign pfifo3_data_byte2_is_nan = _1050_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:683" *) _1093_;
  assign pfifo3_data_byte3_is_nan = _1052_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:684" *) _1094_;
  assign pfifo3_data_byte4_is_nan = _1054_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:685" *) _1095_;
  assign pfifo3_data_byte5_is_nan = _1056_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:686" *) _1096_;
  assign pfifo3_data_byte6_is_nan = _1058_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:687" *) _1097_;
  assign pfifo3_data_byte7_is_nan = _1060_ && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:688" *) _1098_;
  assign _1063_ = cfg_mode_16to8 && (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:730" *) _1064_;
  assign _1064_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:730" *) cfg_mode_1x1_pack;
  assign _1065_ = inf_input_cnt_nxt_c || (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:647" *) _1115_;
  assign _1066_ = nan_input_cnt_nxt_c || (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:701" *) _1116_;
  assign _1067_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:657" *) pfifo0_rd_data[9:0];
  assign _1068_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:658" *) pfifo0_rd_data[25:16];
  assign _1069_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:659" *) pfifo0_rd_data[41:32];
  assign _1070_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:660" *) pfifo0_rd_data[57:48];
  assign _1071_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:661" *) pfifo0_rd_data[73:64];
  assign _1072_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:662" *) pfifo0_rd_data[89:80];
  assign _1073_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:663" *) pfifo0_rd_data[105:96];
  assign _1074_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:664" *) pfifo0_rd_data[121:112];
  assign _1075_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:665" *) pfifo1_rd_data[9:0];
  assign _1076_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:666" *) pfifo1_rd_data[25:16];
  assign _1077_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:667" *) pfifo1_rd_data[41:32];
  assign _1078_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:668" *) pfifo1_rd_data[57:48];
  assign _1079_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:669" *) pfifo1_rd_data[73:64];
  assign _1080_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:670" *) pfifo1_rd_data[89:80];
  assign _1081_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:671" *) pfifo1_rd_data[105:96];
  assign _1082_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:672" *) pfifo1_rd_data[121:112];
  assign _1083_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:673" *) pfifo2_rd_data[9:0];
  assign _1084_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:674" *) pfifo2_rd_data[25:16];
  assign _1085_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:675" *) pfifo2_rd_data[41:32];
  assign _1086_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:676" *) pfifo2_rd_data[57:48];
  assign _1087_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:677" *) pfifo2_rd_data[73:64];
  assign _1088_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:678" *) pfifo2_rd_data[89:80];
  assign _1089_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:679" *) pfifo2_rd_data[105:96];
  assign _1090_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:680" *) pfifo2_rd_data[121:112];
  assign _1091_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:681" *) pfifo3_rd_data[9:0];
  assign _1092_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:682" *) pfifo3_rd_data[25:16];
  assign _1093_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:683" *) pfifo3_rd_data[41:32];
  assign _1094_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:684" *) pfifo3_rd_data[57:48];
  assign _1095_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:685" *) pfifo3_rd_data[73:64];
  assign _1096_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:686" *) pfifo3_rd_data[89:80];
  assign _1097_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:687" *) pfifo3_rd_data[105:96];
  assign _1098_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:688" *) pfifo3_rd_data[121:112];
  assign _0782_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[9], _1149_, _1181_, _1213_, _1245_, _1277_, _1309_, _1341_, _1373_, _0932_ };
  assign _0783_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[25], _1150_, _1182_, _1214_, _1246_, _1278_, _1310_, _1342_, _1374_, _0933_ };
  assign _0784_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[41], _1151_, _1183_, _1215_, _1247_, _1279_, _1311_, _1343_, _1375_, _0934_ };
  assign _0785_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[57], _1152_, _1184_, _1216_, _1248_, _1280_, _1312_, _1344_, _1376_, _0935_ };
  assign _0786_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[73], _1153_, _1185_, _1217_, _1249_, _1281_, _1313_, _1345_, _1377_, _0936_ };
  assign _0787_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[89], _1154_, _1186_, _1218_, _1250_, _1282_, _1314_, _1346_, _1378_, _0937_ };
  assign _0788_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[105], _1155_, _1187_, _1219_, _1251_, _1283_, _1315_, _1347_, _1379_, _0938_ };
  assign _0789_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo0_rd_data[121], _1156_, _1188_, _1220_, _1252_, _1284_, _1316_, _1348_, _1380_, _0939_ };
  assign _0790_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[9], _1157_, _1189_, _1221_, _1253_, _1285_, _1317_, _1349_, _1381_, _0940_ };
  assign _0791_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[25], _1158_, _1190_, _1222_, _1254_, _1286_, _1318_, _1350_, _1382_, _0941_ };
  assign _0792_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[41], _1159_, _1191_, _1223_, _1255_, _1287_, _1319_, _1351_, _1383_, _0942_ };
  assign _0793_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[57], _1160_, _1192_, _1224_, _1256_, _1288_, _1320_, _1352_, _1384_, _0943_ };
  assign _0794_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[73], _1161_, _1193_, _1225_, _1257_, _1289_, _1321_, _1353_, _1385_, _0944_ };
  assign _0795_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[89], _1162_, _1194_, _1226_, _1258_, _1290_, _1322_, _1354_, _1386_, _0945_ };
  assign _0796_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[105], _1163_, _1195_, _1227_, _1259_, _1291_, _1323_, _1355_, _1387_, _0946_ };
  assign _0797_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo1_rd_data[121], _1164_, _1196_, _1228_, _1260_, _1292_, _1324_, _1356_, _1388_, _0947_ };
  assign _0798_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[9], _1165_, _1197_, _1229_, _1261_, _1293_, _1325_, _1357_, _1389_, _0948_ };
  assign _0799_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[25], _1166_, _1198_, _1230_, _1262_, _1294_, _1326_, _1358_, _1390_, _0949_ };
  assign _0800_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[41], _1167_, _1199_, _1231_, _1263_, _1295_, _1327_, _1359_, _1391_, _0950_ };
  assign _0801_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[57], _1168_, _1200_, _1232_, _1264_, _1296_, _1328_, _1360_, _1392_, _0951_ };
  assign _0802_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[73], _1169_, _1201_, _1233_, _1265_, _1297_, _1329_, _1361_, _1393_, _0952_ };
  assign _0803_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[89], _1170_, _1202_, _1234_, _1266_, _1298_, _1330_, _1362_, _1394_, _0953_ };
  assign _0804_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[105], _1171_, _1203_, _1235_, _1267_, _1299_, _1331_, _1363_, _1395_, _0954_ };
  assign _0805_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo2_rd_data[121], _1172_, _1204_, _1236_, _1268_, _1300_, _1332_, _1364_, _1396_, _0955_ };
  assign _0806_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[9], _1173_, _1205_, _1237_, _1269_, _1301_, _1333_, _1365_, _1397_, _0956_ };
  assign _0807_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[25], _1174_, _1206_, _1238_, _1270_, _1302_, _1334_, _1366_, _1398_, _0957_ };
  assign _0808_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[41], _1175_, _1207_, _1239_, _1271_, _1303_, _1335_, _1367_, _1399_, _0958_ };
  assign _0809_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[57], _1176_, _1208_, _1240_, _1272_, _1304_, _1336_, _1368_, _1400_, _0959_ };
  assign _0810_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[73], _1177_, _1209_, _1241_, _1273_, _1305_, _1337_, _1369_, _1401_, _0960_ };
  assign _0811_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[89], _1178_, _1210_, _1242_, _1274_, _1306_, _1338_, _1370_, _1402_, _0961_ };
  assign _0812_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[105], _1179_, _1211_, _1243_, _1275_, _1307_, _1339_, _1371_, _1403_, _0962_ };
  assign _0813_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1484" *) { pfifo3_rd_data[121], _1180_, _1212_, _1244_, _1276_, _1308_, _1340_, _1372_, _1404_, _0963_ };
  assign _1099_ = pfifo3_sel | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1156" *) pfifo2_sel;
  assign _1100_ = _1099_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1156" *) pfifo1_sel;
  assign pfifo_sel = _1100_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1156" *) pfifo0_sel;
  assign sfifo_sel = sfifo1_sel | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1157" *) sfifo0_sel;
  assign cfg_di_16 = cfg_di_int16 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:574" *) cfg_di_fp16;
  assign _1101_ = _0768_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) _0769_;
  assign _1102_ = _1101_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) _0770_;
  assign pfifo_vld = _1102_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:737" *) _0771_;
  assign sfifo_vld = _0772_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:738" *) _0773_;
  assign fifo_vld = pfifo_vld | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:739" *) sfifo_vld;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      eg_done <= 1'b0;
    else
      eg_done <= _0129_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      nan_input_cnt <= 32'd0;
    else
      nan_input_cnt <= _0131_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      inf_input_cnt <= 32'd0;
    else
      inf_input_cnt <= _0130_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      beat_cnt <= 14'b00000000000000;
    else
      beat_cnt <= _0128_;
  assign _0323_ = _0125_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[121:112], 13'b0000000000000 };
  assign _0322_ = _0125_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0387_;
  assign _0259_ = _0126_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[121:112] } : _0323_;
  assign _0258_ = _0126_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0322_;
  assign _0194_ = _0124_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0867_[7:0] : _0258_;
  assign _0195_ = _0124_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0843_[22:0] : _0259_;
  assign pfifo3_data_ext_byte7_fp16[22:0] = _0127_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0195_;
  assign pfifo3_data_ext_byte7_fp16[30:23] = _0127_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0194_;
  assign _0321_ = _0121_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[105:96], 13'b0000000000000 };
  assign _0320_ = _0121_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0386_;
  assign _0257_ = _0122_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[105:96] } : _0321_;
  assign _0256_ = _0122_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0320_;
  assign _0192_ = _0120_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0866_[7:0] : _0256_;
  assign _0193_ = _0120_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0842_[22:0] : _0257_;
  assign pfifo3_data_ext_byte6_fp16[22:0] = _0123_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0193_;
  assign pfifo3_data_ext_byte6_fp16[30:23] = _0123_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0192_;
  assign _0319_ = _0117_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[89:80], 13'b0000000000000 };
  assign _0318_ = _0117_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0385_;
  assign _0255_ = _0118_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[89:80] } : _0319_;
  assign _0254_ = _0118_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0318_;
  assign _0190_ = _0116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0865_[7:0] : _0254_;
  assign _0191_ = _0116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0841_[22:0] : _0255_;
  assign pfifo3_data_ext_byte5_fp16[22:0] = _0119_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0191_;
  assign pfifo3_data_ext_byte5_fp16[30:23] = _0119_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0190_;
  assign _0317_ = _0113_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[73:64], 13'b0000000000000 };
  assign _0316_ = _0113_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0384_;
  assign _0253_ = _0114_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[73:64] } : _0317_;
  assign _0252_ = _0114_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0316_;
  assign _0188_ = _0112_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0864_[7:0] : _0252_;
  assign _0189_ = _0112_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0840_[22:0] : _0253_;
  assign pfifo3_data_ext_byte4_fp16[22:0] = _0115_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0189_;
  assign pfifo3_data_ext_byte4_fp16[30:23] = _0115_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0188_;
  assign _0315_ = _0109_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[57:48], 13'b0000000000000 };
  assign _0314_ = _0109_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0383_;
  assign _0251_ = _0110_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[57:48] } : _0315_;
  assign _0250_ = _0110_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0314_;
  assign _0186_ = _0108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1414_[7:0] : _0250_;
  assign _0187_ = _0108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0839_[22:0] : _0251_;
  assign pfifo3_data_ext_byte3_fp16[22:0] = _0111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0187_;
  assign pfifo3_data_ext_byte3_fp16[30:23] = _0111_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0186_;
  assign _0313_ = _0105_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[41:32], 13'b0000000000000 };
  assign _0312_ = _0105_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0382_;
  assign _0249_ = _0106_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[41:32] } : _0313_;
  assign _0248_ = _0106_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0312_;
  assign _0184_ = _0104_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1413_[7:0] : _0248_;
  assign _0185_ = _0104_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0838_[22:0] : _0249_;
  assign pfifo3_data_ext_byte2_fp16[22:0] = _0107_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0185_;
  assign pfifo3_data_ext_byte2_fp16[30:23] = _0107_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0184_;
  assign _0311_ = _0101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[25:16], 13'b0000000000000 };
  assign _0310_ = _0101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0381_;
  assign _0247_ = _0102_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[25:16] } : _0311_;
  assign _0246_ = _0102_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0310_;
  assign _0182_ = _0100_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1412_[7:0] : _0246_;
  assign _0183_ = _0100_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0837_[22:0] : _0247_;
  assign pfifo3_data_ext_byte1_fp16[22:0] = _0103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0183_;
  assign pfifo3_data_ext_byte1_fp16[30:23] = _0103_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0182_;
  assign _0309_ = _0097_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo3_rd_data[9:0], 13'b0000000000000 };
  assign _0308_ = _0097_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0380_;
  assign _0245_ = _0098_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo3_rd_data[9:0] } : _0309_;
  assign _0244_ = _0098_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0308_;
  assign _0180_ = _0096_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1411_[7:0] : _0244_;
  assign _0181_ = _0096_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0836_[22:0] : _0245_;
  assign pfifo3_data_ext_byte0_fp16[22:0] = _0099_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0181_;
  assign pfifo3_data_ext_byte0_fp16[30:23] = _0099_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0180_;
  assign _0307_ = _0093_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[121:112], 13'b0000000000000 };
  assign _0306_ = _0093_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0379_;
  assign _0243_ = _0094_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[121:112] } : _0307_;
  assign _0242_ = _0094_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0306_;
  assign _0178_ = _0092_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0863_[7:0] : _0242_;
  assign _0179_ = _0092_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0835_[22:0] : _0243_;
  assign pfifo2_data_ext_byte7_fp16[22:0] = _0095_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0179_;
  assign pfifo2_data_ext_byte7_fp16[30:23] = _0095_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0178_;
  assign _0305_ = _0089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[105:96], 13'b0000000000000 };
  assign _0304_ = _0089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0378_;
  assign _0241_ = _0090_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[105:96] } : _0305_;
  assign _0240_ = _0090_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0304_;
  assign _0176_ = _0088_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0862_[7:0] : _0240_;
  assign _0177_ = _0088_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0834_[22:0] : _0241_;
  assign pfifo2_data_ext_byte6_fp16[22:0] = _0091_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0177_;
  assign pfifo2_data_ext_byte6_fp16[30:23] = _0091_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0176_;
  assign _0303_ = _0085_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[89:80], 13'b0000000000000 };
  assign _0302_ = _0085_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0377_;
  assign _0239_ = _0086_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[89:80] } : _0303_;
  assign _0238_ = _0086_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0302_;
  assign _0174_ = _0084_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0861_[7:0] : _0238_;
  assign _0175_ = _0084_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0833_[22:0] : _0239_;
  assign pfifo2_data_ext_byte5_fp16[22:0] = _0087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0175_;
  assign pfifo2_data_ext_byte5_fp16[30:23] = _0087_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0174_;
  assign _0301_ = _0081_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[73:64], 13'b0000000000000 };
  assign _0300_ = _0081_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0376_;
  assign _0237_ = _0082_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[73:64] } : _0301_;
  assign _0236_ = _0082_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0300_;
  assign _0172_ = _0080_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1410_[7:0] : _0236_;
  assign _0173_ = _0080_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1406_[22:0] : _0237_;
  assign pfifo2_data_ext_byte4_fp16[22:0] = _0083_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0173_;
  assign pfifo2_data_ext_byte4_fp16[30:23] = _0083_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0172_;
  assign _0299_ = _0077_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[57:48], 13'b0000000000000 };
  assign _0298_ = _0077_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0375_;
  assign _0235_ = _0078_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[57:48] } : _0299_;
  assign _0234_ = _0078_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0298_;
  assign _0170_ = _0076_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0860_[7:0] : _0234_;
  assign _0171_ = _0076_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0832_[22:0] : _0235_;
  assign pfifo2_data_ext_byte3_fp16[22:0] = _0079_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0171_;
  assign pfifo2_data_ext_byte3_fp16[30:23] = _0079_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0170_;
  assign _0297_ = _0073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[41:32], 13'b0000000000000 };
  assign _0296_ = _0073_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0374_;
  assign _0233_ = _0074_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[41:32] } : _0297_;
  assign _0232_ = _0074_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0296_;
  assign _0168_ = _0072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0859_[7:0] : _0232_;
  assign _0169_ = _0072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0831_[22:0] : _0233_;
  assign pfifo2_data_ext_byte2_fp16[22:0] = _0075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0169_;
  assign pfifo2_data_ext_byte2_fp16[30:23] = _0075_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0168_;
  assign _0295_ = _0069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[25:16], 13'b0000000000000 };
  assign _0294_ = _0069_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0373_;
  assign _0231_ = _0070_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[25:16] } : _0295_;
  assign _0230_ = _0070_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0294_;
  assign _0166_ = _0068_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0858_[7:0] : _0230_;
  assign _0167_ = _0068_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0830_[22:0] : _0231_;
  assign pfifo2_data_ext_byte1_fp16[22:0] = _0071_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0167_;
  assign pfifo2_data_ext_byte1_fp16[30:23] = _0071_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0166_;
  assign _0293_ = _0065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo2_rd_data[9:0], 13'b0000000000000 };
  assign _0292_ = _0065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0372_;
  assign _0229_ = _0066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo2_rd_data[9:0] } : _0293_;
  assign _0228_ = _0066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0292_;
  assign _0164_ = _0064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0857_[7:0] : _0228_;
  assign _0165_ = _0064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0829_[22:0] : _0229_;
  assign pfifo2_data_ext_byte0_fp16[22:0] = _0067_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0165_;
  assign pfifo2_data_ext_byte0_fp16[30:23] = _0067_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0164_;
  assign _0291_ = _0061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[121:112], 13'b0000000000000 };
  assign _0290_ = _0061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0371_;
  assign _0227_ = _0062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[121:112] } : _0291_;
  assign _0226_ = _0062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0290_;
  assign _0162_ = _0060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0856_[7:0] : _0226_;
  assign _0163_ = _0060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0828_[22:0] : _0227_;
  assign pfifo1_data_ext_byte7_fp16[22:0] = _0063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0163_;
  assign pfifo1_data_ext_byte7_fp16[30:23] = _0063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0162_;
  assign _0289_ = _0057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[105:96], 13'b0000000000000 };
  assign _0288_ = _0057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0370_;
  assign _0225_ = _0058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[105:96] } : _0289_;
  assign _0224_ = _0058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0288_;
  assign _0160_ = _0056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0855_[7:0] : _0224_;
  assign _0161_ = _0056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0827_[22:0] : _0225_;
  assign pfifo1_data_ext_byte6_fp16[22:0] = _0059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0161_;
  assign pfifo1_data_ext_byte6_fp16[30:23] = _0059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0160_;
  assign _0287_ = _0053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[89:80], 13'b0000000000000 };
  assign _0286_ = _0053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0369_;
  assign _0223_ = _0054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[89:80] } : _0287_;
  assign _0222_ = _0054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0286_;
  assign _0158_ = _0052_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0854_[7:0] : _0222_;
  assign _0159_ = _0052_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0826_[22:0] : _0223_;
  assign pfifo1_data_ext_byte5_fp16[22:0] = _0055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0159_;
  assign pfifo1_data_ext_byte5_fp16[30:23] = _0055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0158_;
  assign _0285_ = _0049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[73:64], 13'b0000000000000 };
  assign _0284_ = _0049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0368_;
  assign _0221_ = _0050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[73:64] } : _0285_;
  assign _0220_ = _0050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0284_;
  assign _0156_ = _0048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0853_[7:0] : _0220_;
  assign _0157_ = _0048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0825_[22:0] : _0221_;
  assign pfifo1_data_ext_byte4_fp16[22:0] = _0051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0157_;
  assign pfifo1_data_ext_byte4_fp16[30:23] = _0051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0156_;
  assign _0283_ = _0045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[57:48], 13'b0000000000000 };
  assign _0282_ = _0045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0367_;
  assign _0219_ = _0046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[57:48] } : _0283_;
  assign _0218_ = _0046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0282_;
  assign _0154_ = _0044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1409_[7:0] : _0218_;
  assign _0155_ = _0044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0824_[22:0] : _0219_;
  assign pfifo1_data_ext_byte3_fp16[22:0] = _0047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0155_;
  assign pfifo1_data_ext_byte3_fp16[30:23] = _0047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0154_;
  assign _0281_ = _0041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[41:32], 13'b0000000000000 };
  assign _0280_ = _0041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0366_;
  assign _0217_ = _0042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[41:32] } : _0281_;
  assign _0216_ = _0042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0280_;
  assign _0152_ = _0040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1408_[7:0] : _0216_;
  assign _0153_ = _0040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0823_[22:0] : _0217_;
  assign pfifo1_data_ext_byte2_fp16[22:0] = _0043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0153_;
  assign pfifo1_data_ext_byte2_fp16[30:23] = _0043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0152_;
  assign _0279_ = _0037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[25:16], 13'b0000000000000 };
  assign _0278_ = _0037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0365_;
  assign _0215_ = _0038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[25:16] } : _0279_;
  assign _0214_ = _0038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0278_;
  assign _0150_ = _0036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0852_[7:0] : _0214_;
  assign _0151_ = _0036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0822_[22:0] : _0215_;
  assign pfifo1_data_ext_byte1_fp16[22:0] = _0039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0151_;
  assign pfifo1_data_ext_byte1_fp16[30:23] = _0039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0150_;
  assign _0277_ = _0033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo1_rd_data[9:0], 13'b0000000000000 };
  assign _0276_ = _0033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0364_;
  assign _0213_ = _0034_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo1_rd_data[9:0] } : _0277_;
  assign _0212_ = _0034_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0276_;
  assign _0148_ = _0032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0851_[7:0] : _0212_;
  assign _0149_ = _0032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0821_[22:0] : _0213_;
  assign pfifo1_data_ext_byte0_fp16[22:0] = _0035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0149_;
  assign pfifo1_data_ext_byte0_fp16[30:23] = _0035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0148_;
  assign _0275_ = _0029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[121:112], 13'b0000000000000 };
  assign _0274_ = _0029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0363_;
  assign _0211_ = _0030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[121:112] } : _0275_;
  assign _0210_ = _0030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0274_;
  assign _0146_ = _0028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0850_[7:0] : _0210_;
  assign _0147_ = _0028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0820_[22:0] : _0211_;
  assign pfifo0_data_ext_byte7_fp16[22:0] = _0031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0147_;
  assign pfifo0_data_ext_byte7_fp16[30:23] = _0031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0146_;
  assign _0273_ = _0025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[105:96], 13'b0000000000000 };
  assign _0272_ = _0025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0362_;
  assign _0209_ = _0026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[105:96] } : _0273_;
  assign _0208_ = _0026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0272_;
  assign _0144_ = _0024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0849_[7:0] : _0208_;
  assign _0145_ = _0024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0819_[22:0] : _0209_;
  assign pfifo0_data_ext_byte6_fp16[22:0] = _0027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0145_;
  assign pfifo0_data_ext_byte6_fp16[30:23] = _0027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0144_;
  assign _0271_ = _0021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[89:80], 13'b0000000000000 };
  assign _0270_ = _0021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0361_;
  assign _0207_ = _0022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[89:80] } : _0271_;
  assign _0206_ = _0022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0270_;
  assign _0142_ = _0020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0848_[7:0] : _0206_;
  assign _0143_ = _0020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0818_[22:0] : _0207_;
  assign pfifo0_data_ext_byte5_fp16[22:0] = _0023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0143_;
  assign pfifo0_data_ext_byte5_fp16[30:23] = _0023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0142_;
  assign _0269_ = _0017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[73:64], 13'b0000000000000 };
  assign _0268_ = _0017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0360_;
  assign _0205_ = _0018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[73:64] } : _0269_;
  assign _0204_ = _0018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0268_;
  assign _0140_ = _0016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1407_[7:0] : _0204_;
  assign _0141_ = _0016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _1405_[22:0] : _0205_;
  assign pfifo0_data_ext_byte4_fp16[22:0] = _0019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0141_;
  assign pfifo0_data_ext_byte4_fp16[30:23] = _0019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0140_;
  assign _0267_ = _0013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[57:48], 13'b0000000000000 };
  assign _0266_ = _0013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0359_;
  assign _0203_ = _0014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[57:48] } : _0267_;
  assign _0202_ = _0014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0266_;
  assign _0138_ = _0012_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0847_[7:0] : _0202_;
  assign _0139_ = _0012_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0817_[22:0] : _0203_;
  assign pfifo0_data_ext_byte3_fp16[22:0] = _0015_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0139_;
  assign pfifo0_data_ext_byte3_fp16[30:23] = _0015_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0138_;
  assign _0265_ = _0009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[41:32], 13'b0000000000000 };
  assign _0264_ = _0009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0358_;
  assign _0201_ = _0010_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[41:32] } : _0265_;
  assign _0200_ = _0010_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0264_;
  assign _0136_ = _0008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0846_[7:0] : _0200_;
  assign _0137_ = _0008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0816_[22:0] : _0201_;
  assign pfifo0_data_ext_byte2_fp16[22:0] = _0011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0137_;
  assign pfifo0_data_ext_byte2_fp16[30:23] = _0011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0136_;
  assign _0263_ = _0005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[25:16], 13'b0000000000000 };
  assign _0262_ = _0005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0357_;
  assign _0199_ = _0006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[25:16] } : _0263_;
  assign _0198_ = _0006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0262_;
  assign _0134_ = _0004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0845_[7:0] : _0198_;
  assign _0135_ = _0004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0815_[22:0] : _0199_;
  assign pfifo0_data_ext_byte1_fp16[22:0] = _0007_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0135_;
  assign pfifo0_data_ext_byte1_fp16[30:23] = _0007_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0134_;
  assign _0261_ = _0001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 23'b11111111111111111111111 : { pfifo0_rd_data[9:0], 13'b0000000000000 };
  assign _0260_ = _0001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1455" *) 8'b11111110 : _0356_;
  assign _0197_ = _0002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) { 13'b0000000000000, pfifo0_rd_data[9:0] } : _0261_;
  assign _0196_ = _0002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1452" *) 8'b11111111 : _0260_;
  assign _0132_ = _0000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0844_[7:0] : _0196_;
  assign _0133_ = _0000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1445" *) _0814_[22:0] : _0197_;
  assign pfifo0_data_ext_byte0_fp16[22:0] = _0003_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 23'b00000000000000000000000 : _0133_;
  assign pfifo0_data_ext_byte0_fp16[30:23] = _0003_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1442" *) 8'b00000000 : _0132_;
  assign _1103_ = sfifo1_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1148|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1146" *) { sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16, sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16, sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16, sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16, sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16, sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[334:319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[302:287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[270:255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[238:223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[206:191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[174:159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[142:127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[110:95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[78:63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[46:31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[14:0] } : 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign sfifo_data = sfifo0_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1147|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1146" *) { sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255:239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239:223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223:207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207:191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191:175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175:159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159:143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143:127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127:111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111:95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95:79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79:63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63:47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47:31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31:15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15:0] } : _1103_;
  assign _1104_ = pfifo2_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1131|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1129" *) { pfifo3_rd_data[127], pfifo3_data_ext_byte7_16[30:0], pfifo3_rd_data[111], pfifo3_data_ext_byte6_16[30:0], pfifo3_rd_data[95], pfifo3_data_ext_byte5_16[30:0], pfifo3_rd_data[79], pfifo3_data_ext_byte4_16[30:0], pfifo3_rd_data[63], pfifo3_data_ext_byte3_16[30:0], pfifo3_rd_data[47], pfifo3_data_ext_byte2_16[30:0], pfifo3_rd_data[31], pfifo3_data_ext_byte1_16[30:0], pfifo3_rd_data[15], pfifo3_data_ext_byte0_16[30:0], pfifo2_rd_data[127], pfifo2_data_ext_byte7_16[30:0], pfifo2_rd_data[111], pfifo2_data_ext_byte6_16[30:0], pfifo2_rd_data[95], pfifo2_data_ext_byte5_16[30:0], pfifo2_rd_data[79], pfifo2_data_ext_byte4_16[30:0], pfifo2_rd_data[63], pfifo2_data_ext_byte3_16[30:0], pfifo2_rd_data[47], pfifo2_data_ext_byte2_16[30:0], pfifo2_rd_data[31], pfifo2_data_ext_byte1_16[30:0], pfifo2_rd_data[15], pfifo2_data_ext_byte0_16[30:0] } : 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign pfifo_data_16 = pfifo0_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1130|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1129" *) { pfifo1_rd_data[127], pfifo1_data_ext_byte7_16[30:0], pfifo1_rd_data[111], pfifo1_data_ext_byte6_16[30:0], pfifo1_rd_data[95], pfifo1_data_ext_byte5_16[30:0], pfifo1_rd_data[79], pfifo1_data_ext_byte4_16[30:0], pfifo1_rd_data[63], pfifo1_data_ext_byte3_16[30:0], pfifo1_rd_data[47], pfifo1_data_ext_byte2_16[30:0], pfifo1_rd_data[31], pfifo1_data_ext_byte1_16[30:0], pfifo1_rd_data[15], pfifo1_data_ext_byte0_16[30:0], pfifo0_rd_data[127], pfifo0_data_ext_byte7_16[30:0], pfifo0_rd_data[111], pfifo0_data_ext_byte6_16[30:0], pfifo0_rd_data[95], pfifo0_data_ext_byte5_16[30:0], pfifo0_rd_data[79], pfifo0_data_ext_byte4_16[30:0], pfifo0_rd_data[63], pfifo0_data_ext_byte3_16[30:0], pfifo0_rd_data[47], pfifo0_data_ext_byte2_16[30:0], pfifo0_rd_data[31], pfifo0_data_ext_byte1_16[30:0], pfifo0_rd_data[15], pfifo0_data_ext_byte0_16[30:0] } : _1104_;
  assign _1105_ = pfifo3_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1115|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1111" *) { pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127:119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119:111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111:103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103:95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95:87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87:79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79:71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71:63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63:55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55:47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47:39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39:31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31:23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23:15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15:7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7:0] } : 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _1106_ = pfifo2_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1114|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1111" *) { pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127:119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119:111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111:103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103:95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95:87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87:79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79:71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71:63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63:55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55:47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47:39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39:31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31:23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23:15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15:7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7:0] } : _1105_;
  assign _1107_ = pfifo1_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1113|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1111" *) { pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127:119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119:111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111:103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103:95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95:87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87:79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79:71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71:63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63:55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55:47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47:39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39:31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31:23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23:15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15:7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7:0] } : _1106_;
  assign pfifo_data_8 = pfifo0_sel ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1112|./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1111" *) { pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127:119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119:111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111:103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103:95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95:87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87:79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79:71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71:63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63:55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55:47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47:39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39:31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31:23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23:15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15:7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7:0] } : _1107_;
  assign _1108_ = _1066_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:701" *) 32'd4294967295 : nan_input_cnt_nxt;
  assign _1109_ = dat_accept ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:700" *) _1108_ : nan_input_cnt;
  assign _1110_ = op_load ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:698" *) 32'd0 : _1109_;
  assign _0131_ = _1062_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:697" *) _1110_ : nan_input_cnt;
  assign _1111_ = _1065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:647" *) 32'd4294967295 : inf_input_cnt_nxt;
  assign _1112_ = dat_accept ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:646" *) _1111_ : inf_input_cnt;
  assign _1113_ = op_load ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:644" *) 32'd0 : _1112_;
  assign _0130_ = _1062_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:643" *) _1113_ : inf_input_cnt;
  assign _1114_ = is_last_beat ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:592" *) 14'b00000000000000 : _0708_;
  assign _0128_ = dat_accept ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:591" *) _1114_ : beat_cnt;
  assign _0964_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[10], pfifo0_rd_data[11], pfifo0_rd_data[12], pfifo0_rd_data[13], pfifo0_rd_data[14] };
  assign _0965_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[26], pfifo0_rd_data[27], pfifo0_rd_data[28], pfifo0_rd_data[29], pfifo0_rd_data[30] };
  assign _0966_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[42], pfifo0_rd_data[43], pfifo0_rd_data[44], pfifo0_rd_data[45], pfifo0_rd_data[46] };
  assign _0967_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[58], pfifo0_rd_data[59], pfifo0_rd_data[60], pfifo0_rd_data[61], pfifo0_rd_data[62] };
  assign _0968_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[74], pfifo0_rd_data[75], pfifo0_rd_data[76], pfifo0_rd_data[77], pfifo0_rd_data[78] };
  assign _0969_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[90], pfifo0_rd_data[91], pfifo0_rd_data[92], pfifo0_rd_data[93], pfifo0_rd_data[94] };
  assign _0970_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[106], pfifo0_rd_data[107], pfifo0_rd_data[108], pfifo0_rd_data[109], pfifo0_rd_data[110] };
  assign _0971_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo0_rd_data[122], pfifo0_rd_data[123], pfifo0_rd_data[124], pfifo0_rd_data[125], pfifo0_rd_data[126] };
  assign _0972_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[10], pfifo1_rd_data[11], pfifo1_rd_data[12], pfifo1_rd_data[13], pfifo1_rd_data[14] };
  assign _0973_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[26], pfifo1_rd_data[27], pfifo1_rd_data[28], pfifo1_rd_data[29], pfifo1_rd_data[30] };
  assign _0974_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[42], pfifo1_rd_data[43], pfifo1_rd_data[44], pfifo1_rd_data[45], pfifo1_rd_data[46] };
  assign _0975_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[58], pfifo1_rd_data[59], pfifo1_rd_data[60], pfifo1_rd_data[61], pfifo1_rd_data[62] };
  assign _0976_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[74], pfifo1_rd_data[75], pfifo1_rd_data[76], pfifo1_rd_data[77], pfifo1_rd_data[78] };
  assign _0977_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[90], pfifo1_rd_data[91], pfifo1_rd_data[92], pfifo1_rd_data[93], pfifo1_rd_data[94] };
  assign _0978_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[106], pfifo1_rd_data[107], pfifo1_rd_data[108], pfifo1_rd_data[109], pfifo1_rd_data[110] };
  assign _0979_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo1_rd_data[122], pfifo1_rd_data[123], pfifo1_rd_data[124], pfifo1_rd_data[125], pfifo1_rd_data[126] };
  assign _0980_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[10], pfifo2_rd_data[11], pfifo2_rd_data[12], pfifo2_rd_data[13], pfifo2_rd_data[14] };
  assign _0981_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[26], pfifo2_rd_data[27], pfifo2_rd_data[28], pfifo2_rd_data[29], pfifo2_rd_data[30] };
  assign _0982_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[42], pfifo2_rd_data[43], pfifo2_rd_data[44], pfifo2_rd_data[45], pfifo2_rd_data[46] };
  assign _0983_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[58], pfifo2_rd_data[59], pfifo2_rd_data[60], pfifo2_rd_data[61], pfifo2_rd_data[62] };
  assign _0984_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[74], pfifo2_rd_data[75], pfifo2_rd_data[76], pfifo2_rd_data[77], pfifo2_rd_data[78] };
  assign _0985_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[90], pfifo2_rd_data[91], pfifo2_rd_data[92], pfifo2_rd_data[93], pfifo2_rd_data[94] };
  assign _0986_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[106], pfifo2_rd_data[107], pfifo2_rd_data[108], pfifo2_rd_data[109], pfifo2_rd_data[110] };
  assign _0987_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo2_rd_data[122], pfifo2_rd_data[123], pfifo2_rd_data[124], pfifo2_rd_data[125], pfifo2_rd_data[126] };
  assign _0988_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[10], pfifo3_rd_data[11], pfifo3_rd_data[12], pfifo3_rd_data[13], pfifo3_rd_data[14] };
  assign _0989_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[26], pfifo3_rd_data[27], pfifo3_rd_data[28], pfifo3_rd_data[29], pfifo3_rd_data[30] };
  assign _0990_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[42], pfifo3_rd_data[43], pfifo3_rd_data[44], pfifo3_rd_data[45], pfifo3_rd_data[46] };
  assign _0991_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[58], pfifo3_rd_data[59], pfifo3_rd_data[60], pfifo3_rd_data[61], pfifo3_rd_data[62] };
  assign _0992_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[74], pfifo3_rd_data[75], pfifo3_rd_data[76], pfifo3_rd_data[77], pfifo3_rd_data[78] };
  assign _0993_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[90], pfifo3_rd_data[91], pfifo3_rd_data[92], pfifo3_rd_data[93], pfifo3_rd_data[94] };
  assign _0994_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[106], pfifo3_rd_data[107], pfifo3_rd_data[108], pfifo3_rd_data[109], pfifo3_rd_data[110] };
  assign _0995_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1439" *) { pfifo3_rd_data[122], pfifo3_rd_data[123], pfifo3_rd_data[124], pfifo3_rd_data[125], pfifo3_rd_data[126] };
  assign _1115_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:647" *) { inf_input_cnt[0], inf_input_cnt[1], inf_input_cnt[2], inf_input_cnt[3], inf_input_cnt[4], inf_input_cnt[5], inf_input_cnt[6], inf_input_cnt[7], inf_input_cnt[8], inf_input_cnt[9], inf_input_cnt[10], inf_input_cnt[11], inf_input_cnt[12], inf_input_cnt[13], inf_input_cnt[14], inf_input_cnt[15], inf_input_cnt[16], inf_input_cnt[17], inf_input_cnt[18], inf_input_cnt[19], inf_input_cnt[20], inf_input_cnt[21], inf_input_cnt[22], inf_input_cnt[23], inf_input_cnt[24], inf_input_cnt[25], inf_input_cnt[26], inf_input_cnt[27], inf_input_cnt[28], inf_input_cnt[29], inf_input_cnt[30], inf_input_cnt[31] };
  assign _1116_ = & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:701" *) { nan_input_cnt[0], nan_input_cnt[1], nan_input_cnt[2], nan_input_cnt[3], nan_input_cnt[4], nan_input_cnt[5], nan_input_cnt[6], nan_input_cnt[7], nan_input_cnt[8], nan_input_cnt[9], nan_input_cnt[10], nan_input_cnt[11], nan_input_cnt[12], nan_input_cnt[13], nan_input_cnt[14], nan_input_cnt[15], nan_input_cnt[16], nan_input_cnt[17], nan_input_cnt[18], nan_input_cnt[19], nan_input_cnt[20], nan_input_cnt[21], nan_input_cnt[22], nan_input_cnt[23], nan_input_cnt[24], nan_input_cnt[25], nan_input_cnt[26], nan_input_cnt[27], nan_input_cnt[28], nan_input_cnt[29], nan_input_cnt[30], nan_input_cnt[31] };
  assign _1117_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[10], pfifo0_rd_data[11], pfifo0_rd_data[12], pfifo0_rd_data[13], pfifo0_rd_data[14] };
  assign _0932_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[0], pfifo0_rd_data[1], pfifo0_rd_data[2], pfifo0_rd_data[3], pfifo0_rd_data[4], pfifo0_rd_data[5], pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1118_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[26], pfifo0_rd_data[27], pfifo0_rd_data[28], pfifo0_rd_data[29], pfifo0_rd_data[30] };
  assign _0933_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[16], pfifo0_rd_data[17], pfifo0_rd_data[18], pfifo0_rd_data[19], pfifo0_rd_data[20], pfifo0_rd_data[21], pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1119_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[42], pfifo0_rd_data[43], pfifo0_rd_data[44], pfifo0_rd_data[45], pfifo0_rd_data[46] };
  assign _0934_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[32], pfifo0_rd_data[33], pfifo0_rd_data[34], pfifo0_rd_data[35], pfifo0_rd_data[36], pfifo0_rd_data[37], pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1120_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[58], pfifo0_rd_data[59], pfifo0_rd_data[60], pfifo0_rd_data[61], pfifo0_rd_data[62] };
  assign _0935_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[48], pfifo0_rd_data[49], pfifo0_rd_data[50], pfifo0_rd_data[51], pfifo0_rd_data[52], pfifo0_rd_data[53], pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1121_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[74], pfifo0_rd_data[75], pfifo0_rd_data[76], pfifo0_rd_data[77], pfifo0_rd_data[78] };
  assign _0936_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[64], pfifo0_rd_data[65], pfifo0_rd_data[66], pfifo0_rd_data[67], pfifo0_rd_data[68], pfifo0_rd_data[69], pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1122_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[90], pfifo0_rd_data[91], pfifo0_rd_data[92], pfifo0_rd_data[93], pfifo0_rd_data[94] };
  assign _0937_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[80], pfifo0_rd_data[81], pfifo0_rd_data[82], pfifo0_rd_data[83], pfifo0_rd_data[84], pfifo0_rd_data[85], pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1123_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[106], pfifo0_rd_data[107], pfifo0_rd_data[108], pfifo0_rd_data[109], pfifo0_rd_data[110] };
  assign _0938_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[96], pfifo0_rd_data[97], pfifo0_rd_data[98], pfifo0_rd_data[99], pfifo0_rd_data[100], pfifo0_rd_data[101], pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1124_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[122], pfifo0_rd_data[123], pfifo0_rd_data[124], pfifo0_rd_data[125], pfifo0_rd_data[126] };
  assign _0939_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo0_rd_data[112], pfifo0_rd_data[113], pfifo0_rd_data[114], pfifo0_rd_data[115], pfifo0_rd_data[116], pfifo0_rd_data[117], pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1125_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[10], pfifo1_rd_data[11], pfifo1_rd_data[12], pfifo1_rd_data[13], pfifo1_rd_data[14] };
  assign _0940_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[0], pfifo1_rd_data[1], pfifo1_rd_data[2], pfifo1_rd_data[3], pfifo1_rd_data[4], pfifo1_rd_data[5], pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1126_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[26], pfifo1_rd_data[27], pfifo1_rd_data[28], pfifo1_rd_data[29], pfifo1_rd_data[30] };
  assign _0941_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[16], pfifo1_rd_data[17], pfifo1_rd_data[18], pfifo1_rd_data[19], pfifo1_rd_data[20], pfifo1_rd_data[21], pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1127_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[42], pfifo1_rd_data[43], pfifo1_rd_data[44], pfifo1_rd_data[45], pfifo1_rd_data[46] };
  assign _0942_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[32], pfifo1_rd_data[33], pfifo1_rd_data[34], pfifo1_rd_data[35], pfifo1_rd_data[36], pfifo1_rd_data[37], pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1128_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[58], pfifo1_rd_data[59], pfifo1_rd_data[60], pfifo1_rd_data[61], pfifo1_rd_data[62] };
  assign _0943_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[48], pfifo1_rd_data[49], pfifo1_rd_data[50], pfifo1_rd_data[51], pfifo1_rd_data[52], pfifo1_rd_data[53], pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1129_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[74], pfifo1_rd_data[75], pfifo1_rd_data[76], pfifo1_rd_data[77], pfifo1_rd_data[78] };
  assign _0944_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[64], pfifo1_rd_data[65], pfifo1_rd_data[66], pfifo1_rd_data[67], pfifo1_rd_data[68], pfifo1_rd_data[69], pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1130_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[90], pfifo1_rd_data[91], pfifo1_rd_data[92], pfifo1_rd_data[93], pfifo1_rd_data[94] };
  assign _0945_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[80], pfifo1_rd_data[81], pfifo1_rd_data[82], pfifo1_rd_data[83], pfifo1_rd_data[84], pfifo1_rd_data[85], pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1131_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[106], pfifo1_rd_data[107], pfifo1_rd_data[108], pfifo1_rd_data[109], pfifo1_rd_data[110] };
  assign _0946_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[96], pfifo1_rd_data[97], pfifo1_rd_data[98], pfifo1_rd_data[99], pfifo1_rd_data[100], pfifo1_rd_data[101], pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1132_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[122], pfifo1_rd_data[123], pfifo1_rd_data[124], pfifo1_rd_data[125], pfifo1_rd_data[126] };
  assign _0947_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo1_rd_data[112], pfifo1_rd_data[113], pfifo1_rd_data[114], pfifo1_rd_data[115], pfifo1_rd_data[116], pfifo1_rd_data[117], pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1133_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[10], pfifo2_rd_data[11], pfifo2_rd_data[12], pfifo2_rd_data[13], pfifo2_rd_data[14] };
  assign _0948_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[0], pfifo2_rd_data[1], pfifo2_rd_data[2], pfifo2_rd_data[3], pfifo2_rd_data[4], pfifo2_rd_data[5], pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1134_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[26], pfifo2_rd_data[27], pfifo2_rd_data[28], pfifo2_rd_data[29], pfifo2_rd_data[30] };
  assign _0949_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[16], pfifo2_rd_data[17], pfifo2_rd_data[18], pfifo2_rd_data[19], pfifo2_rd_data[20], pfifo2_rd_data[21], pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1135_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[42], pfifo2_rd_data[43], pfifo2_rd_data[44], pfifo2_rd_data[45], pfifo2_rd_data[46] };
  assign _0950_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[32], pfifo2_rd_data[33], pfifo2_rd_data[34], pfifo2_rd_data[35], pfifo2_rd_data[36], pfifo2_rd_data[37], pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1136_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[58], pfifo2_rd_data[59], pfifo2_rd_data[60], pfifo2_rd_data[61], pfifo2_rd_data[62] };
  assign _0951_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[48], pfifo2_rd_data[49], pfifo2_rd_data[50], pfifo2_rd_data[51], pfifo2_rd_data[52], pfifo2_rd_data[53], pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1137_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[74], pfifo2_rd_data[75], pfifo2_rd_data[76], pfifo2_rd_data[77], pfifo2_rd_data[78] };
  assign _0952_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[64], pfifo2_rd_data[65], pfifo2_rd_data[66], pfifo2_rd_data[67], pfifo2_rd_data[68], pfifo2_rd_data[69], pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1138_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[90], pfifo2_rd_data[91], pfifo2_rd_data[92], pfifo2_rd_data[93], pfifo2_rd_data[94] };
  assign _0953_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[80], pfifo2_rd_data[81], pfifo2_rd_data[82], pfifo2_rd_data[83], pfifo2_rd_data[84], pfifo2_rd_data[85], pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1139_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[106], pfifo2_rd_data[107], pfifo2_rd_data[108], pfifo2_rd_data[109], pfifo2_rd_data[110] };
  assign _0954_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[96], pfifo2_rd_data[97], pfifo2_rd_data[98], pfifo2_rd_data[99], pfifo2_rd_data[100], pfifo2_rd_data[101], pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1140_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[122], pfifo2_rd_data[123], pfifo2_rd_data[124], pfifo2_rd_data[125], pfifo2_rd_data[126] };
  assign _0955_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo2_rd_data[112], pfifo2_rd_data[113], pfifo2_rd_data[114], pfifo2_rd_data[115], pfifo2_rd_data[116], pfifo2_rd_data[117], pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1141_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[10], pfifo3_rd_data[11], pfifo3_rd_data[12], pfifo3_rd_data[13], pfifo3_rd_data[14] };
  assign _0956_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[0], pfifo3_rd_data[1], pfifo3_rd_data[2], pfifo3_rd_data[3], pfifo3_rd_data[4], pfifo3_rd_data[5], pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1142_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[26], pfifo3_rd_data[27], pfifo3_rd_data[28], pfifo3_rd_data[29], pfifo3_rd_data[30] };
  assign _0957_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[16], pfifo3_rd_data[17], pfifo3_rd_data[18], pfifo3_rd_data[19], pfifo3_rd_data[20], pfifo3_rd_data[21], pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1143_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[42], pfifo3_rd_data[43], pfifo3_rd_data[44], pfifo3_rd_data[45], pfifo3_rd_data[46] };
  assign _0958_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[32], pfifo3_rd_data[33], pfifo3_rd_data[34], pfifo3_rd_data[35], pfifo3_rd_data[36], pfifo3_rd_data[37], pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1144_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[58], pfifo3_rd_data[59], pfifo3_rd_data[60], pfifo3_rd_data[61], pfifo3_rd_data[62] };
  assign _0959_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[48], pfifo3_rd_data[49], pfifo3_rd_data[50], pfifo3_rd_data[51], pfifo3_rd_data[52], pfifo3_rd_data[53], pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1145_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[74], pfifo3_rd_data[75], pfifo3_rd_data[76], pfifo3_rd_data[77], pfifo3_rd_data[78] };
  assign _0960_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[64], pfifo3_rd_data[65], pfifo3_rd_data[66], pfifo3_rd_data[67], pfifo3_rd_data[68], pfifo3_rd_data[69], pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1146_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[90], pfifo3_rd_data[91], pfifo3_rd_data[92], pfifo3_rd_data[93], pfifo3_rd_data[94] };
  assign _0961_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[80], pfifo3_rd_data[81], pfifo3_rd_data[82], pfifo3_rd_data[83], pfifo3_rd_data[84], pfifo3_rd_data[85], pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1147_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[106], pfifo3_rd_data[107], pfifo3_rd_data[108], pfifo3_rd_data[109], pfifo3_rd_data[110] };
  assign _0962_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[96], pfifo3_rd_data[97], pfifo3_rd_data[98], pfifo3_rd_data[99], pfifo3_rd_data[100], pfifo3_rd_data[101], pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1148_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[122], pfifo3_rd_data[123], pfifo3_rd_data[124], pfifo3_rd_data[125], pfifo3_rd_data[126] };
  assign _0963_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1437" *) { pfifo3_rd_data[112], pfifo3_rd_data[113], pfifo3_rd_data[114], pfifo3_rd_data[115], pfifo3_rd_data[116], pfifo3_rd_data[117], pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1149_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1150_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1151_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1152_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1153_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1154_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1155_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1156_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1157_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1158_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1159_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1160_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1161_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1162_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1163_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1164_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1165_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1166_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1167_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1168_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1169_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1170_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1171_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1172_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1173_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1174_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1175_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1176_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1177_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1178_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1179_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1180_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1475" *) { pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1181_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1182_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1183_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1184_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1185_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1186_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1187_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1188_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1189_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1190_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1191_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1192_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1193_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1194_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1195_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1196_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1197_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1198_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1199_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1200_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1201_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1202_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1203_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1204_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1205_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1206_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1207_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1208_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1209_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1210_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1211_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1212_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1476" *) { pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1213_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1214_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1215_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1216_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1217_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1218_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1219_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1220_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1221_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1222_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1223_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1224_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1225_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1226_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1227_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1228_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1229_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1230_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1231_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1232_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1233_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1234_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1235_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1236_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1237_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1238_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1239_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1240_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1241_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1242_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1243_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1244_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1477" *) { pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1245_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[5], pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1246_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[21], pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1247_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[37], pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1248_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[53], pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1249_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[69], pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1250_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[85], pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1251_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[101], pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1252_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo0_rd_data[117], pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1253_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[5], pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1254_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[21], pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1255_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[37], pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1256_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[53], pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1257_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[69], pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1258_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[85], pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1259_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[101], pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1260_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo1_rd_data[117], pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1261_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[5], pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1262_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[21], pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1263_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[37], pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1264_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[53], pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1265_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[69], pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1266_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[85], pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1267_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[101], pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1268_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo2_rd_data[117], pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1269_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[5], pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1270_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[21], pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1271_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[37], pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1272_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[53], pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1273_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[69], pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1274_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[85], pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1275_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[101], pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1276_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1478" *) { pfifo3_rd_data[117], pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1277_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[4], pfifo0_rd_data[5], pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1278_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[20], pfifo0_rd_data[21], pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1279_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[36], pfifo0_rd_data[37], pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1280_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[52], pfifo0_rd_data[53], pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1281_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[68], pfifo0_rd_data[69], pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1282_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[84], pfifo0_rd_data[85], pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1283_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[100], pfifo0_rd_data[101], pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1284_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo0_rd_data[116], pfifo0_rd_data[117], pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1285_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[4], pfifo1_rd_data[5], pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1286_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[20], pfifo1_rd_data[21], pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1287_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[36], pfifo1_rd_data[37], pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1288_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[52], pfifo1_rd_data[53], pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1289_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[68], pfifo1_rd_data[69], pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1290_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[84], pfifo1_rd_data[85], pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1291_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[100], pfifo1_rd_data[101], pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1292_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo1_rd_data[116], pfifo1_rd_data[117], pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1293_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[4], pfifo2_rd_data[5], pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1294_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[20], pfifo2_rd_data[21], pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1295_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[36], pfifo2_rd_data[37], pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1296_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[52], pfifo2_rd_data[53], pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1297_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[68], pfifo2_rd_data[69], pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1298_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[84], pfifo2_rd_data[85], pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1299_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[100], pfifo2_rd_data[101], pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1300_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo2_rd_data[116], pfifo2_rd_data[117], pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1301_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[4], pfifo3_rd_data[5], pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1302_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[20], pfifo3_rd_data[21], pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1303_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[36], pfifo3_rd_data[37], pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1304_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[52], pfifo3_rd_data[53], pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1305_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[68], pfifo3_rd_data[69], pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1306_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[84], pfifo3_rd_data[85], pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1307_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[100], pfifo3_rd_data[101], pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1308_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1479" *) { pfifo3_rd_data[116], pfifo3_rd_data[117], pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1309_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[3], pfifo0_rd_data[4], pfifo0_rd_data[5], pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1310_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[19], pfifo0_rd_data[20], pfifo0_rd_data[21], pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1311_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[35], pfifo0_rd_data[36], pfifo0_rd_data[37], pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1312_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[51], pfifo0_rd_data[52], pfifo0_rd_data[53], pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1313_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[67], pfifo0_rd_data[68], pfifo0_rd_data[69], pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1314_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[83], pfifo0_rd_data[84], pfifo0_rd_data[85], pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1315_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[99], pfifo0_rd_data[100], pfifo0_rd_data[101], pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1316_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo0_rd_data[115], pfifo0_rd_data[116], pfifo0_rd_data[117], pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1317_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[3], pfifo1_rd_data[4], pfifo1_rd_data[5], pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1318_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[19], pfifo1_rd_data[20], pfifo1_rd_data[21], pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1319_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[35], pfifo1_rd_data[36], pfifo1_rd_data[37], pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1320_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[51], pfifo1_rd_data[52], pfifo1_rd_data[53], pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1321_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[67], pfifo1_rd_data[68], pfifo1_rd_data[69], pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1322_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[83], pfifo1_rd_data[84], pfifo1_rd_data[85], pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1323_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[99], pfifo1_rd_data[100], pfifo1_rd_data[101], pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1324_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo1_rd_data[115], pfifo1_rd_data[116], pfifo1_rd_data[117], pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1325_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[3], pfifo2_rd_data[4], pfifo2_rd_data[5], pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1326_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[19], pfifo2_rd_data[20], pfifo2_rd_data[21], pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1327_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[35], pfifo2_rd_data[36], pfifo2_rd_data[37], pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1328_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[51], pfifo2_rd_data[52], pfifo2_rd_data[53], pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1329_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[67], pfifo2_rd_data[68], pfifo2_rd_data[69], pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1330_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[83], pfifo2_rd_data[84], pfifo2_rd_data[85], pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1331_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[99], pfifo2_rd_data[100], pfifo2_rd_data[101], pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1332_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo2_rd_data[115], pfifo2_rd_data[116], pfifo2_rd_data[117], pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1333_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[3], pfifo3_rd_data[4], pfifo3_rd_data[5], pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1334_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[19], pfifo3_rd_data[20], pfifo3_rd_data[21], pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1335_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[35], pfifo3_rd_data[36], pfifo3_rd_data[37], pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1336_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[51], pfifo3_rd_data[52], pfifo3_rd_data[53], pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1337_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[67], pfifo3_rd_data[68], pfifo3_rd_data[69], pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1338_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[83], pfifo3_rd_data[84], pfifo3_rd_data[85], pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1339_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[99], pfifo3_rd_data[100], pfifo3_rd_data[101], pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1340_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1480" *) { pfifo3_rd_data[115], pfifo3_rd_data[116], pfifo3_rd_data[117], pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1341_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[2], pfifo0_rd_data[3], pfifo0_rd_data[4], pfifo0_rd_data[5], pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1342_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[18], pfifo0_rd_data[19], pfifo0_rd_data[20], pfifo0_rd_data[21], pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1343_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[34], pfifo0_rd_data[35], pfifo0_rd_data[36], pfifo0_rd_data[37], pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1344_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[50], pfifo0_rd_data[51], pfifo0_rd_data[52], pfifo0_rd_data[53], pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1345_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[66], pfifo0_rd_data[67], pfifo0_rd_data[68], pfifo0_rd_data[69], pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1346_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[82], pfifo0_rd_data[83], pfifo0_rd_data[84], pfifo0_rd_data[85], pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1347_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[98], pfifo0_rd_data[99], pfifo0_rd_data[100], pfifo0_rd_data[101], pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1348_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo0_rd_data[114], pfifo0_rd_data[115], pfifo0_rd_data[116], pfifo0_rd_data[117], pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1349_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[2], pfifo1_rd_data[3], pfifo1_rd_data[4], pfifo1_rd_data[5], pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1350_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[18], pfifo1_rd_data[19], pfifo1_rd_data[20], pfifo1_rd_data[21], pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1351_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[34], pfifo1_rd_data[35], pfifo1_rd_data[36], pfifo1_rd_data[37], pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1352_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[50], pfifo1_rd_data[51], pfifo1_rd_data[52], pfifo1_rd_data[53], pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1353_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[66], pfifo1_rd_data[67], pfifo1_rd_data[68], pfifo1_rd_data[69], pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1354_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[82], pfifo1_rd_data[83], pfifo1_rd_data[84], pfifo1_rd_data[85], pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1355_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[98], pfifo1_rd_data[99], pfifo1_rd_data[100], pfifo1_rd_data[101], pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1356_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo1_rd_data[114], pfifo1_rd_data[115], pfifo1_rd_data[116], pfifo1_rd_data[117], pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1357_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[2], pfifo2_rd_data[3], pfifo2_rd_data[4], pfifo2_rd_data[5], pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1358_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[18], pfifo2_rd_data[19], pfifo2_rd_data[20], pfifo2_rd_data[21], pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1359_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[34], pfifo2_rd_data[35], pfifo2_rd_data[36], pfifo2_rd_data[37], pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1360_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[50], pfifo2_rd_data[51], pfifo2_rd_data[52], pfifo2_rd_data[53], pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1361_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[66], pfifo2_rd_data[67], pfifo2_rd_data[68], pfifo2_rd_data[69], pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1362_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[82], pfifo2_rd_data[83], pfifo2_rd_data[84], pfifo2_rd_data[85], pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1363_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[98], pfifo2_rd_data[99], pfifo2_rd_data[100], pfifo2_rd_data[101], pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1364_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo2_rd_data[114], pfifo2_rd_data[115], pfifo2_rd_data[116], pfifo2_rd_data[117], pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1365_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[2], pfifo3_rd_data[3], pfifo3_rd_data[4], pfifo3_rd_data[5], pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1366_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[18], pfifo3_rd_data[19], pfifo3_rd_data[20], pfifo3_rd_data[21], pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1367_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[34], pfifo3_rd_data[35], pfifo3_rd_data[36], pfifo3_rd_data[37], pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1368_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[50], pfifo3_rd_data[51], pfifo3_rd_data[52], pfifo3_rd_data[53], pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1369_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[66], pfifo3_rd_data[67], pfifo3_rd_data[68], pfifo3_rd_data[69], pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1370_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[82], pfifo3_rd_data[83], pfifo3_rd_data[84], pfifo3_rd_data[85], pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1371_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[98], pfifo3_rd_data[99], pfifo3_rd_data[100], pfifo3_rd_data[101], pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1372_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1481" *) { pfifo3_rd_data[114], pfifo3_rd_data[115], pfifo3_rd_data[116], pfifo3_rd_data[117], pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _1373_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[1], pfifo0_rd_data[2], pfifo0_rd_data[3], pfifo0_rd_data[4], pfifo0_rd_data[5], pfifo0_rd_data[6], pfifo0_rd_data[7], pfifo0_rd_data[8], pfifo0_rd_data[9] };
  assign _1374_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[17], pfifo0_rd_data[18], pfifo0_rd_data[19], pfifo0_rd_data[20], pfifo0_rd_data[21], pfifo0_rd_data[22], pfifo0_rd_data[23], pfifo0_rd_data[24], pfifo0_rd_data[25] };
  assign _1375_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[33], pfifo0_rd_data[34], pfifo0_rd_data[35], pfifo0_rd_data[36], pfifo0_rd_data[37], pfifo0_rd_data[38], pfifo0_rd_data[39], pfifo0_rd_data[40], pfifo0_rd_data[41] };
  assign _1376_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[49], pfifo0_rd_data[50], pfifo0_rd_data[51], pfifo0_rd_data[52], pfifo0_rd_data[53], pfifo0_rd_data[54], pfifo0_rd_data[55], pfifo0_rd_data[56], pfifo0_rd_data[57] };
  assign _1377_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[65], pfifo0_rd_data[66], pfifo0_rd_data[67], pfifo0_rd_data[68], pfifo0_rd_data[69], pfifo0_rd_data[70], pfifo0_rd_data[71], pfifo0_rd_data[72], pfifo0_rd_data[73] };
  assign _1378_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[81], pfifo0_rd_data[82], pfifo0_rd_data[83], pfifo0_rd_data[84], pfifo0_rd_data[85], pfifo0_rd_data[86], pfifo0_rd_data[87], pfifo0_rd_data[88], pfifo0_rd_data[89] };
  assign _1379_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[97], pfifo0_rd_data[98], pfifo0_rd_data[99], pfifo0_rd_data[100], pfifo0_rd_data[101], pfifo0_rd_data[102], pfifo0_rd_data[103], pfifo0_rd_data[104], pfifo0_rd_data[105] };
  assign _1380_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo0_rd_data[113], pfifo0_rd_data[114], pfifo0_rd_data[115], pfifo0_rd_data[116], pfifo0_rd_data[117], pfifo0_rd_data[118], pfifo0_rd_data[119], pfifo0_rd_data[120], pfifo0_rd_data[121] };
  assign _1381_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[1], pfifo1_rd_data[2], pfifo1_rd_data[3], pfifo1_rd_data[4], pfifo1_rd_data[5], pfifo1_rd_data[6], pfifo1_rd_data[7], pfifo1_rd_data[8], pfifo1_rd_data[9] };
  assign _1382_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[17], pfifo1_rd_data[18], pfifo1_rd_data[19], pfifo1_rd_data[20], pfifo1_rd_data[21], pfifo1_rd_data[22], pfifo1_rd_data[23], pfifo1_rd_data[24], pfifo1_rd_data[25] };
  assign _1383_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[33], pfifo1_rd_data[34], pfifo1_rd_data[35], pfifo1_rd_data[36], pfifo1_rd_data[37], pfifo1_rd_data[38], pfifo1_rd_data[39], pfifo1_rd_data[40], pfifo1_rd_data[41] };
  assign _1384_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[49], pfifo1_rd_data[50], pfifo1_rd_data[51], pfifo1_rd_data[52], pfifo1_rd_data[53], pfifo1_rd_data[54], pfifo1_rd_data[55], pfifo1_rd_data[56], pfifo1_rd_data[57] };
  assign _1385_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[65], pfifo1_rd_data[66], pfifo1_rd_data[67], pfifo1_rd_data[68], pfifo1_rd_data[69], pfifo1_rd_data[70], pfifo1_rd_data[71], pfifo1_rd_data[72], pfifo1_rd_data[73] };
  assign _1386_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[81], pfifo1_rd_data[82], pfifo1_rd_data[83], pfifo1_rd_data[84], pfifo1_rd_data[85], pfifo1_rd_data[86], pfifo1_rd_data[87], pfifo1_rd_data[88], pfifo1_rd_data[89] };
  assign _1387_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[97], pfifo1_rd_data[98], pfifo1_rd_data[99], pfifo1_rd_data[100], pfifo1_rd_data[101], pfifo1_rd_data[102], pfifo1_rd_data[103], pfifo1_rd_data[104], pfifo1_rd_data[105] };
  assign _1388_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo1_rd_data[113], pfifo1_rd_data[114], pfifo1_rd_data[115], pfifo1_rd_data[116], pfifo1_rd_data[117], pfifo1_rd_data[118], pfifo1_rd_data[119], pfifo1_rd_data[120], pfifo1_rd_data[121] };
  assign _1389_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[1], pfifo2_rd_data[2], pfifo2_rd_data[3], pfifo2_rd_data[4], pfifo2_rd_data[5], pfifo2_rd_data[6], pfifo2_rd_data[7], pfifo2_rd_data[8], pfifo2_rd_data[9] };
  assign _1390_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[17], pfifo2_rd_data[18], pfifo2_rd_data[19], pfifo2_rd_data[20], pfifo2_rd_data[21], pfifo2_rd_data[22], pfifo2_rd_data[23], pfifo2_rd_data[24], pfifo2_rd_data[25] };
  assign _1391_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[33], pfifo2_rd_data[34], pfifo2_rd_data[35], pfifo2_rd_data[36], pfifo2_rd_data[37], pfifo2_rd_data[38], pfifo2_rd_data[39], pfifo2_rd_data[40], pfifo2_rd_data[41] };
  assign _1392_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[49], pfifo2_rd_data[50], pfifo2_rd_data[51], pfifo2_rd_data[52], pfifo2_rd_data[53], pfifo2_rd_data[54], pfifo2_rd_data[55], pfifo2_rd_data[56], pfifo2_rd_data[57] };
  assign _1393_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[65], pfifo2_rd_data[66], pfifo2_rd_data[67], pfifo2_rd_data[68], pfifo2_rd_data[69], pfifo2_rd_data[70], pfifo2_rd_data[71], pfifo2_rd_data[72], pfifo2_rd_data[73] };
  assign _1394_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[81], pfifo2_rd_data[82], pfifo2_rd_data[83], pfifo2_rd_data[84], pfifo2_rd_data[85], pfifo2_rd_data[86], pfifo2_rd_data[87], pfifo2_rd_data[88], pfifo2_rd_data[89] };
  assign _1395_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[97], pfifo2_rd_data[98], pfifo2_rd_data[99], pfifo2_rd_data[100], pfifo2_rd_data[101], pfifo2_rd_data[102], pfifo2_rd_data[103], pfifo2_rd_data[104], pfifo2_rd_data[105] };
  assign _1396_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo2_rd_data[113], pfifo2_rd_data[114], pfifo2_rd_data[115], pfifo2_rd_data[116], pfifo2_rd_data[117], pfifo2_rd_data[118], pfifo2_rd_data[119], pfifo2_rd_data[120], pfifo2_rd_data[121] };
  assign _1397_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[1], pfifo3_rd_data[2], pfifo3_rd_data[3], pfifo3_rd_data[4], pfifo3_rd_data[5], pfifo3_rd_data[6], pfifo3_rd_data[7], pfifo3_rd_data[8], pfifo3_rd_data[9] };
  assign _1398_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[17], pfifo3_rd_data[18], pfifo3_rd_data[19], pfifo3_rd_data[20], pfifo3_rd_data[21], pfifo3_rd_data[22], pfifo3_rd_data[23], pfifo3_rd_data[24], pfifo3_rd_data[25] };
  assign _1399_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[33], pfifo3_rd_data[34], pfifo3_rd_data[35], pfifo3_rd_data[36], pfifo3_rd_data[37], pfifo3_rd_data[38], pfifo3_rd_data[39], pfifo3_rd_data[40], pfifo3_rd_data[41] };
  assign _1400_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[49], pfifo3_rd_data[50], pfifo3_rd_data[51], pfifo3_rd_data[52], pfifo3_rd_data[53], pfifo3_rd_data[54], pfifo3_rd_data[55], pfifo3_rd_data[56], pfifo3_rd_data[57] };
  assign _1401_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[65], pfifo3_rd_data[66], pfifo3_rd_data[67], pfifo3_rd_data[68], pfifo3_rd_data[69], pfifo3_rd_data[70], pfifo3_rd_data[71], pfifo3_rd_data[72], pfifo3_rd_data[73] };
  assign _1402_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[81], pfifo3_rd_data[82], pfifo3_rd_data[83], pfifo3_rd_data[84], pfifo3_rd_data[85], pfifo3_rd_data[86], pfifo3_rd_data[87], pfifo3_rd_data[88], pfifo3_rd_data[89] };
  assign _1403_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[97], pfifo3_rd_data[98], pfifo3_rd_data[99], pfifo3_rd_data[100], pfifo3_rd_data[101], pfifo3_rd_data[102], pfifo3_rd_data[103], pfifo3_rd_data[104], pfifo3_rd_data[105] };
  assign _1404_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1482" *) { pfifo3_rd_data[113], pfifo3_rd_data[114], pfifo3_rd_data[115], pfifo3_rd_data[116], pfifo3_rd_data[117], pfifo3_rd_data[118], pfifo3_rd_data[119], pfifo3_rd_data[120], pfifo3_rd_data[121] };
  assign _0814_[22:0] = pfifo0_rd_data[9:0] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0324_;
  assign _0815_[22:0] = pfifo0_rd_data[25:16] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0325_;
  assign _0816_[22:0] = pfifo0_rd_data[41:32] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0326_;
  assign _0817_[22:0] = pfifo0_rd_data[57:48] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0327_;
  assign _1405_[22:0] = pfifo0_rd_data[73:64] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0328_;
  assign _0818_[22:0] = pfifo0_rd_data[89:80] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0329_;
  assign _0819_[22:0] = pfifo0_rd_data[105:96] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0330_;
  assign _0820_[22:0] = pfifo0_rd_data[121:112] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0331_;
  assign _0821_[22:0] = pfifo1_rd_data[9:0] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0332_;
  assign _0822_[22:0] = pfifo1_rd_data[25:16] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0333_;
  assign _0823_[22:0] = pfifo1_rd_data[41:32] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0334_;
  assign _0824_[22:0] = pfifo1_rd_data[57:48] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0335_;
  assign _0825_[22:0] = pfifo1_rd_data[73:64] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0336_;
  assign _0826_[22:0] = pfifo1_rd_data[89:80] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0337_;
  assign _0827_[22:0] = pfifo1_rd_data[105:96] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0338_;
  assign _0828_[22:0] = pfifo1_rd_data[121:112] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0339_;
  assign _0829_[22:0] = pfifo2_rd_data[9:0] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0340_;
  assign _0830_[22:0] = pfifo2_rd_data[25:16] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0341_;
  assign _0831_[22:0] = pfifo2_rd_data[41:32] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0342_;
  assign _0832_[22:0] = pfifo2_rd_data[57:48] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0343_;
  assign _1406_[22:0] = pfifo2_rd_data[73:64] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0344_;
  assign _0833_[22:0] = pfifo2_rd_data[89:80] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0345_;
  assign _0834_[22:0] = pfifo2_rd_data[105:96] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0346_;
  assign _0835_[22:0] = pfifo2_rd_data[121:112] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0347_;
  assign _0836_[22:0] = pfifo3_rd_data[9:0] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0348_;
  assign _0837_[22:0] = pfifo3_rd_data[25:16] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0349_;
  assign _0838_[22:0] = pfifo3_rd_data[41:32] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0350_;
  assign _0839_[22:0] = pfifo3_rd_data[57:48] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0351_;
  assign _0840_[22:0] = pfifo3_rd_data[73:64] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0352_;
  assign _0841_[22:0] = pfifo3_rd_data[89:80] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0353_;
  assign _0842_[22:0] = pfifo3_rd_data[105:96] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0354_;
  assign _0843_[22:0] = pfifo3_rd_data[121:112] << (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1450" *) _0355_;
  assign _0844_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0676_;
  assign _0845_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0677_;
  assign _0846_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0678_;
  assign _0847_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0679_;
  assign _1407_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) { _0780_[3:1], _0680_ };
  assign _0848_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0681_;
  assign _0849_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0682_;
  assign _0850_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0683_;
  assign _0851_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0684_;
  assign _0852_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0685_;
  assign _1408_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0686_;
  assign _1409_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0687_;
  assign _0853_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0688_;
  assign _0854_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0689_;
  assign _0855_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0690_;
  assign _0856_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0691_;
  assign _0857_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0692_;
  assign _0858_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0693_;
  assign _0859_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0694_;
  assign _0860_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0695_;
  assign _1410_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) { _0781_[3:1], _0696_ };
  assign _0861_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0697_;
  assign _0862_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0698_;
  assign _0863_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0699_;
  assign _1411_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0700_;
  assign _1412_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0701_;
  assign _1413_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0702_;
  assign _1414_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0703_;
  assign _0864_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0704_;
  assign _0865_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0705_;
  assign _0866_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0706_;
  assign _0867_[7:0] = 7'b1110001 - (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1448" *) _0707_;
  assign pfifo_data = cfg_di_16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1139" *) pfifo_data_16 : pfifo_data_8;
  assign _1415_ = sfifo_sel ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1158" *) sfifo_data : 512'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign dat_data = pfifo_sel ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1158" *) pfifo_data : _1415_;
  assign sum_of_inf = beat_cnt[0] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:637" *) sum1_of_inf : sum0_of_inf;
  assign sum_of_nan = beat_cnt[0] ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:691" *) sum1_of_nan : sum0_of_nan;
  assign mode_norm_pfifo0_sel = cfg_di_int8 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:720" *) mode_norm_pfifo0_sel_8 : mode_norm_pfifo0_sel_16;
  assign mode_norm_pfifo1_sel = cfg_di_int8 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:721" *) mode_norm_pfifo1_sel_8 : mode_norm_pfifo0_sel_16;
  assign mode_norm_pfifo2_sel = cfg_di_int8 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:722" *) mode_norm_pfifo2_sel_8 : beat_cnt[0];
  assign mode_norm_pfifo3_sel = cfg_di_int8 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:723" *) mode_norm_pfifo3_sel_8 : beat_cnt[0];
  assign pfifo0_sel = _1063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:730" *) mode_norm_pfifo0_sel_8 : mode_norm_pfifo0_sel;
  assign pfifo1_sel = _1063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:731" *) mode_norm_pfifo0_sel_8 : mode_norm_pfifo1_sel;
  assign pfifo2_sel = _1063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:732" *) mode_norm_pfifo2_sel_8 : mode_norm_pfifo2_sel;
  assign pfifo3_sel = _1063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:733" *) mode_norm_pfifo2_sel_8 : mode_norm_pfifo3_sel;
  assign sfifo0_sel = _1063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:734" *) mode_norm_pfifo1_sel_8 : 1'b0;
  assign sfifo1_sel = _1063_ ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:735" *) mode_norm_pfifo3_sel_8 : 1'b0;
  assign pfifo0_data_ext_byte0_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:852" *) pfifo0_data_ext_byte0_fp16[30:0] : { pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15:0] };
  assign pfifo0_data_ext_byte1_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:853" *) pfifo0_data_ext_byte1_fp16[30:0] : { pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31:16] };
  assign pfifo0_data_ext_byte2_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:854" *) pfifo0_data_ext_byte2_fp16[30:0] : { pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47:32] };
  assign pfifo0_data_ext_byte3_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:855" *) pfifo0_data_ext_byte3_fp16[30:0] : { pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63:48] };
  assign pfifo0_data_ext_byte4_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:856" *) pfifo0_data_ext_byte4_fp16[30:0] : { pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79:64] };
  assign pfifo0_data_ext_byte5_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:857" *) pfifo0_data_ext_byte5_fp16[30:0] : { pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95:80] };
  assign pfifo0_data_ext_byte6_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:858" *) pfifo0_data_ext_byte6_fp16[30:0] : { pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111:96] };
  assign pfifo0_data_ext_byte7_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:859" *) pfifo0_data_ext_byte7_fp16[30:0] : { pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127:112] };
  assign pfifo1_data_ext_byte0_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:860" *) pfifo1_data_ext_byte0_fp16[30:0] : { pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15:0] };
  assign pfifo1_data_ext_byte1_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:861" *) pfifo1_data_ext_byte1_fp16[30:0] : { pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31:16] };
  assign pfifo1_data_ext_byte2_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:862" *) pfifo1_data_ext_byte2_fp16[30:0] : { pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47:32] };
  assign pfifo1_data_ext_byte3_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:863" *) pfifo1_data_ext_byte3_fp16[30:0] : { pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63:48] };
  assign pfifo1_data_ext_byte4_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:864" *) pfifo1_data_ext_byte4_fp16[30:0] : { pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79:64] };
  assign pfifo1_data_ext_byte5_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:865" *) pfifo1_data_ext_byte5_fp16[30:0] : { pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95:80] };
  assign pfifo1_data_ext_byte6_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:866" *) pfifo1_data_ext_byte6_fp16[30:0] : { pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111:96] };
  assign pfifo1_data_ext_byte7_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:867" *) pfifo1_data_ext_byte7_fp16[30:0] : { pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127:112] };
  assign pfifo2_data_ext_byte0_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:868" *) pfifo2_data_ext_byte0_fp16[30:0] : { pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15:0] };
  assign pfifo2_data_ext_byte1_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:869" *) pfifo2_data_ext_byte1_fp16[30:0] : { pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31:16] };
  assign pfifo2_data_ext_byte2_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:870" *) pfifo2_data_ext_byte2_fp16[30:0] : { pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47:32] };
  assign pfifo2_data_ext_byte3_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:871" *) pfifo2_data_ext_byte3_fp16[30:0] : { pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63:48] };
  assign pfifo2_data_ext_byte4_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:872" *) pfifo2_data_ext_byte4_fp16[30:0] : { pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79:64] };
  assign pfifo2_data_ext_byte5_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:873" *) pfifo2_data_ext_byte5_fp16[30:0] : { pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95:80] };
  assign pfifo2_data_ext_byte6_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:874" *) pfifo2_data_ext_byte6_fp16[30:0] : { pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111:96] };
  assign pfifo2_data_ext_byte7_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:875" *) pfifo2_data_ext_byte7_fp16[30:0] : { pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127:112] };
  assign pfifo3_data_ext_byte0_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:876" *) pfifo3_data_ext_byte0_fp16[30:0] : { pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15:0] };
  assign pfifo3_data_ext_byte1_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:877" *) pfifo3_data_ext_byte1_fp16[30:0] : { pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31:16] };
  assign pfifo3_data_ext_byte2_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:878" *) pfifo3_data_ext_byte2_fp16[30:0] : { pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47:32] };
  assign pfifo3_data_ext_byte3_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:879" *) pfifo3_data_ext_byte3_fp16[30:0] : { pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63:48] };
  assign pfifo3_data_ext_byte4_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:880" *) pfifo3_data_ext_byte4_fp16[30:0] : { pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79:64] };
  assign pfifo3_data_ext_byte5_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:881" *) pfifo3_data_ext_byte5_fp16[30:0] : { pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95:80] };
  assign pfifo3_data_ext_byte6_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:882" *) pfifo3_data_ext_byte6_fp16[30:0] : { pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111:96] };
  assign pfifo3_data_ext_byte7_16[30:0] = cfg_di_fp16 ? (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:883" *) pfifo3_data_ext_byte7_fp16[30:0] : { pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127:112] };
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_MRDMA_EG_dout.v:1169" *)
  NV_NVDLA_SDP_MRDMA_EG_DOUT_pipe_p1 pipe_p1 (
    .dat_pd({ dat_batch_end, dat_batch_end, dat_data }),
    .dat_rdy(dat_rdy),
    .dat_vld(dat_vld),
    .nvdla_core_clk(nvdla_core_clk),
    .nvdla_core_rstn(nvdla_core_rstn),
    .sdp_mrdma2cmux_pd(sdp_mrdma2cmux_pd),
    .sdp_mrdma2cmux_ready(sdp_mrdma2cmux_ready),
    .sdp_mrdma2cmux_valid(sdp_mrdma2cmux_valid)
  );
  assign _0780_[0] = _0680_;
  assign _0781_[0] = _0696_;
  assign cfg_perf_nan_inf_count_en = reg2dp_perf_nan_inf_count_en;
  assign cmd2dat_dma_cube_end = cmd2dat_dma_pd[14];
  assign cmd2dat_dma_size = cmd2dat_dma_pd[13:0];
  assign dat_layer_end = dat_batch_end;
  assign dat_pd = { dat_batch_end, dat_batch_end, dat_data };
  assign dp2reg_status_inf_input_num = inf_input_cnt;
  assign dp2reg_status_nan_input_num = nan_input_cnt;
  assign mode_16to8_pfifo0_sel = mode_norm_pfifo0_sel_8;
  assign mode_16to8_pfifo1_sel = mode_norm_pfifo0_sel_8;
  assign mode_16to8_pfifo2_sel = mode_norm_pfifo2_sel_8;
  assign mode_16to8_pfifo3_sel = mode_norm_pfifo2_sel_8;
  assign mode_16to8_sfifo0_sel = mode_norm_pfifo1_sel_8;
  assign mode_16to8_sfifo1_sel = mode_norm_pfifo3_sel_8;
  assign mode_norm_pfifo1_sel_16 = mode_norm_pfifo0_sel_16;
  assign mode_norm_pfifo2_sel_16 = beat_cnt[0];
  assign mode_norm_pfifo3_sel_16 = beat_cnt[0];
  assign pfifo0_data_16 = { pfifo0_rd_data[127], pfifo0_data_ext_byte7_16[30:0], pfifo0_rd_data[111], pfifo0_data_ext_byte6_16[30:0], pfifo0_rd_data[95], pfifo0_data_ext_byte5_16[30:0], pfifo0_rd_data[79], pfifo0_data_ext_byte4_16[30:0], pfifo0_rd_data[63], pfifo0_data_ext_byte3_16[30:0], pfifo0_rd_data[47], pfifo0_data_ext_byte2_16[30:0], pfifo0_rd_data[31], pfifo0_data_ext_byte1_16[30:0], pfifo0_rd_data[15], pfifo0_data_ext_byte0_16[30:0] };
  assign pfifo0_data_byte0_16 = pfifo0_rd_data[15:0];
  assign pfifo0_data_byte0_8 = pfifo0_rd_data[7:0];
  assign pfifo0_data_byte10_8 = pfifo0_rd_data[87:80];
  assign pfifo0_data_byte11_8 = pfifo0_rd_data[95:88];
  assign pfifo0_data_byte12_8 = pfifo0_rd_data[103:96];
  assign pfifo0_data_byte13_8 = pfifo0_rd_data[111:104];
  assign pfifo0_data_byte14_8 = pfifo0_rd_data[119:112];
  assign pfifo0_data_byte15_8 = pfifo0_rd_data[127:120];
  assign pfifo0_data_byte1_16 = pfifo0_rd_data[31:16];
  assign pfifo0_data_byte1_8 = pfifo0_rd_data[15:8];
  assign pfifo0_data_byte2_16 = pfifo0_rd_data[47:32];
  assign pfifo0_data_byte2_8 = pfifo0_rd_data[23:16];
  assign pfifo0_data_byte3_16 = pfifo0_rd_data[63:48];
  assign pfifo0_data_byte3_8 = pfifo0_rd_data[31:24];
  assign pfifo0_data_byte4_16 = pfifo0_rd_data[79:64];
  assign pfifo0_data_byte4_8 = pfifo0_rd_data[39:32];
  assign pfifo0_data_byte5_16 = pfifo0_rd_data[95:80];
  assign pfifo0_data_byte5_8 = pfifo0_rd_data[47:40];
  assign pfifo0_data_byte6_16 = pfifo0_rd_data[111:96];
  assign pfifo0_data_byte6_8 = pfifo0_rd_data[55:48];
  assign pfifo0_data_byte7_16 = pfifo0_rd_data[127:112];
  assign pfifo0_data_byte7_8 = pfifo0_rd_data[63:56];
  assign pfifo0_data_byte8_8 = pfifo0_rd_data[71:64];
  assign pfifo0_data_byte9_8 = pfifo0_rd_data[79:72];
  assign pfifo0_data_ext_byte0_16[31] = pfifo0_rd_data[15];
  assign pfifo0_data_ext_byte0_8 = { pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7:0] };
  assign pfifo0_data_ext_byte0_fp16[31] = pfifo0_rd_data[15];
  assign pfifo0_data_ext_byte0_int16 = { pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15:0] };
  assign pfifo0_data_ext_byte10_8 = { pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87:80] };
  assign pfifo0_data_ext_byte11_8 = { pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95:88] };
  assign pfifo0_data_ext_byte12_8 = { pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103:96] };
  assign pfifo0_data_ext_byte13_8 = { pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111:104] };
  assign pfifo0_data_ext_byte14_8 = { pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119:112] };
  assign pfifo0_data_ext_byte15_8 = { pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127:120] };
  assign pfifo0_data_ext_byte1_16[31] = pfifo0_rd_data[31];
  assign pfifo0_data_ext_byte1_8 = { pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15:8] };
  assign pfifo0_data_ext_byte1_fp16[31] = pfifo0_rd_data[31];
  assign pfifo0_data_ext_byte1_int16 = { pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31:16] };
  assign pfifo0_data_ext_byte2_16[31] = pfifo0_rd_data[47];
  assign pfifo0_data_ext_byte2_8 = { pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23:16] };
  assign pfifo0_data_ext_byte2_fp16[31] = pfifo0_rd_data[47];
  assign pfifo0_data_ext_byte2_int16 = { pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47:32] };
  assign pfifo0_data_ext_byte3_16[31] = pfifo0_rd_data[63];
  assign pfifo0_data_ext_byte3_8 = { pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31:24] };
  assign pfifo0_data_ext_byte3_fp16[31] = pfifo0_rd_data[63];
  assign pfifo0_data_ext_byte3_int16 = { pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63:48] };
  assign pfifo0_data_ext_byte4_16[31] = pfifo0_rd_data[79];
  assign pfifo0_data_ext_byte4_8 = { pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39:32] };
  assign pfifo0_data_ext_byte4_fp16[31] = pfifo0_rd_data[79];
  assign pfifo0_data_ext_byte4_int16 = { pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79:64] };
  assign pfifo0_data_ext_byte5_16[31] = pfifo0_rd_data[95];
  assign pfifo0_data_ext_byte5_8 = { pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47:40] };
  assign pfifo0_data_ext_byte5_fp16[31] = pfifo0_rd_data[95];
  assign pfifo0_data_ext_byte5_int16 = { pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95:80] };
  assign pfifo0_data_ext_byte6_16[31] = pfifo0_rd_data[111];
  assign pfifo0_data_ext_byte6_8 = { pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55:48] };
  assign pfifo0_data_ext_byte6_fp16[31] = pfifo0_rd_data[111];
  assign pfifo0_data_ext_byte6_int16 = { pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111:96] };
  assign pfifo0_data_ext_byte7_16[31] = pfifo0_rd_data[127];
  assign pfifo0_data_ext_byte7_8 = { pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63:56] };
  assign pfifo0_data_ext_byte7_fp16[31] = pfifo0_rd_data[127];
  assign pfifo0_data_ext_byte7_int16 = { pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127:112] };
  assign pfifo0_data_ext_byte8_8 = { pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71:64] };
  assign pfifo0_data_ext_byte9_8 = { pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79:72] };
  assign pfifo1_data_16 = { pfifo1_rd_data[127], pfifo1_data_ext_byte7_16[30:0], pfifo1_rd_data[111], pfifo1_data_ext_byte6_16[30:0], pfifo1_rd_data[95], pfifo1_data_ext_byte5_16[30:0], pfifo1_rd_data[79], pfifo1_data_ext_byte4_16[30:0], pfifo1_rd_data[63], pfifo1_data_ext_byte3_16[30:0], pfifo1_rd_data[47], pfifo1_data_ext_byte2_16[30:0], pfifo1_rd_data[31], pfifo1_data_ext_byte1_16[30:0], pfifo1_rd_data[15], pfifo1_data_ext_byte0_16[30:0] };
  assign pfifo1_data_byte0_16 = pfifo1_rd_data[15:0];
  assign pfifo1_data_byte0_8 = pfifo1_rd_data[7:0];
  assign pfifo1_data_byte10_8 = pfifo1_rd_data[87:80];
  assign pfifo1_data_byte11_8 = pfifo1_rd_data[95:88];
  assign pfifo1_data_byte12_8 = pfifo1_rd_data[103:96];
  assign pfifo1_data_byte13_8 = pfifo1_rd_data[111:104];
  assign pfifo1_data_byte14_8 = pfifo1_rd_data[119:112];
  assign pfifo1_data_byte15_8 = pfifo1_rd_data[127:120];
  assign pfifo1_data_byte1_16 = pfifo1_rd_data[31:16];
  assign pfifo1_data_byte1_8 = pfifo1_rd_data[15:8];
  assign pfifo1_data_byte2_16 = pfifo1_rd_data[47:32];
  assign pfifo1_data_byte2_8 = pfifo1_rd_data[23:16];
  assign pfifo1_data_byte3_16 = pfifo1_rd_data[63:48];
  assign pfifo1_data_byte3_8 = pfifo1_rd_data[31:24];
  assign pfifo1_data_byte4_16 = pfifo1_rd_data[79:64];
  assign pfifo1_data_byte4_8 = pfifo1_rd_data[39:32];
  assign pfifo1_data_byte5_16 = pfifo1_rd_data[95:80];
  assign pfifo1_data_byte5_8 = pfifo1_rd_data[47:40];
  assign pfifo1_data_byte6_16 = pfifo1_rd_data[111:96];
  assign pfifo1_data_byte6_8 = pfifo1_rd_data[55:48];
  assign pfifo1_data_byte7_16 = pfifo1_rd_data[127:112];
  assign pfifo1_data_byte7_8 = pfifo1_rd_data[63:56];
  assign pfifo1_data_byte8_8 = pfifo1_rd_data[71:64];
  assign pfifo1_data_byte9_8 = pfifo1_rd_data[79:72];
  assign pfifo1_data_ext_byte0_16[31] = pfifo1_rd_data[15];
  assign pfifo1_data_ext_byte0_8 = { pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7:0] };
  assign pfifo1_data_ext_byte0_fp16[31] = pfifo1_rd_data[15];
  assign pfifo1_data_ext_byte0_int16 = { pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15:0] };
  assign pfifo1_data_ext_byte10_8 = { pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87:80] };
  assign pfifo1_data_ext_byte11_8 = { pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95:88] };
  assign pfifo1_data_ext_byte12_8 = { pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103:96] };
  assign pfifo1_data_ext_byte13_8 = { pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111:104] };
  assign pfifo1_data_ext_byte14_8 = { pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119:112] };
  assign pfifo1_data_ext_byte15_8 = { pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127:120] };
  assign pfifo1_data_ext_byte1_16[31] = pfifo1_rd_data[31];
  assign pfifo1_data_ext_byte1_8 = { pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15:8] };
  assign pfifo1_data_ext_byte1_fp16[31] = pfifo1_rd_data[31];
  assign pfifo1_data_ext_byte1_int16 = { pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31:16] };
  assign pfifo1_data_ext_byte2_16[31] = pfifo1_rd_data[47];
  assign pfifo1_data_ext_byte2_8 = { pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23:16] };
  assign pfifo1_data_ext_byte2_fp16[31] = pfifo1_rd_data[47];
  assign pfifo1_data_ext_byte2_int16 = { pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47:32] };
  assign pfifo1_data_ext_byte3_16[31] = pfifo1_rd_data[63];
  assign pfifo1_data_ext_byte3_8 = { pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31:24] };
  assign pfifo1_data_ext_byte3_fp16[31] = pfifo1_rd_data[63];
  assign pfifo1_data_ext_byte3_int16 = { pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63:48] };
  assign pfifo1_data_ext_byte4_16[31] = pfifo1_rd_data[79];
  assign pfifo1_data_ext_byte4_8 = { pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39:32] };
  assign pfifo1_data_ext_byte4_fp16[31] = pfifo1_rd_data[79];
  assign pfifo1_data_ext_byte4_int16 = { pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79:64] };
  assign pfifo1_data_ext_byte5_16[31] = pfifo1_rd_data[95];
  assign pfifo1_data_ext_byte5_8 = { pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47:40] };
  assign pfifo1_data_ext_byte5_fp16[31] = pfifo1_rd_data[95];
  assign pfifo1_data_ext_byte5_int16 = { pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95:80] };
  assign pfifo1_data_ext_byte6_16[31] = pfifo1_rd_data[111];
  assign pfifo1_data_ext_byte6_8 = { pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55:48] };
  assign pfifo1_data_ext_byte6_fp16[31] = pfifo1_rd_data[111];
  assign pfifo1_data_ext_byte6_int16 = { pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111:96] };
  assign pfifo1_data_ext_byte7_16[31] = pfifo1_rd_data[127];
  assign pfifo1_data_ext_byte7_8 = { pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63:56] };
  assign pfifo1_data_ext_byte7_fp16[31] = pfifo1_rd_data[127];
  assign pfifo1_data_ext_byte7_int16 = { pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127:112] };
  assign pfifo1_data_ext_byte8_8 = { pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71:64] };
  assign pfifo1_data_ext_byte9_8 = { pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79:72] };
  assign pfifo2_data_16 = { pfifo2_rd_data[127], pfifo2_data_ext_byte7_16[30:0], pfifo2_rd_data[111], pfifo2_data_ext_byte6_16[30:0], pfifo2_rd_data[95], pfifo2_data_ext_byte5_16[30:0], pfifo2_rd_data[79], pfifo2_data_ext_byte4_16[30:0], pfifo2_rd_data[63], pfifo2_data_ext_byte3_16[30:0], pfifo2_rd_data[47], pfifo2_data_ext_byte2_16[30:0], pfifo2_rd_data[31], pfifo2_data_ext_byte1_16[30:0], pfifo2_rd_data[15], pfifo2_data_ext_byte0_16[30:0] };
  assign pfifo2_data_byte0_16 = pfifo2_rd_data[15:0];
  assign pfifo2_data_byte0_8 = pfifo2_rd_data[7:0];
  assign pfifo2_data_byte10_8 = pfifo2_rd_data[87:80];
  assign pfifo2_data_byte11_8 = pfifo2_rd_data[95:88];
  assign pfifo2_data_byte12_8 = pfifo2_rd_data[103:96];
  assign pfifo2_data_byte13_8 = pfifo2_rd_data[111:104];
  assign pfifo2_data_byte14_8 = pfifo2_rd_data[119:112];
  assign pfifo2_data_byte15_8 = pfifo2_rd_data[127:120];
  assign pfifo2_data_byte1_16 = pfifo2_rd_data[31:16];
  assign pfifo2_data_byte1_8 = pfifo2_rd_data[15:8];
  assign pfifo2_data_byte2_16 = pfifo2_rd_data[47:32];
  assign pfifo2_data_byte2_8 = pfifo2_rd_data[23:16];
  assign pfifo2_data_byte3_16 = pfifo2_rd_data[63:48];
  assign pfifo2_data_byte3_8 = pfifo2_rd_data[31:24];
  assign pfifo2_data_byte4_16 = pfifo2_rd_data[79:64];
  assign pfifo2_data_byte4_8 = pfifo2_rd_data[39:32];
  assign pfifo2_data_byte5_16 = pfifo2_rd_data[95:80];
  assign pfifo2_data_byte5_8 = pfifo2_rd_data[47:40];
  assign pfifo2_data_byte6_16 = pfifo2_rd_data[111:96];
  assign pfifo2_data_byte6_8 = pfifo2_rd_data[55:48];
  assign pfifo2_data_byte7_16 = pfifo2_rd_data[127:112];
  assign pfifo2_data_byte7_8 = pfifo2_rd_data[63:56];
  assign pfifo2_data_byte8_8 = pfifo2_rd_data[71:64];
  assign pfifo2_data_byte9_8 = pfifo2_rd_data[79:72];
  assign pfifo2_data_ext_byte0_16[31] = pfifo2_rd_data[15];
  assign pfifo2_data_ext_byte0_8 = { pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7:0] };
  assign pfifo2_data_ext_byte0_fp16[31] = pfifo2_rd_data[15];
  assign pfifo2_data_ext_byte0_int16 = { pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15:0] };
  assign pfifo2_data_ext_byte10_8 = { pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87:80] };
  assign pfifo2_data_ext_byte11_8 = { pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95:88] };
  assign pfifo2_data_ext_byte12_8 = { pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103:96] };
  assign pfifo2_data_ext_byte13_8 = { pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111:104] };
  assign pfifo2_data_ext_byte14_8 = { pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119:112] };
  assign pfifo2_data_ext_byte15_8 = { pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127:120] };
  assign pfifo2_data_ext_byte1_16[31] = pfifo2_rd_data[31];
  assign pfifo2_data_ext_byte1_8 = { pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15:8] };
  assign pfifo2_data_ext_byte1_fp16[31] = pfifo2_rd_data[31];
  assign pfifo2_data_ext_byte1_int16 = { pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31:16] };
  assign pfifo2_data_ext_byte2_16[31] = pfifo2_rd_data[47];
  assign pfifo2_data_ext_byte2_8 = { pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23:16] };
  assign pfifo2_data_ext_byte2_fp16[31] = pfifo2_rd_data[47];
  assign pfifo2_data_ext_byte2_int16 = { pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47:32] };
  assign pfifo2_data_ext_byte3_16[31] = pfifo2_rd_data[63];
  assign pfifo2_data_ext_byte3_8 = { pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31:24] };
  assign pfifo2_data_ext_byte3_fp16[31] = pfifo2_rd_data[63];
  assign pfifo2_data_ext_byte3_int16 = { pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63:48] };
  assign pfifo2_data_ext_byte4_16[31] = pfifo2_rd_data[79];
  assign pfifo2_data_ext_byte4_8 = { pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39:32] };
  assign pfifo2_data_ext_byte4_fp16[31] = pfifo2_rd_data[79];
  assign pfifo2_data_ext_byte4_int16 = { pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79:64] };
  assign pfifo2_data_ext_byte5_16[31] = pfifo2_rd_data[95];
  assign pfifo2_data_ext_byte5_8 = { pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47:40] };
  assign pfifo2_data_ext_byte5_fp16[31] = pfifo2_rd_data[95];
  assign pfifo2_data_ext_byte5_int16 = { pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95:80] };
  assign pfifo2_data_ext_byte6_16[31] = pfifo2_rd_data[111];
  assign pfifo2_data_ext_byte6_8 = { pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55:48] };
  assign pfifo2_data_ext_byte6_fp16[31] = pfifo2_rd_data[111];
  assign pfifo2_data_ext_byte6_int16 = { pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111:96] };
  assign pfifo2_data_ext_byte7_16[31] = pfifo2_rd_data[127];
  assign pfifo2_data_ext_byte7_8 = { pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63:56] };
  assign pfifo2_data_ext_byte7_fp16[31] = pfifo2_rd_data[127];
  assign pfifo2_data_ext_byte7_int16 = { pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127:112] };
  assign pfifo2_data_ext_byte8_8 = { pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71:64] };
  assign pfifo2_data_ext_byte9_8 = { pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79:72] };
  assign pfifo3_data_16 = { pfifo3_rd_data[127], pfifo3_data_ext_byte7_16[30:0], pfifo3_rd_data[111], pfifo3_data_ext_byte6_16[30:0], pfifo3_rd_data[95], pfifo3_data_ext_byte5_16[30:0], pfifo3_rd_data[79], pfifo3_data_ext_byte4_16[30:0], pfifo3_rd_data[63], pfifo3_data_ext_byte3_16[30:0], pfifo3_rd_data[47], pfifo3_data_ext_byte2_16[30:0], pfifo3_rd_data[31], pfifo3_data_ext_byte1_16[30:0], pfifo3_rd_data[15], pfifo3_data_ext_byte0_16[30:0] };
  assign pfifo3_data_byte0_16 = pfifo3_rd_data[15:0];
  assign pfifo3_data_byte0_8 = pfifo3_rd_data[7:0];
  assign pfifo3_data_byte10_8 = pfifo3_rd_data[87:80];
  assign pfifo3_data_byte11_8 = pfifo3_rd_data[95:88];
  assign pfifo3_data_byte12_8 = pfifo3_rd_data[103:96];
  assign pfifo3_data_byte13_8 = pfifo3_rd_data[111:104];
  assign pfifo3_data_byte14_8 = pfifo3_rd_data[119:112];
  assign pfifo3_data_byte15_8 = pfifo3_rd_data[127:120];
  assign pfifo3_data_byte1_16 = pfifo3_rd_data[31:16];
  assign pfifo3_data_byte1_8 = pfifo3_rd_data[15:8];
  assign pfifo3_data_byte2_16 = pfifo3_rd_data[47:32];
  assign pfifo3_data_byte2_8 = pfifo3_rd_data[23:16];
  assign pfifo3_data_byte3_16 = pfifo3_rd_data[63:48];
  assign pfifo3_data_byte3_8 = pfifo3_rd_data[31:24];
  assign pfifo3_data_byte4_16 = pfifo3_rd_data[79:64];
  assign pfifo3_data_byte4_8 = pfifo3_rd_data[39:32];
  assign pfifo3_data_byte5_16 = pfifo3_rd_data[95:80];
  assign pfifo3_data_byte5_8 = pfifo3_rd_data[47:40];
  assign pfifo3_data_byte6_16 = pfifo3_rd_data[111:96];
  assign pfifo3_data_byte6_8 = pfifo3_rd_data[55:48];
  assign pfifo3_data_byte7_16 = pfifo3_rd_data[127:112];
  assign pfifo3_data_byte7_8 = pfifo3_rd_data[63:56];
  assign pfifo3_data_byte8_8 = pfifo3_rd_data[71:64];
  assign pfifo3_data_byte9_8 = pfifo3_rd_data[79:72];
  assign pfifo3_data_ext_byte0_16[31] = pfifo3_rd_data[15];
  assign pfifo3_data_ext_byte0_8 = { pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7:0] };
  assign pfifo3_data_ext_byte0_fp16[31] = pfifo3_rd_data[15];
  assign pfifo3_data_ext_byte0_int16 = { pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15:0] };
  assign pfifo3_data_ext_byte10_8 = { pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87:80] };
  assign pfifo3_data_ext_byte11_8 = { pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95:88] };
  assign pfifo3_data_ext_byte12_8 = { pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103:96] };
  assign pfifo3_data_ext_byte13_8 = { pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111:104] };
  assign pfifo3_data_ext_byte14_8 = { pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119:112] };
  assign pfifo3_data_ext_byte15_8 = { pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127:120] };
  assign pfifo3_data_ext_byte1_16[31] = pfifo3_rd_data[31];
  assign pfifo3_data_ext_byte1_8 = { pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15:8] };
  assign pfifo3_data_ext_byte1_fp16[31] = pfifo3_rd_data[31];
  assign pfifo3_data_ext_byte1_int16 = { pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31:16] };
  assign pfifo3_data_ext_byte2_16[31] = pfifo3_rd_data[47];
  assign pfifo3_data_ext_byte2_8 = { pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23:16] };
  assign pfifo3_data_ext_byte2_fp16[31] = pfifo3_rd_data[47];
  assign pfifo3_data_ext_byte2_int16 = { pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47:32] };
  assign pfifo3_data_ext_byte3_16[31] = pfifo3_rd_data[63];
  assign pfifo3_data_ext_byte3_8 = { pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31:24] };
  assign pfifo3_data_ext_byte3_fp16[31] = pfifo3_rd_data[63];
  assign pfifo3_data_ext_byte3_int16 = { pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63:48] };
  assign pfifo3_data_ext_byte4_16[31] = pfifo3_rd_data[79];
  assign pfifo3_data_ext_byte4_8 = { pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39:32] };
  assign pfifo3_data_ext_byte4_fp16[31] = pfifo3_rd_data[79];
  assign pfifo3_data_ext_byte4_int16 = { pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79:64] };
  assign pfifo3_data_ext_byte5_16[31] = pfifo3_rd_data[95];
  assign pfifo3_data_ext_byte5_8 = { pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47:40] };
  assign pfifo3_data_ext_byte5_fp16[31] = pfifo3_rd_data[95];
  assign pfifo3_data_ext_byte5_int16 = { pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95:80] };
  assign pfifo3_data_ext_byte6_16[31] = pfifo3_rd_data[111];
  assign pfifo3_data_ext_byte6_8 = { pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55:48] };
  assign pfifo3_data_ext_byte6_fp16[31] = pfifo3_rd_data[111];
  assign pfifo3_data_ext_byte6_int16 = { pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111:96] };
  assign pfifo3_data_ext_byte7_16[31] = pfifo3_rd_data[127];
  assign pfifo3_data_ext_byte7_8 = { pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63:56] };
  assign pfifo3_data_ext_byte7_fp16[31] = pfifo3_rd_data[127];
  assign pfifo3_data_ext_byte7_int16 = { pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127:112] };
  assign pfifo3_data_ext_byte8_8 = { pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71:64] };
  assign pfifo3_data_ext_byte9_8 = { pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79:72] };
  assign pfifo_data0_16 = { pfifo1_rd_data[127], pfifo1_data_ext_byte7_16[30:0], pfifo1_rd_data[111], pfifo1_data_ext_byte6_16[30:0], pfifo1_rd_data[95], pfifo1_data_ext_byte5_16[30:0], pfifo1_rd_data[79], pfifo1_data_ext_byte4_16[30:0], pfifo1_rd_data[63], pfifo1_data_ext_byte3_16[30:0], pfifo1_rd_data[47], pfifo1_data_ext_byte2_16[30:0], pfifo1_rd_data[31], pfifo1_data_ext_byte1_16[30:0], pfifo1_rd_data[15], pfifo1_data_ext_byte0_16[30:0], pfifo0_rd_data[127], pfifo0_data_ext_byte7_16[30:0], pfifo0_rd_data[111], pfifo0_data_ext_byte6_16[30:0], pfifo0_rd_data[95], pfifo0_data_ext_byte5_16[30:0], pfifo0_rd_data[79], pfifo0_data_ext_byte4_16[30:0], pfifo0_rd_data[63], pfifo0_data_ext_byte3_16[30:0], pfifo0_rd_data[47], pfifo0_data_ext_byte2_16[30:0], pfifo0_rd_data[31], pfifo0_data_ext_byte1_16[30:0], pfifo0_rd_data[15], pfifo0_data_ext_byte0_16[30:0] };
  assign pfifo_data0_8 = { pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127], pfifo0_rd_data[127:119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119], pfifo0_rd_data[119:111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111], pfifo0_rd_data[111:103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103], pfifo0_rd_data[103:95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95], pfifo0_rd_data[95:87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87], pfifo0_rd_data[87:79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79], pfifo0_rd_data[79:71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71], pfifo0_rd_data[71:63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63], pfifo0_rd_data[63:55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55], pfifo0_rd_data[55:47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47], pfifo0_rd_data[47:39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39], pfifo0_rd_data[39:31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31], pfifo0_rd_data[31:23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23], pfifo0_rd_data[23:15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15], pfifo0_rd_data[15:7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7], pfifo0_rd_data[7:0] };
  assign pfifo_data1_16 = { pfifo3_rd_data[127], pfifo3_data_ext_byte7_16[30:0], pfifo3_rd_data[111], pfifo3_data_ext_byte6_16[30:0], pfifo3_rd_data[95], pfifo3_data_ext_byte5_16[30:0], pfifo3_rd_data[79], pfifo3_data_ext_byte4_16[30:0], pfifo3_rd_data[63], pfifo3_data_ext_byte3_16[30:0], pfifo3_rd_data[47], pfifo3_data_ext_byte2_16[30:0], pfifo3_rd_data[31], pfifo3_data_ext_byte1_16[30:0], pfifo3_rd_data[15], pfifo3_data_ext_byte0_16[30:0], pfifo2_rd_data[127], pfifo2_data_ext_byte7_16[30:0], pfifo2_rd_data[111], pfifo2_data_ext_byte6_16[30:0], pfifo2_rd_data[95], pfifo2_data_ext_byte5_16[30:0], pfifo2_rd_data[79], pfifo2_data_ext_byte4_16[30:0], pfifo2_rd_data[63], pfifo2_data_ext_byte3_16[30:0], pfifo2_rd_data[47], pfifo2_data_ext_byte2_16[30:0], pfifo2_rd_data[31], pfifo2_data_ext_byte1_16[30:0], pfifo2_rd_data[15], pfifo2_data_ext_byte0_16[30:0] };
  assign pfifo_data1_8 = { pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127], pfifo1_rd_data[127:119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119], pfifo1_rd_data[119:111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111], pfifo1_rd_data[111:103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103], pfifo1_rd_data[103:95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95], pfifo1_rd_data[95:87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87], pfifo1_rd_data[87:79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79], pfifo1_rd_data[79:71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71], pfifo1_rd_data[71:63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63], pfifo1_rd_data[63:55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55], pfifo1_rd_data[55:47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47], pfifo1_rd_data[47:39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39], pfifo1_rd_data[39:31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31], pfifo1_rd_data[31:23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23], pfifo1_rd_data[23:15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15], pfifo1_rd_data[15:7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7], pfifo1_rd_data[7:0] };
  assign pfifo_data2_8 = { pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127], pfifo2_rd_data[127:119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119], pfifo2_rd_data[119:111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111], pfifo2_rd_data[111:103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103], pfifo2_rd_data[103:95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95], pfifo2_rd_data[95:87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87], pfifo2_rd_data[87:79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79], pfifo2_rd_data[79:71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71], pfifo2_rd_data[71:63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63], pfifo2_rd_data[63:55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55], pfifo2_rd_data[55:47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47], pfifo2_rd_data[47:39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39], pfifo2_rd_data[39:31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31], pfifo2_rd_data[31:23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23], pfifo2_rd_data[23:15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15], pfifo2_rd_data[15:7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7], pfifo2_rd_data[7:0] };
  assign pfifo_data3_8 = { pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127], pfifo3_rd_data[127:119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119], pfifo3_rd_data[119:111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111], pfifo3_rd_data[111:103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103], pfifo3_rd_data[103:95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95], pfifo3_rd_data[95:87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87], pfifo3_rd_data[87:79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79], pfifo3_rd_data[79:71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71], pfifo3_rd_data[71:63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63], pfifo3_rd_data[63:55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55], pfifo3_rd_data[55:47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47], pfifo3_rd_data[47:39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39], pfifo3_rd_data[39:31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31], pfifo3_rd_data[31:23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23], pfifo3_rd_data[23:15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15], pfifo3_rd_data[15:7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7], pfifo3_rd_data[7:0] };
  assign sdp_mrdma2cmux_layer_end = sdp_mrdma2cmux_pd[513];
  assign sfifo0_data_16 = { sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255:239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239:223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223:207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207:191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191:175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175:159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159:143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143:127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127:111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111:95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95:79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79:63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63:47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47:31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31:15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15:0] };
  assign sfifo0_data_byte0_16 = sfifo0_rd_data[15:0];
  assign sfifo0_data_byte10_16 = sfifo0_rd_data[175:160];
  assign sfifo0_data_byte11_16 = sfifo0_rd_data[191:176];
  assign sfifo0_data_byte12_16 = sfifo0_rd_data[207:192];
  assign sfifo0_data_byte13_16 = sfifo0_rd_data[223:208];
  assign sfifo0_data_byte14_16 = sfifo0_rd_data[239:224];
  assign sfifo0_data_byte15_16 = sfifo0_rd_data[255:240];
  assign sfifo0_data_byte1_16 = sfifo0_rd_data[31:16];
  assign sfifo0_data_byte2_16 = sfifo0_rd_data[47:32];
  assign sfifo0_data_byte3_16 = sfifo0_rd_data[63:48];
  assign sfifo0_data_byte4_16 = sfifo0_rd_data[79:64];
  assign sfifo0_data_byte5_16 = sfifo0_rd_data[95:80];
  assign sfifo0_data_byte6_16 = sfifo0_rd_data[111:96];
  assign sfifo0_data_byte7_16 = sfifo0_rd_data[127:112];
  assign sfifo0_data_byte8_16 = sfifo0_rd_data[143:128];
  assign sfifo0_data_byte9_16 = sfifo0_rd_data[159:144];
  assign sfifo0_data_ext_byte0_16 = { sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15:0] };
  assign sfifo0_data_ext_byte10_16 = { sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175:160] };
  assign sfifo0_data_ext_byte11_16 = { sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191], sfifo0_rd_data[191:176] };
  assign sfifo0_data_ext_byte12_16 = { sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207], sfifo0_rd_data[207:192] };
  assign sfifo0_data_ext_byte13_16 = { sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223], sfifo0_rd_data[223:208] };
  assign sfifo0_data_ext_byte14_16 = { sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239], sfifo0_rd_data[239:224] };
  assign sfifo0_data_ext_byte15_16 = { sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255], sfifo0_rd_data[255:240] };
  assign sfifo0_data_ext_byte1_16 = { sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31:16] };
  assign sfifo0_data_ext_byte2_16 = { sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47:32] };
  assign sfifo0_data_ext_byte3_16 = { sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63:48] };
  assign sfifo0_data_ext_byte4_16 = { sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79:64] };
  assign sfifo0_data_ext_byte5_16 = { sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95:80] };
  assign sfifo0_data_ext_byte6_16 = { sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111:96] };
  assign sfifo0_data_ext_byte7_16 = { sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127:112] };
  assign sfifo0_data_ext_byte8_16 = { sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143:128] };
  assign sfifo0_data_ext_byte9_16 = { sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159:144] };
  assign { sfifo1_data_16[350:335], sfifo1_data_16[318:303], sfifo1_data_16[286:271], sfifo1_data_16[254:239], sfifo1_data_16[222:207], sfifo1_data_16[190:175], sfifo1_data_16[158:143], sfifo1_data_16[126:111], sfifo1_data_16[94:79], sfifo1_data_16[62:47], sfifo1_data_16[30:15] } = { sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31] };
  assign sfifo1_data_byte0_16 = { sfifo1_data_16[31], sfifo1_data_16[14:0] };
  assign sfifo1_data_byte10_16 = { sfifo1_data_16[351], sfifo1_data_16[334:320] };
  assign sfifo1_data_byte1_16 = { sfifo1_data_16[63], sfifo1_data_16[46:32] };
  assign sfifo1_data_byte2_16 = { sfifo1_data_16[95], sfifo1_data_16[78:64] };
  assign sfifo1_data_byte3_16 = { sfifo1_data_16[127], sfifo1_data_16[110:96] };
  assign sfifo1_data_byte4_16 = { sfifo1_data_16[159], sfifo1_data_16[142:128] };
  assign sfifo1_data_byte5_16 = { sfifo1_data_16[191], sfifo1_data_16[174:160] };
  assign sfifo1_data_byte6_16 = { sfifo1_data_16[223], sfifo1_data_16[206:192] };
  assign sfifo1_data_byte7_16 = { sfifo1_data_16[255], sfifo1_data_16[238:224] };
  assign sfifo1_data_byte8_16 = { sfifo1_data_16[287], sfifo1_data_16[270:256] };
  assign sfifo1_data_byte9_16 = { sfifo1_data_16[319], sfifo1_data_16[302:288] };
  assign sfifo1_data_ext_byte0_16 = { sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[14:0] };
  assign sfifo1_data_ext_byte10_16 = { sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[334:320] };
  assign sfifo1_data_ext_byte11_16 = { sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16 };
  assign sfifo1_data_ext_byte12_16 = { sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16 };
  assign sfifo1_data_ext_byte13_16 = { sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16 };
  assign sfifo1_data_ext_byte14_16 = { sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16 };
  assign sfifo1_data_ext_byte15_16 = { sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16 };
  assign sfifo1_data_ext_byte1_16 = { sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[46:32] };
  assign sfifo1_data_ext_byte2_16 = { sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[78:64] };
  assign sfifo1_data_ext_byte3_16 = { sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[110:96] };
  assign sfifo1_data_ext_byte4_16 = { sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[142:128] };
  assign sfifo1_data_ext_byte5_16 = { sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[174:160] };
  assign sfifo1_data_ext_byte6_16 = { sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[206:192] };
  assign sfifo1_data_ext_byte7_16 = { sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[238:224] };
  assign sfifo1_data_ext_byte8_16 = { sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[270:256] };
  assign sfifo1_data_ext_byte9_16 = { sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[302:288] };
  assign sfifo1_rd_data = { sfifo1_data_16[351], sfifo1_data_16[334:319], sfifo1_data_16[302:287], sfifo1_data_16[270:255], sfifo1_data_16[238:223], sfifo1_data_16[206:191], sfifo1_data_16[174:159], sfifo1_data_16[142:127], sfifo1_data_16[110:95], sfifo1_data_16[78:63], sfifo1_data_16[46:31], sfifo1_data_16[14:0] };
  assign sfifo_data0_16 = { sfifo0_rd_data[176:175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175], sfifo0_rd_data[175:159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159], sfifo0_rd_data[159:143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143], sfifo0_rd_data[143:127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127], sfifo0_rd_data[127:111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111], sfifo0_rd_data[111:95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95], sfifo0_rd_data[95:79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79], sfifo0_rd_data[79:63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63], sfifo0_rd_data[63:47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47], sfifo0_rd_data[47:31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31], sfifo0_rd_data[31:15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15], sfifo0_rd_data[15:0] };
  assign sfifo_data1_16 = { sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16[15], sfifo1_data_byte15_16, sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16[15], sfifo1_data_byte14_16, sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16[15], sfifo1_data_byte13_16, sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16[15], sfifo1_data_byte12_16, sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16[15], sfifo1_data_byte11_16, sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[351], sfifo1_data_16[334:319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[319], sfifo1_data_16[302:287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[287], sfifo1_data_16[270:255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[255], sfifo1_data_16[238:223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[223], sfifo1_data_16[206:191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[191], sfifo1_data_16[174:159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[159], sfifo1_data_16[142:127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[127], sfifo1_data_16[110:95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[95], sfifo1_data_16[78:63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[63], sfifo1_data_16[46:31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[31], sfifo1_data_16[14:0] };
  assign sum_of_sel = beat_cnt[0];
endmodule
