module NV_NVDLA_CDMA_shared_buffer(nvdla_core_clk, nvdla_core_rstn, pwrbus_ram_pd, dc2sbuf_p0_wr_en, dc2sbuf_p0_wr_addr, dc2sbuf_p0_wr_data, dc2sbuf_p1_wr_en, dc2sbuf_p1_wr_addr, dc2sbuf_p1_wr_data, wg2sbuf_p0_wr_en, wg2sbuf_p0_wr_addr, wg2sbuf_p0_wr_data, wg2sbuf_p1_wr_en, wg2sbuf_p1_wr_addr, wg2sbuf_p1_wr_data, img2sbuf_p0_wr_en, img2sbuf_p0_wr_addr, img2sbuf_p0_wr_data, img2sbuf_p1_wr_en, img2sbuf_p1_wr_addr, img2sbuf_p1_wr_data, dc2sbuf_p0_rd_en, dc2sbuf_p0_rd_addr, dc2sbuf_p0_rd_data, dc2sbuf_p1_rd_en, dc2sbuf_p1_rd_addr, dc2sbuf_p1_rd_data, wg2sbuf_p0_rd_en, wg2sbuf_p0_rd_addr, wg2sbuf_p0_rd_data, wg2sbuf_p1_rd_en, wg2sbuf_p1_rd_addr, wg2sbuf_p1_rd_data, img2sbuf_p0_rd_en, img2sbuf_p0_rd_addr, img2sbuf_p0_rd_data, img2sbuf_p1_rd_en, img2sbuf_p1_rd_addr, img2sbuf_p1_rd_data);
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3798" *)
  wire _0000_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4082" *)
  wire [255:0] _0001_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3462" *)
  wire _0002_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3686" *)
  wire _0003_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3476" *)
  wire _0004_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3700" *)
  wire _0005_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3490" *)
  wire _0006_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3714" *)
  wire _0007_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3504" *)
  wire _0008_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3728" *)
  wire _0009_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3518" *)
  wire _0010_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3532" *)
  wire _0011_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3546" *)
  wire _0012_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3560" *)
  wire _0013_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3574" *)
  wire _0014_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3588" *)
  wire _0015_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3602" *)
  wire _0016_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3616" *)
  wire _0017_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3630" *)
  wire _0018_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3644" *)
  wire _0019_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3658" *)
  wire _0020_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3672" *)
  wire _0021_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3805" *)
  wire _0022_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4092" *)
  wire [255:0] _0023_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3469" *)
  wire _0024_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3693" *)
  wire _0025_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3483" *)
  wire _0026_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3707" *)
  wire _0027_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3497" *)
  wire _0028_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3721" *)
  wire _0029_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3511" *)
  wire _0030_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3735" *)
  wire _0031_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3525" *)
  wire _0032_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3539" *)
  wire _0033_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3553" *)
  wire _0034_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3567" *)
  wire _0035_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3581" *)
  wire _0036_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3595" *)
  wire _0037_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3609" *)
  wire _0038_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3623" *)
  wire _0039_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3637" *)
  wire _0040_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3651" *)
  wire _0041_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3665" *)
  wire _0042_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3679" *)
  wire _0043_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1343" *)
  wire [3:0] _0044_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1344" *)
  wire [3:0] _0045_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1345" *)
  wire [3:0] _0046_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1346" *)
  wire [3:0] _0047_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1347" *)
  wire [3:0] _0048_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1348" *)
  wire [3:0] _0049_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1364" *)
  wire [3:0] _0050_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1365" *)
  wire [3:0] _0051_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1366" *)
  wire [3:0] _0052_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1367" *)
  wire [3:0] _0053_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1368" *)
  wire [3:0] _0054_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1369" *)
  wire [3:0] _0055_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1385" *)
  wire [3:0] _0056_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1386" *)
  wire [3:0] _0057_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1387" *)
  wire [3:0] _0058_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1388" *)
  wire [3:0] _0059_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1389" *)
  wire [3:0] _0060_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1390" *)
  wire [3:0] _0061_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1406" *)
  wire [3:0] _0062_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1407" *)
  wire [3:0] _0063_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1408" *)
  wire [3:0] _0064_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1409" *)
  wire [3:0] _0065_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1410" *)
  wire [3:0] _0066_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1411" *)
  wire [3:0] _0067_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1427" *)
  wire [3:0] _0068_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1428" *)
  wire [3:0] _0069_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1429" *)
  wire [3:0] _0070_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1430" *)
  wire [3:0] _0071_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1431" *)
  wire [3:0] _0072_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1432" *)
  wire [3:0] _0073_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1448" *)
  wire [3:0] _0074_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1449" *)
  wire [3:0] _0075_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1450" *)
  wire [3:0] _0076_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1451" *)
  wire [3:0] _0077_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1452" *)
  wire [3:0] _0078_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1453" *)
  wire [3:0] _0079_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1469" *)
  wire [3:0] _0080_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1470" *)
  wire [3:0] _0081_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1471" *)
  wire [3:0] _0082_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1472" *)
  wire [3:0] _0083_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1473" *)
  wire [3:0] _0084_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1474" *)
  wire [3:0] _0085_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1490" *)
  wire [3:0] _0086_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1491" *)
  wire [3:0] _0087_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1492" *)
  wire [3:0] _0088_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1493" *)
  wire [3:0] _0089_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1494" *)
  wire [3:0] _0090_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1495" *)
  wire [3:0] _0091_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1511" *)
  wire [3:0] _0092_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1512" *)
  wire [3:0] _0093_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1513" *)
  wire [3:0] _0094_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1514" *)
  wire [3:0] _0095_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1515" *)
  wire [3:0] _0096_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1516" *)
  wire [3:0] _0097_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1532" *)
  wire [3:0] _0098_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1533" *)
  wire [3:0] _0099_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1534" *)
  wire [3:0] _0100_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1535" *)
  wire [3:0] _0101_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1536" *)
  wire [3:0] _0102_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1537" *)
  wire [3:0] _0103_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1553" *)
  wire [3:0] _0104_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1554" *)
  wire [3:0] _0105_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1555" *)
  wire [3:0] _0106_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1556" *)
  wire [3:0] _0107_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1557" *)
  wire [3:0] _0108_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1558" *)
  wire [3:0] _0109_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1574" *)
  wire [3:0] _0110_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1575" *)
  wire [3:0] _0111_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1576" *)
  wire [3:0] _0112_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1577" *)
  wire [3:0] _0113_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1578" *)
  wire [3:0] _0114_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1579" *)
  wire [3:0] _0115_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1595" *)
  wire [3:0] _0116_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1596" *)
  wire [3:0] _0117_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1597" *)
  wire [3:0] _0118_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1598" *)
  wire [3:0] _0119_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1599" *)
  wire [3:0] _0120_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1600" *)
  wire [3:0] _0121_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1616" *)
  wire [3:0] _0122_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1617" *)
  wire [3:0] _0123_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1618" *)
  wire [3:0] _0124_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1619" *)
  wire [3:0] _0125_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1620" *)
  wire [3:0] _0126_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1621" *)
  wire [3:0] _0127_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1637" *)
  wire [3:0] _0128_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1638" *)
  wire [3:0] _0129_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1639" *)
  wire [3:0] _0130_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1640" *)
  wire [3:0] _0131_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1641" *)
  wire [3:0] _0132_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1642" *)
  wire [3:0] _0133_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1658" *)
  wire [3:0] _0134_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1659" *)
  wire [3:0] _0135_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1660" *)
  wire [3:0] _0136_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1661" *)
  wire [3:0] _0137_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1662" *)
  wire [3:0] _0138_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1663" *)
  wire [3:0] _0139_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1679" *)
  wire [255:0] _0140_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1680" *)
  wire [255:0] _0141_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1681" *)
  wire [255:0] _0142_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1682" *)
  wire [255:0] _0143_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1683" *)
  wire [255:0] _0144_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1684" *)
  wire [255:0] _0145_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1700" *)
  wire [255:0] _0146_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1701" *)
  wire [255:0] _0147_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1702" *)
  wire [255:0] _0148_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1703" *)
  wire [255:0] _0149_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1704" *)
  wire [255:0] _0150_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1705" *)
  wire [255:0] _0151_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1721" *)
  wire [255:0] _0152_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1722" *)
  wire [255:0] _0153_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1723" *)
  wire [255:0] _0154_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1724" *)
  wire [255:0] _0155_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1725" *)
  wire [255:0] _0156_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1726" *)
  wire [255:0] _0157_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1742" *)
  wire [255:0] _0158_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1743" *)
  wire [255:0] _0159_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1744" *)
  wire [255:0] _0160_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1745" *)
  wire [255:0] _0161_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1746" *)
  wire [255:0] _0162_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1747" *)
  wire [255:0] _0163_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1763" *)
  wire [255:0] _0164_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1764" *)
  wire [255:0] _0165_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1765" *)
  wire [255:0] _0166_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1766" *)
  wire [255:0] _0167_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1767" *)
  wire [255:0] _0168_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1768" *)
  wire [255:0] _0169_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1784" *)
  wire [255:0] _0170_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1785" *)
  wire [255:0] _0171_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1786" *)
  wire [255:0] _0172_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1787" *)
  wire [255:0] _0173_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1788" *)
  wire [255:0] _0174_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1789" *)
  wire [255:0] _0175_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1805" *)
  wire [255:0] _0176_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1806" *)
  wire [255:0] _0177_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1807" *)
  wire [255:0] _0178_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1808" *)
  wire [255:0] _0179_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1809" *)
  wire [255:0] _0180_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1810" *)
  wire [255:0] _0181_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1826" *)
  wire [255:0] _0182_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1827" *)
  wire [255:0] _0183_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1828" *)
  wire [255:0] _0184_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1829" *)
  wire [255:0] _0185_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1830" *)
  wire [255:0] _0186_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1831" *)
  wire [255:0] _0187_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1847" *)
  wire [255:0] _0188_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1848" *)
  wire [255:0] _0189_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1849" *)
  wire [255:0] _0190_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1850" *)
  wire [255:0] _0191_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1851" *)
  wire [255:0] _0192_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1852" *)
  wire [255:0] _0193_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1868" *)
  wire [255:0] _0194_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1869" *)
  wire [255:0] _0195_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1870" *)
  wire [255:0] _0196_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1871" *)
  wire [255:0] _0197_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1872" *)
  wire [255:0] _0198_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1873" *)
  wire [255:0] _0199_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1889" *)
  wire [255:0] _0200_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1890" *)
  wire [255:0] _0201_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1891" *)
  wire [255:0] _0202_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1892" *)
  wire [255:0] _0203_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1893" *)
  wire [255:0] _0204_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1894" *)
  wire [255:0] _0205_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1910" *)
  wire [255:0] _0206_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1911" *)
  wire [255:0] _0207_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1912" *)
  wire [255:0] _0208_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1913" *)
  wire [255:0] _0209_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1914" *)
  wire [255:0] _0210_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1915" *)
  wire [255:0] _0211_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1931" *)
  wire [255:0] _0212_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1932" *)
  wire [255:0] _0213_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1933" *)
  wire [255:0] _0214_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1934" *)
  wire [255:0] _0215_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1935" *)
  wire [255:0] _0216_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1936" *)
  wire [255:0] _0217_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1952" *)
  wire [255:0] _0218_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1953" *)
  wire [255:0] _0219_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1954" *)
  wire [255:0] _0220_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1955" *)
  wire [255:0] _0221_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1956" *)
  wire [255:0] _0222_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1957" *)
  wire [255:0] _0223_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1973" *)
  wire [255:0] _0224_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1974" *)
  wire [255:0] _0225_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1975" *)
  wire [255:0] _0226_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1976" *)
  wire [255:0] _0227_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1977" *)
  wire [255:0] _0228_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1978" *)
  wire [255:0] _0229_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1994" *)
  wire [255:0] _0230_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1995" *)
  wire [255:0] _0231_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1996" *)
  wire [255:0] _0232_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1997" *)
  wire [255:0] _0233_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1998" *)
  wire [255:0] _0234_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1999" *)
  wire [255:0] _0235_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3089" *)
  wire [3:0] _0236_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3090" *)
  wire [3:0] _0237_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3091" *)
  wire [3:0] _0238_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3092" *)
  wire [3:0] _0239_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3093" *)
  wire [3:0] _0240_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3094" *)
  wire [3:0] _0241_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3110" *)
  wire [3:0] _0242_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3111" *)
  wire [3:0] _0243_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3114" *)
  wire [3:0] _0244_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3115" *)
  wire [3:0] _0245_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3131" *)
  wire [3:0] _0246_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3132" *)
  wire [3:0] _0247_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3135" *)
  wire [3:0] _0248_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3136" *)
  wire [3:0] _0249_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3152" *)
  wire [3:0] _0250_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3153" *)
  wire [3:0] _0251_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3156" *)
  wire [3:0] _0252_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3157" *)
  wire [3:0] _0253_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3173" *)
  wire [3:0] _0254_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3174" *)
  wire [3:0] _0255_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3175" *)
  wire [3:0] _0256_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3176" *)
  wire [3:0] _0257_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3177" *)
  wire [3:0] _0258_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3178" *)
  wire [3:0] _0259_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3194" *)
  wire [3:0] _0260_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3195" *)
  wire [3:0] _0261_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3198" *)
  wire [3:0] _0262_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3199" *)
  wire [3:0] _0263_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3215" *)
  wire [3:0] _0264_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3216" *)
  wire [3:0] _0265_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3219" *)
  wire [3:0] _0266_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3220" *)
  wire [3:0] _0267_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3236" *)
  wire [3:0] _0268_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3237" *)
  wire [3:0] _0269_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3240" *)
  wire [3:0] _0270_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3241" *)
  wire [3:0] _0271_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3257" *)
  wire [3:0] _0272_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3258" *)
  wire [3:0] _0273_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3259" *)
  wire [3:0] _0274_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3260" *)
  wire [3:0] _0275_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3261" *)
  wire [3:0] _0276_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3262" *)
  wire [3:0] _0277_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3278" *)
  wire [3:0] _0278_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3279" *)
  wire [3:0] _0279_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3282" *)
  wire [3:0] _0280_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3283" *)
  wire [3:0] _0281_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3299" *)
  wire [3:0] _0282_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3300" *)
  wire [3:0] _0283_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3303" *)
  wire [3:0] _0284_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3304" *)
  wire [3:0] _0285_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3320" *)
  wire [3:0] _0286_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3321" *)
  wire [3:0] _0287_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3324" *)
  wire [3:0] _0288_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3325" *)
  wire [3:0] _0289_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3341" *)
  wire [3:0] _0290_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3342" *)
  wire [3:0] _0291_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3343" *)
  wire [3:0] _0292_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3344" *)
  wire [3:0] _0293_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3345" *)
  wire [3:0] _0294_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3346" *)
  wire [3:0] _0295_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3362" *)
  wire [3:0] _0296_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3363" *)
  wire [3:0] _0297_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3366" *)
  wire [3:0] _0298_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3367" *)
  wire [3:0] _0299_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3383" *)
  wire [3:0] _0300_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3384" *)
  wire [3:0] _0301_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3387" *)
  wire [3:0] _0302_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3388" *)
  wire [3:0] _0303_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3404" *)
  wire [3:0] _0304_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3405" *)
  wire [3:0] _0305_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3408" *)
  wire [3:0] _0306_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3409" *)
  wire [3:0] _0307_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3849" *)
  wire [255:0] _0308_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3850" *)
  wire [255:0] _0309_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3851" *)
  wire [255:0] _0310_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3852" *)
  wire [255:0] _0311_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3853" *)
  wire [255:0] _0312_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3854" *)
  wire [255:0] _0313_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3855" *)
  wire [255:0] _0314_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3856" *)
  wire [255:0] _0315_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3857" *)
  wire [255:0] _0316_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3858" *)
  wire [255:0] _0317_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3859" *)
  wire [255:0] _0318_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3860" *)
  wire [255:0] _0319_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3861" *)
  wire [255:0] _0320_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3862" *)
  wire [255:0] _0321_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3863" *)
  wire [255:0] _0322_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3864" *)
  wire [255:0] _0323_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3900" *)
  wire [255:0] _0324_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3901" *)
  wire [255:0] _0325_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3902" *)
  wire [255:0] _0326_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3903" *)
  wire [255:0] _0327_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3904" *)
  wire [255:0] _0328_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3905" *)
  wire [255:0] _0329_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3906" *)
  wire [255:0] _0330_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3907" *)
  wire [255:0] _0331_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3908" *)
  wire [255:0] _0332_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3909" *)
  wire [255:0] _0333_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3910" *)
  wire [255:0] _0334_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3911" *)
  wire [255:0] _0335_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3912" *)
  wire [255:0] _0336_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3913" *)
  wire [255:0] _0337_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3914" *)
  wire [255:0] _0338_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3915" *)
  wire [255:0] _0339_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3927" *)
  wire [255:0] _0340_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3928" *)
  wire [255:0] _0341_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3929" *)
  wire [255:0] _0342_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3930" *)
  wire [255:0] _0343_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3942" *)
  wire [255:0] _0344_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3943" *)
  wire [255:0] _0345_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3944" *)
  wire [255:0] _0346_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3945" *)
  wire [255:0] _0347_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3957" *)
  wire [255:0] _0348_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3958" *)
  wire [255:0] _0349_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3959" *)
  wire [255:0] _0350_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3960" *)
  wire [255:0] _0351_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3972" *)
  wire [255:0] _0352_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3973" *)
  wire [255:0] _0353_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3974" *)
  wire [255:0] _0354_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3975" *)
  wire [255:0] _0355_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3987" *)
  wire [255:0] _0356_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3988" *)
  wire [255:0] _0357_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3989" *)
  wire [255:0] _0358_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3990" *)
  wire [255:0] _0359_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4002" *)
  wire [255:0] _0360_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4003" *)
  wire [255:0] _0361_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4004" *)
  wire [255:0] _0362_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4005" *)
  wire [255:0] _0363_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4017" *)
  wire [255:0] _0364_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4018" *)
  wire [255:0] _0365_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4019" *)
  wire [255:0] _0366_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4020" *)
  wire [255:0] _0367_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4032" *)
  wire [255:0] _0368_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4033" *)
  wire [255:0] _0369_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4034" *)
  wire [255:0] _0370_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4035" *)
  wire [255:0] _0371_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4047" *)
  wire [255:0] _0372_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4048" *)
  wire [255:0] _0373_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4049" *)
  wire [255:0] _0374_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4050" *)
  wire [255:0] _0375_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4062" *)
  wire [255:0] _0376_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4063" *)
  wire [255:0] _0377_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4064" *)
  wire [255:0] _0378_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4065" *)
  wire [255:0] _0379_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1003" *)
  wire _0380_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1009" *)
  wire _0381_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1015" *)
  wire _0382_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1021" *)
  wire _0383_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1027" *)
  wire _0384_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1033" *)
  wire _0385_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1039" *)
  wire _0386_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1045" *)
  wire _0387_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1051" *)
  wire _0388_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1057" *)
  wire _0389_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1063" *)
  wire _0390_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1069" *)
  wire _0391_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1075" *)
  wire _0392_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1081" *)
  wire _0393_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1087" *)
  wire _0394_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2177" *)
  wire _0395_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2183" *)
  wire _0396_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2189" *)
  wire _0397_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2195" *)
  wire _0398_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2201" *)
  wire _0399_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2207" *)
  wire _0400_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2213" *)
  wire _0401_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2219" *)
  wire _0402_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2225" *)
  wire _0403_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2231" *)
  wire _0404_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2237" *)
  wire _0405_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2243" *)
  wire _0406_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2249" *)
  wire _0407_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2255" *)
  wire _0408_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2261" *)
  wire _0409_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2267" *)
  wire _0410_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2273" *)
  wire _0411_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2279" *)
  wire _0412_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2285" *)
  wire _0413_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2291" *)
  wire _0414_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2297" *)
  wire _0415_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2303" *)
  wire _0416_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2309" *)
  wire _0417_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2315" *)
  wire _0418_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2321" *)
  wire _0419_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2327" *)
  wire _0420_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2333" *)
  wire _0421_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2339" *)
  wire _0422_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2345" *)
  wire _0423_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2351" *)
  wire _0424_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2357" *)
  wire _0425_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2363" *)
  wire _0426_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2369" *)
  wire _0427_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2375" *)
  wire _0428_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2381" *)
  wire _0429_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2387" *)
  wire _0430_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2393" *)
  wire _0431_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2399" *)
  wire _0432_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2405" *)
  wire _0433_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2411" *)
  wire _0434_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2417" *)
  wire _0435_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2423" *)
  wire _0436_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2429" *)
  wire _0437_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2435" *)
  wire _0438_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2441" *)
  wire _0439_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2447" *)
  wire _0440_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2453" *)
  wire _0441_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2459" *)
  wire _0442_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2465" *)
  wire _0443_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2471" *)
  wire _0444_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2477" *)
  wire _0445_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2483" *)
  wire _0446_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2489" *)
  wire _0447_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2495" *)
  wire _0448_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2501" *)
  wire _0449_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2507" *)
  wire _0450_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2513" *)
  wire _0451_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2519" *)
  wire _0452_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2525" *)
  wire _0453_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2531" *)
  wire _0454_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2537" *)
  wire _0455_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2543" *)
  wire _0456_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2549" *)
  wire _0457_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2555" *)
  wire _0458_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2561" *)
  wire _0459_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2567" *)
  wire _0460_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2609" *)
  wire _0461_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2615" *)
  wire _0462_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2657" *)
  wire _0463_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2663" *)
  wire _0464_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2705" *)
  wire _0465_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2711" *)
  wire _0466_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3415" *)
  wire _0467_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3421" *)
  wire _0468_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3427" *)
  wire _0469_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3433" *)
  wire _0470_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3439" *)
  wire _0471_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3445" *)
  wire _0472_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3451" *)
  wire _0473_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3457" *)
  wire _0474_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:517" *)
  wire _0475_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:523" *)
  wire _0476_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:529" *)
  wire _0477_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:535" *)
  wire _0478_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:541" *)
  wire _0479_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:547" *)
  wire _0480_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:553" *)
  wire _0481_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:559" *)
  wire _0482_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:565" *)
  wire _0483_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:571" *)
  wire _0484_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:577" *)
  wire _0485_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:583" *)
  wire _0486_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:589" *)
  wire _0487_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:595" *)
  wire _0488_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:601" *)
  wire _0489_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:607" *)
  wire _0490_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:613" *)
  wire _0491_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:619" *)
  wire _0492_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:625" *)
  wire _0493_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:631" *)
  wire _0494_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:637" *)
  wire _0495_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:643" *)
  wire _0496_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:649" *)
  wire _0497_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:655" *)
  wire _0498_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:661" *)
  wire _0499_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:667" *)
  wire _0500_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:673" *)
  wire _0501_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:679" *)
  wire _0502_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:685" *)
  wire _0503_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:691" *)
  wire _0504_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:697" *)
  wire _0505_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:703" *)
  wire _0506_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:709" *)
  wire _0507_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:715" *)
  wire _0508_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:721" *)
  wire _0509_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:727" *)
  wire _0510_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:733" *)
  wire _0511_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:739" *)
  wire _0512_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:745" *)
  wire _0513_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:751" *)
  wire _0514_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:757" *)
  wire _0515_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:763" *)
  wire _0516_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:769" *)
  wire _0517_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:775" *)
  wire _0518_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:781" *)
  wire _0519_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:787" *)
  wire _0520_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:793" *)
  wire _0521_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:799" *)
  wire _0522_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:805" *)
  wire _0523_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:811" *)
  wire _0524_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:817" *)
  wire _0525_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:823" *)
  wire _0526_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:829" *)
  wire _0527_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:835" *)
  wire _0528_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:841" *)
  wire _0529_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:847" *)
  wire _0530_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:853" *)
  wire _0531_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:859" *)
  wire _0532_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:865" *)
  wire _0533_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:871" *)
  wire _0534_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:877" *)
  wire _0535_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:883" *)
  wire _0536_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:889" *)
  wire _0537_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:895" *)
  wire _0538_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:901" *)
  wire _0539_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:907" *)
  wire _0540_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:913" *)
  wire _0541_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:919" *)
  wire _0542_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:925" *)
  wire _0543_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:931" *)
  wire _0544_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:937" *)
  wire _0545_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:943" *)
  wire _0546_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:949" *)
  wire _0547_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:955" *)
  wire _0548_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:961" *)
  wire _0549_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:967" *)
  wire _0550_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:973" *)
  wire _0551_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:979" *)
  wire _0552_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:985" *)
  wire _0553_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:991" *)
  wire _0554_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:997" *)
  wire _0555_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3466" *)
  wire _0556_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3473" *)
  wire _0557_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1098" *)
  wire _0558_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1099" *)
  wire _0559_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1100" *)
  wire _0560_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1101" *)
  wire _0561_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1113" *)
  wire _0562_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1114" *)
  wire _0563_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1115" *)
  wire _0564_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1116" *)
  wire _0565_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1128" *)
  wire _0566_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1129" *)
  wire _0567_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1130" *)
  wire _0568_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1131" *)
  wire _0569_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1143" *)
  wire _0570_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1144" *)
  wire _0571_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1145" *)
  wire _0572_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1146" *)
  wire _0573_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1158" *)
  wire _0574_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1159" *)
  wire _0575_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1160" *)
  wire _0576_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1161" *)
  wire _0577_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1173" *)
  wire _0578_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1174" *)
  wire _0579_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1175" *)
  wire _0580_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1176" *)
  wire _0581_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1188" *)
  wire _0582_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1189" *)
  wire _0583_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1190" *)
  wire _0584_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1191" *)
  wire _0585_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1203" *)
  wire _0586_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1204" *)
  wire _0587_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1205" *)
  wire _0588_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1206" *)
  wire _0589_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1218" *)
  wire _0590_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1219" *)
  wire _0591_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1220" *)
  wire _0592_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1221" *)
  wire _0593_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1233" *)
  wire _0594_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1234" *)
  wire _0595_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1235" *)
  wire _0596_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1236" *)
  wire _0597_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1248" *)
  wire _0598_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1249" *)
  wire _0599_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1250" *)
  wire _0600_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1251" *)
  wire _0601_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1263" *)
  wire _0602_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1264" *)
  wire _0603_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1265" *)
  wire _0604_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1266" *)
  wire _0605_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1278" *)
  wire _0606_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1279" *)
  wire _0607_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1280" *)
  wire _0608_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1281" *)
  wire _0609_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1293" *)
  wire _0610_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1294" *)
  wire _0611_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1295" *)
  wire _0612_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1296" *)
  wire _0613_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1308" *)
  wire _0614_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1309" *)
  wire _0615_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1310" *)
  wire _0616_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1311" *)
  wire _0617_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1323" *)
  wire _0618_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1324" *)
  wire _0619_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1325" *)
  wire _0620_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1326" *)
  wire _0621_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1344" *)
  wire [3:0] _0622_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1345" *)
  wire [3:0] _0623_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1346" *)
  wire [3:0] _0624_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1347" *)
  wire [3:0] _0625_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1365" *)
  wire [3:0] _0626_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1366" *)
  wire [3:0] _0627_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1367" *)
  wire [3:0] _0628_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1368" *)
  wire [3:0] _0629_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1386" *)
  wire [3:0] _0630_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1387" *)
  wire [3:0] _0631_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1388" *)
  wire [3:0] _0632_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1389" *)
  wire [3:0] _0633_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1407" *)
  wire [3:0] _0634_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1408" *)
  wire [3:0] _0635_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1409" *)
  wire [3:0] _0636_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1410" *)
  wire [3:0] _0637_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1428" *)
  wire [3:0] _0638_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1429" *)
  wire [3:0] _0639_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1430" *)
  wire [3:0] _0640_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1431" *)
  wire [3:0] _0641_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1449" *)
  wire [3:0] _0642_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1450" *)
  wire [3:0] _0643_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1451" *)
  wire [3:0] _0644_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1452" *)
  wire [3:0] _0645_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1470" *)
  wire [3:0] _0646_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1471" *)
  wire [3:0] _0647_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1472" *)
  wire [3:0] _0648_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1473" *)
  wire [3:0] _0649_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1491" *)
  wire [3:0] _0650_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1492" *)
  wire [3:0] _0651_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1493" *)
  wire [3:0] _0652_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1494" *)
  wire [3:0] _0653_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1512" *)
  wire [3:0] _0654_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1513" *)
  wire [3:0] _0655_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1514" *)
  wire [3:0] _0656_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1515" *)
  wire [3:0] _0657_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1533" *)
  wire [3:0] _0658_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1534" *)
  wire [3:0] _0659_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1535" *)
  wire [3:0] _0660_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1536" *)
  wire [3:0] _0661_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1554" *)
  wire [3:0] _0662_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1555" *)
  wire [3:0] _0663_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1556" *)
  wire [3:0] _0664_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1557" *)
  wire [3:0] _0665_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1575" *)
  wire [3:0] _0666_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1576" *)
  wire [3:0] _0667_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1577" *)
  wire [3:0] _0668_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1578" *)
  wire [3:0] _0669_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1596" *)
  wire [3:0] _0670_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1597" *)
  wire [3:0] _0671_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1598" *)
  wire [3:0] _0672_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1599" *)
  wire [3:0] _0673_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1617" *)
  wire [3:0] _0674_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1618" *)
  wire [3:0] _0675_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1619" *)
  wire [3:0] _0676_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1620" *)
  wire [3:0] _0677_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1638" *)
  wire [3:0] _0678_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1639" *)
  wire [3:0] _0679_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1640" *)
  wire [3:0] _0680_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1641" *)
  wire [3:0] _0681_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1659" *)
  wire [3:0] _0682_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1660" *)
  wire [3:0] _0683_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1661" *)
  wire [3:0] _0684_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1662" *)
  wire [3:0] _0685_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1680" *)
  wire [255:0] _0686_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1681" *)
  wire [255:0] _0687_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1682" *)
  wire [255:0] _0688_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1683" *)
  wire [255:0] _0689_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1701" *)
  wire [255:0] _0690_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1702" *)
  wire [255:0] _0691_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1703" *)
  wire [255:0] _0692_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1704" *)
  wire [255:0] _0693_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1722" *)
  wire [255:0] _0694_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1723" *)
  wire [255:0] _0695_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1724" *)
  wire [255:0] _0696_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1725" *)
  wire [255:0] _0697_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1743" *)
  wire [255:0] _0698_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1744" *)
  wire [255:0] _0699_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1745" *)
  wire [255:0] _0700_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1746" *)
  wire [255:0] _0701_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1764" *)
  wire [255:0] _0702_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1765" *)
  wire [255:0] _0703_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1766" *)
  wire [255:0] _0704_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1767" *)
  wire [255:0] _0705_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1785" *)
  wire [255:0] _0706_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1786" *)
  wire [255:0] _0707_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1787" *)
  wire [255:0] _0708_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1788" *)
  wire [255:0] _0709_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1806" *)
  wire [255:0] _0710_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1807" *)
  wire [255:0] _0711_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1808" *)
  wire [255:0] _0712_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1809" *)
  wire [255:0] _0713_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1827" *)
  wire [255:0] _0714_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1828" *)
  wire [255:0] _0715_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1829" *)
  wire [255:0] _0716_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1830" *)
  wire [255:0] _0717_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1848" *)
  wire [255:0] _0718_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1849" *)
  wire [255:0] _0719_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1850" *)
  wire [255:0] _0720_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1851" *)
  wire [255:0] _0721_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1869" *)
  wire [255:0] _0722_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1870" *)
  wire [255:0] _0723_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1871" *)
  wire [255:0] _0724_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1872" *)
  wire [255:0] _0725_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1890" *)
  wire [255:0] _0726_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1891" *)
  wire [255:0] _0727_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1892" *)
  wire [255:0] _0728_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1893" *)
  wire [255:0] _0729_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1911" *)
  wire [255:0] _0730_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1912" *)
  wire [255:0] _0731_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1913" *)
  wire [255:0] _0732_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1914" *)
  wire [255:0] _0733_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1932" *)
  wire [255:0] _0734_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1933" *)
  wire [255:0] _0735_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1934" *)
  wire [255:0] _0736_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1935" *)
  wire [255:0] _0737_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1953" *)
  wire [255:0] _0738_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1954" *)
  wire [255:0] _0739_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1955" *)
  wire [255:0] _0740_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1956" *)
  wire [255:0] _0741_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1974" *)
  wire [255:0] _0742_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1975" *)
  wire [255:0] _0743_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1976" *)
  wire [255:0] _0744_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1977" *)
  wire [255:0] _0745_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1995" *)
  wire [255:0] _0746_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1996" *)
  wire [255:0] _0747_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1997" *)
  wire [255:0] _0748_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1998" *)
  wire [255:0] _0749_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2754" *)
  wire _0750_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2761" *)
  wire _0751_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2768" *)
  wire _0752_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2775" *)
  wire _0753_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2782" *)
  wire _0754_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2789" *)
  wire _0755_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2796" *)
  wire _0756_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2803" *)
  wire _0757_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2810" *)
  wire _0758_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2817" *)
  wire _0759_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2824" *)
  wire _0760_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2831" *)
  wire _0761_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2838" *)
  wire _0762_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2845" *)
  wire _0763_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2852" *)
  wire _0764_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2859" *)
  wire _0765_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2866" *)
  wire _0766_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2873" *)
  wire _0767_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2880" *)
  wire _0768_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2887" *)
  wire _0769_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2894" *)
  wire _0770_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2901" *)
  wire _0771_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2908" *)
  wire _0772_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2915" *)
  wire _0773_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2922" *)
  wire _0774_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2929" *)
  wire _0775_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2936" *)
  wire _0776_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2943" *)
  wire _0777_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2950" *)
  wire _0778_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2957" *)
  wire _0779_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2964" *)
  wire _0780_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2971" *)
  wire _0781_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3090" *)
  wire [3:0] _0782_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3091" *)
  wire [3:0] _0783_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3092" *)
  wire [3:0] _0784_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3093" *)
  wire [3:0] _0785_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3111" *)
  wire [3:0] _0786_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3112" *)
  wire [3:0] _0787_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3113" *)
  wire [3:0] _0788_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3114" *)
  wire [3:0] _0789_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3132" *)
  wire [3:0] _0790_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3133" *)
  wire [3:0] _0791_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3134" *)
  wire [3:0] _0792_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3135" *)
  wire [3:0] _0793_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3153" *)
  wire [3:0] _0794_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3154" *)
  wire [3:0] _0795_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3155" *)
  wire [3:0] _0796_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3156" *)
  wire [3:0] _0797_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3174" *)
  wire [3:0] _0798_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3175" *)
  wire [3:0] _0799_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3176" *)
  wire [3:0] _0800_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3177" *)
  wire [3:0] _0801_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3195" *)
  wire [3:0] _0802_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3196" *)
  wire [3:0] _0803_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3197" *)
  wire [3:0] _0804_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3198" *)
  wire [3:0] _0805_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3216" *)
  wire [3:0] _0806_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3217" *)
  wire [3:0] _0807_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3218" *)
  wire [3:0] _0808_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3219" *)
  wire [3:0] _0809_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3237" *)
  wire [3:0] _0810_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3238" *)
  wire [3:0] _0811_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3239" *)
  wire [3:0] _0812_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3240" *)
  wire [3:0] _0813_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3258" *)
  wire [3:0] _0814_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3259" *)
  wire [3:0] _0815_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3260" *)
  wire [3:0] _0816_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3261" *)
  wire [3:0] _0817_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3279" *)
  wire [3:0] _0818_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3280" *)
  wire [3:0] _0819_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3281" *)
  wire [3:0] _0820_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3282" *)
  wire [3:0] _0821_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3300" *)
  wire [3:0] _0822_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3301" *)
  wire [3:0] _0823_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3302" *)
  wire [3:0] _0824_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3303" *)
  wire [3:0] _0825_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3321" *)
  wire [3:0] _0826_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3322" *)
  wire [3:0] _0827_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3323" *)
  wire [3:0] _0828_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3324" *)
  wire [3:0] _0829_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3342" *)
  wire [3:0] _0830_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3343" *)
  wire [3:0] _0831_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3344" *)
  wire [3:0] _0832_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3345" *)
  wire [3:0] _0833_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3363" *)
  wire [3:0] _0834_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3364" *)
  wire [3:0] _0835_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3365" *)
  wire [3:0] _0836_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3366" *)
  wire [3:0] _0837_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3384" *)
  wire [3:0] _0838_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3385" *)
  wire [3:0] _0839_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3386" *)
  wire [3:0] _0840_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3387" *)
  wire [3:0] _0841_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3405" *)
  wire [3:0] _0842_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3406" *)
  wire [3:0] _0843_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3407" *)
  wire [3:0] _0844_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3408" *)
  wire [3:0] _0845_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3802" *)
  wire _0846_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3809" *)
  wire _0847_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3850" *)
  wire [255:0] _0848_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3851" *)
  wire [255:0] _0849_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3852" *)
  wire [255:0] _0850_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3853" *)
  wire [255:0] _0851_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3854" *)
  wire [255:0] _0852_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3855" *)
  wire [255:0] _0853_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3856" *)
  wire [255:0] _0854_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3857" *)
  wire [255:0] _0855_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3858" *)
  wire [255:0] _0856_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3859" *)
  wire [255:0] _0857_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3860" *)
  wire [255:0] _0858_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3861" *)
  wire [255:0] _0859_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3862" *)
  wire [255:0] _0860_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3863" *)
  wire [255:0] _0861_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3901" *)
  wire [255:0] _0862_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3902" *)
  wire [255:0] _0863_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3903" *)
  wire [255:0] _0864_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3904" *)
  wire [255:0] _0865_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3905" *)
  wire [255:0] _0866_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3906" *)
  wire [255:0] _0867_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3907" *)
  wire [255:0] _0868_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3908" *)
  wire [255:0] _0869_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3909" *)
  wire [255:0] _0870_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3910" *)
  wire [255:0] _0871_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3911" *)
  wire [255:0] _0872_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3912" *)
  wire [255:0] _0873_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3913" *)
  wire [255:0] _0874_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3914" *)
  wire [255:0] _0875_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3928" *)
  wire [255:0] _0876_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3929" *)
  wire [255:0] _0877_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3943" *)
  wire [255:0] _0878_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3944" *)
  wire [255:0] _0879_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3958" *)
  wire [255:0] _0880_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3959" *)
  wire [255:0] _0881_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3973" *)
  wire [255:0] _0882_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3974" *)
  wire [255:0] _0883_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3988" *)
  wire [255:0] _0884_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3989" *)
  wire [255:0] _0885_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4003" *)
  wire [255:0] _0886_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4004" *)
  wire [255:0] _0887_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4018" *)
  wire [255:0] _0888_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4019" *)
  wire [255:0] _0889_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4033" *)
  wire [255:0] _0890_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4034" *)
  wire [255:0] _0891_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4048" *)
  wire [255:0] _0892_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4049" *)
  wire [255:0] _0893_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4063" *)
  wire [255:0] _0894_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4064" *)
  wire [255:0] _0895_;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:75" *)
  input [7:0] dc2sbuf_p0_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:92" *)
  wire [3:0] dc2sbuf_p0_rd_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:76" *)
  output [255:0] dc2sbuf_p0_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:74" *)
  input dc2sbuf_p0_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:93" *)
  wire [3:0] dc2sbuf_p0_rd_esel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:126" *)
  wire dc2sbuf_p0_rd_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:127" *)
  wire dc2sbuf_p0_rd_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:128" *)
  wire dc2sbuf_p0_rd_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:129" *)
  wire dc2sbuf_p0_rd_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:130" *)
  wire dc2sbuf_p0_rd_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:131" *)
  wire dc2sbuf_p0_rd_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:132" *)
  wire dc2sbuf_p0_rd_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:133" *)
  wire dc2sbuf_p0_rd_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:134" *)
  wire dc2sbuf_p0_rd_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:135" *)
  wire dc2sbuf_p0_rd_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:136" *)
  wire dc2sbuf_p0_rd_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:137" *)
  wire dc2sbuf_p0_rd_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:138" *)
  wire dc2sbuf_p0_rd_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:139" *)
  wire dc2sbuf_p0_rd_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:140" *)
  wire dc2sbuf_p0_rd_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:141" *)
  wire dc2sbuf_p0_rd_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:57" *)
  input [7:0] dc2sbuf_p0_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:94" *)
  wire [3:0] dc2sbuf_p0_wr_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:58" *)
  input [255:0] dc2sbuf_p0_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:56" *)
  input dc2sbuf_p0_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:142" *)
  wire dc2sbuf_p0_wr_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:143" *)
  wire dc2sbuf_p0_wr_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:144" *)
  wire dc2sbuf_p0_wr_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:145" *)
  wire dc2sbuf_p0_wr_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:146" *)
  wire dc2sbuf_p0_wr_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:147" *)
  wire dc2sbuf_p0_wr_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:148" *)
  wire dc2sbuf_p0_wr_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:149" *)
  wire dc2sbuf_p0_wr_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:150" *)
  wire dc2sbuf_p0_wr_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:151" *)
  wire dc2sbuf_p0_wr_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:152" *)
  wire dc2sbuf_p0_wr_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:153" *)
  wire dc2sbuf_p0_wr_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:154" *)
  wire dc2sbuf_p0_wr_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:155" *)
  wire dc2sbuf_p0_wr_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:156" *)
  wire dc2sbuf_p0_wr_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:157" *)
  wire dc2sbuf_p0_wr_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:78" *)
  input [7:0] dc2sbuf_p1_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:95" *)
  wire [3:0] dc2sbuf_p1_rd_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:79" *)
  output [255:0] dc2sbuf_p1_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:77" *)
  input dc2sbuf_p1_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:96" *)
  wire [3:0] dc2sbuf_p1_rd_esel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:158" *)
  wire dc2sbuf_p1_rd_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:159" *)
  wire dc2sbuf_p1_rd_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:160" *)
  wire dc2sbuf_p1_rd_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:161" *)
  wire dc2sbuf_p1_rd_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:162" *)
  wire dc2sbuf_p1_rd_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:163" *)
  wire dc2sbuf_p1_rd_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:164" *)
  wire dc2sbuf_p1_rd_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:165" *)
  wire dc2sbuf_p1_rd_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:166" *)
  wire dc2sbuf_p1_rd_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:167" *)
  wire dc2sbuf_p1_rd_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:168" *)
  wire dc2sbuf_p1_rd_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:169" *)
  wire dc2sbuf_p1_rd_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:170" *)
  wire dc2sbuf_p1_rd_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:171" *)
  wire dc2sbuf_p1_rd_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:172" *)
  wire dc2sbuf_p1_rd_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:173" *)
  wire dc2sbuf_p1_rd_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:60" *)
  input [7:0] dc2sbuf_p1_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:97" *)
  wire [3:0] dc2sbuf_p1_wr_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:61" *)
  input [255:0] dc2sbuf_p1_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:59" *)
  input dc2sbuf_p1_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:174" *)
  wire dc2sbuf_p1_wr_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:175" *)
  wire dc2sbuf_p1_wr_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:176" *)
  wire dc2sbuf_p1_wr_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:177" *)
  wire dc2sbuf_p1_wr_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:178" *)
  wire dc2sbuf_p1_wr_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:179" *)
  wire dc2sbuf_p1_wr_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:180" *)
  wire dc2sbuf_p1_wr_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:181" *)
  wire dc2sbuf_p1_wr_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:182" *)
  wire dc2sbuf_p1_wr_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:183" *)
  wire dc2sbuf_p1_wr_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:184" *)
  wire dc2sbuf_p1_wr_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:185" *)
  wire dc2sbuf_p1_wr_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:186" *)
  wire dc2sbuf_p1_wr_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:187" *)
  wire dc2sbuf_p1_wr_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:188" *)
  wire dc2sbuf_p1_wr_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:189" *)
  wire dc2sbuf_p1_wr_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:87" *)
  input [7:0] img2sbuf_p0_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:98" *)
  wire [3:0] img2sbuf_p0_rd_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:88" *)
  output [255:0] img2sbuf_p0_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:86" *)
  input img2sbuf_p0_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:99" *)
  wire [3:0] img2sbuf_p0_rd_esel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:190" *)
  wire img2sbuf_p0_rd_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:191" *)
  wire img2sbuf_p0_rd_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:192" *)
  wire img2sbuf_p0_rd_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:193" *)
  wire img2sbuf_p0_rd_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:194" *)
  wire img2sbuf_p0_rd_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:195" *)
  wire img2sbuf_p0_rd_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:196" *)
  wire img2sbuf_p0_rd_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:197" *)
  wire img2sbuf_p0_rd_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:198" *)
  wire img2sbuf_p0_rd_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:199" *)
  wire img2sbuf_p0_rd_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:200" *)
  wire img2sbuf_p0_rd_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:201" *)
  wire img2sbuf_p0_rd_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:202" *)
  wire img2sbuf_p0_rd_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:203" *)
  wire img2sbuf_p0_rd_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:204" *)
  wire img2sbuf_p0_rd_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:205" *)
  wire img2sbuf_p0_rd_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:69" *)
  input [7:0] img2sbuf_p0_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:100" *)
  wire [3:0] img2sbuf_p0_wr_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:70" *)
  input [255:0] img2sbuf_p0_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:68" *)
  input img2sbuf_p0_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:206" *)
  wire img2sbuf_p0_wr_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:207" *)
  wire img2sbuf_p0_wr_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:208" *)
  wire img2sbuf_p0_wr_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:209" *)
  wire img2sbuf_p0_wr_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:210" *)
  wire img2sbuf_p0_wr_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:211" *)
  wire img2sbuf_p0_wr_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:212" *)
  wire img2sbuf_p0_wr_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:213" *)
  wire img2sbuf_p0_wr_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:214" *)
  wire img2sbuf_p0_wr_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:215" *)
  wire img2sbuf_p0_wr_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:216" *)
  wire img2sbuf_p0_wr_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:217" *)
  wire img2sbuf_p0_wr_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:218" *)
  wire img2sbuf_p0_wr_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:219" *)
  wire img2sbuf_p0_wr_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:220" *)
  wire img2sbuf_p0_wr_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:221" *)
  wire img2sbuf_p0_wr_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:90" *)
  input [7:0] img2sbuf_p1_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:101" *)
  wire [3:0] img2sbuf_p1_rd_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:91" *)
  output [255:0] img2sbuf_p1_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:89" *)
  input img2sbuf_p1_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:102" *)
  wire [3:0] img2sbuf_p1_rd_esel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:222" *)
  wire img2sbuf_p1_rd_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:223" *)
  wire img2sbuf_p1_rd_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:224" *)
  wire img2sbuf_p1_rd_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:225" *)
  wire img2sbuf_p1_rd_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:226" *)
  wire img2sbuf_p1_rd_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:227" *)
  wire img2sbuf_p1_rd_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:228" *)
  wire img2sbuf_p1_rd_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:229" *)
  wire img2sbuf_p1_rd_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:230" *)
  wire img2sbuf_p1_rd_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:231" *)
  wire img2sbuf_p1_rd_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:232" *)
  wire img2sbuf_p1_rd_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:233" *)
  wire img2sbuf_p1_rd_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:234" *)
  wire img2sbuf_p1_rd_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:235" *)
  wire img2sbuf_p1_rd_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:236" *)
  wire img2sbuf_p1_rd_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:237" *)
  wire img2sbuf_p1_rd_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:72" *)
  input [7:0] img2sbuf_p1_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:103" *)
  wire [3:0] img2sbuf_p1_wr_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:73" *)
  input [255:0] img2sbuf_p1_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:71" *)
  input img2sbuf_p1_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:238" *)
  wire img2sbuf_p1_wr_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:239" *)
  wire img2sbuf_p1_wr_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:240" *)
  wire img2sbuf_p1_wr_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:241" *)
  wire img2sbuf_p1_wr_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:242" *)
  wire img2sbuf_p1_wr_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:243" *)
  wire img2sbuf_p1_wr_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:244" *)
  wire img2sbuf_p1_wr_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:245" *)
  wire img2sbuf_p1_wr_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:246" *)
  wire img2sbuf_p1_wr_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:247" *)
  wire img2sbuf_p1_wr_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:248" *)
  wire img2sbuf_p1_wr_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:249" *)
  wire img2sbuf_p1_wr_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:250" *)
  wire img2sbuf_p1_wr_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:251" *)
  wire img2sbuf_p1_wr_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:252" *)
  wire img2sbuf_p1_wr_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:253" *)
  wire img2sbuf_p1_wr_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:53" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:54" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:55" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:254" *)
  wire [255:0] sbuf_p0_norm_rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:255" *)
  reg sbuf_p0_rd_en_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:256" *)
  wire [255:0] sbuf_p0_rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:257" *)
  reg [255:0] sbuf_p0_rdat_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:258" *)
  wire sbuf_p0_re_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:259" *)
  reg sbuf_p0_re_00_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:260" *)
  reg sbuf_p0_re_00_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:261" *)
  wire sbuf_p0_re_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:262" *)
  reg sbuf_p0_re_01_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:263" *)
  reg sbuf_p0_re_01_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:264" *)
  wire sbuf_p0_re_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:265" *)
  reg sbuf_p0_re_02_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:266" *)
  reg sbuf_p0_re_02_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:267" *)
  wire sbuf_p0_re_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:268" *)
  reg sbuf_p0_re_03_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:269" *)
  reg sbuf_p0_re_03_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:270" *)
  wire sbuf_p0_re_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:271" *)
  reg sbuf_p0_re_04_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:272" *)
  wire sbuf_p0_re_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:273" *)
  reg sbuf_p0_re_05_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:274" *)
  wire sbuf_p0_re_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:275" *)
  reg sbuf_p0_re_06_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:276" *)
  wire sbuf_p0_re_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:277" *)
  reg sbuf_p0_re_07_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:278" *)
  wire sbuf_p0_re_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:279" *)
  reg sbuf_p0_re_08_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:280" *)
  wire sbuf_p0_re_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:281" *)
  reg sbuf_p0_re_09_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:282" *)
  wire sbuf_p0_re_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:283" *)
  reg sbuf_p0_re_10_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:284" *)
  wire sbuf_p0_re_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:285" *)
  reg sbuf_p0_re_11_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:286" *)
  wire sbuf_p0_re_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:287" *)
  reg sbuf_p0_re_12_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:288" *)
  wire sbuf_p0_re_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:289" *)
  reg sbuf_p0_re_13_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:290" *)
  wire sbuf_p0_re_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:291" *)
  reg sbuf_p0_re_14_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:292" *)
  wire sbuf_p0_re_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:293" *)
  reg sbuf_p0_re_15_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:294" *)
  wire [255:0] sbuf_p0_wg_rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:295" *)
  wire [255:0] sbuf_p0_wg_rdat_src_0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:296" *)
  wire [255:0] sbuf_p0_wg_rdat_src_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:297" *)
  wire [255:0] sbuf_p0_wg_rdat_src_2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:298" *)
  wire [255:0] sbuf_p0_wg_rdat_src_3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:299" *)
  wire sbuf_p0_wg_sel_q0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:300" *)
  reg sbuf_p0_wg_sel_q0_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:301" *)
  wire sbuf_p0_wg_sel_q1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:302" *)
  reg sbuf_p0_wg_sel_q1_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:303" *)
  wire sbuf_p0_wg_sel_q2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:304" *)
  reg sbuf_p0_wg_sel_q2_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:305" *)
  wire sbuf_p0_wg_sel_q3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:306" *)
  reg sbuf_p0_wg_sel_q3_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:307" *)
  wire [255:0] sbuf_p1_norm_rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:308" *)
  reg sbuf_p1_rd_en_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:309" *)
  wire [255:0] sbuf_p1_rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:310" *)
  reg [255:0] sbuf_p1_rdat_d2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:311" *)
  wire sbuf_p1_re_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:312" *)
  reg sbuf_p1_re_00_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:313" *)
  reg sbuf_p1_re_00_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:314" *)
  wire sbuf_p1_re_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:315" *)
  reg sbuf_p1_re_01_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:316" *)
  reg sbuf_p1_re_01_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:317" *)
  wire sbuf_p1_re_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:318" *)
  reg sbuf_p1_re_02_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:319" *)
  reg sbuf_p1_re_02_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:320" *)
  wire sbuf_p1_re_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:321" *)
  reg sbuf_p1_re_03_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:322" *)
  reg sbuf_p1_re_03_wg_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:323" *)
  wire sbuf_p1_re_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:324" *)
  reg sbuf_p1_re_04_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:325" *)
  wire sbuf_p1_re_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:326" *)
  reg sbuf_p1_re_05_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:327" *)
  wire sbuf_p1_re_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:328" *)
  reg sbuf_p1_re_06_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:329" *)
  wire sbuf_p1_re_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:330" *)
  reg sbuf_p1_re_07_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:331" *)
  wire sbuf_p1_re_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:332" *)
  reg sbuf_p1_re_08_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:333" *)
  wire sbuf_p1_re_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:334" *)
  reg sbuf_p1_re_09_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:335" *)
  wire sbuf_p1_re_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:336" *)
  reg sbuf_p1_re_10_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:337" *)
  wire sbuf_p1_re_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:338" *)
  reg sbuf_p1_re_11_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:339" *)
  wire sbuf_p1_re_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:340" *)
  reg sbuf_p1_re_12_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:341" *)
  wire sbuf_p1_re_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:342" *)
  reg sbuf_p1_re_13_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:343" *)
  wire sbuf_p1_re_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:344" *)
  reg sbuf_p1_re_14_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:345" *)
  wire sbuf_p1_re_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:346" *)
  reg sbuf_p1_re_15_norm_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:347" *)
  wire [255:0] sbuf_p1_wg_rdat;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:348" *)
  wire [255:0] sbuf_p1_wg_rdat_src_0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:349" *)
  wire [255:0] sbuf_p1_wg_rdat_src_1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:350" *)
  wire [255:0] sbuf_p1_wg_rdat_src_2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:351" *)
  wire [255:0] sbuf_p1_wg_rdat_src_3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:352" *)
  wire sbuf_p1_wg_sel_q0;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:353" *)
  reg sbuf_p1_wg_sel_q0_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:354" *)
  wire sbuf_p1_wg_sel_q1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:355" *)
  reg sbuf_p1_wg_sel_q1_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:356" *)
  wire sbuf_p1_wg_sel_q2;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:357" *)
  reg sbuf_p1_wg_sel_q2_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:358" *)
  wire sbuf_p1_wg_sel_q3;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:359" *)
  reg sbuf_p1_wg_sel_q3_d1;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:360" *)
  wire [3:0] sbuf_ra_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:361" *)
  wire [3:0] sbuf_ra_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:362" *)
  wire [3:0] sbuf_ra_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:363" *)
  wire [3:0] sbuf_ra_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:364" *)
  wire [3:0] sbuf_ra_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:365" *)
  wire [3:0] sbuf_ra_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:366" *)
  wire [3:0] sbuf_ra_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:367" *)
  wire [3:0] sbuf_ra_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:368" *)
  wire [3:0] sbuf_ra_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:369" *)
  wire [3:0] sbuf_ra_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:370" *)
  wire [3:0] sbuf_ra_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:371" *)
  wire [3:0] sbuf_ra_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:372" *)
  wire [3:0] sbuf_ra_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:373" *)
  wire [3:0] sbuf_ra_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:374" *)
  wire [3:0] sbuf_ra_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:375" *)
  wire [3:0] sbuf_ra_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:104" *)
  wire [255:0] sbuf_rdat_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:105" *)
  wire [255:0] sbuf_rdat_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:106" *)
  wire [255:0] sbuf_rdat_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:107" *)
  wire [255:0] sbuf_rdat_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:108" *)
  wire [255:0] sbuf_rdat_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:109" *)
  wire [255:0] sbuf_rdat_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:110" *)
  wire [255:0] sbuf_rdat_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:111" *)
  wire [255:0] sbuf_rdat_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:112" *)
  wire [255:0] sbuf_rdat_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:113" *)
  wire [255:0] sbuf_rdat_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:114" *)
  wire [255:0] sbuf_rdat_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:115" *)
  wire [255:0] sbuf_rdat_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:116" *)
  wire [255:0] sbuf_rdat_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:117" *)
  wire [255:0] sbuf_rdat_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:118" *)
  wire [255:0] sbuf_rdat_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:119" *)
  wire [255:0] sbuf_rdat_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:376" *)
  wire sbuf_re_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:377" *)
  wire sbuf_re_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:378" *)
  wire sbuf_re_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:379" *)
  wire sbuf_re_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:380" *)
  wire sbuf_re_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:381" *)
  wire sbuf_re_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:382" *)
  wire sbuf_re_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:383" *)
  wire sbuf_re_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:384" *)
  wire sbuf_re_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:385" *)
  wire sbuf_re_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:386" *)
  wire sbuf_re_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:387" *)
  wire sbuf_re_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:388" *)
  wire sbuf_re_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:389" *)
  wire sbuf_re_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:390" *)
  wire sbuf_re_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:391" *)
  wire sbuf_re_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:392" *)
  wire [3:0] sbuf_wa_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:393" *)
  wire [3:0] sbuf_wa_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:394" *)
  wire [3:0] sbuf_wa_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:395" *)
  wire [3:0] sbuf_wa_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:396" *)
  wire [3:0] sbuf_wa_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:397" *)
  wire [3:0] sbuf_wa_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:398" *)
  wire [3:0] sbuf_wa_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:399" *)
  wire [3:0] sbuf_wa_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:400" *)
  wire [3:0] sbuf_wa_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:401" *)
  wire [3:0] sbuf_wa_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:402" *)
  wire [3:0] sbuf_wa_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:403" *)
  wire [3:0] sbuf_wa_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:404" *)
  wire [3:0] sbuf_wa_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:405" *)
  wire [3:0] sbuf_wa_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:406" *)
  wire [3:0] sbuf_wa_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:407" *)
  wire [3:0] sbuf_wa_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:408" *)
  wire [255:0] sbuf_wdat_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:409" *)
  wire [255:0] sbuf_wdat_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:410" *)
  wire [255:0] sbuf_wdat_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:411" *)
  wire [255:0] sbuf_wdat_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:412" *)
  wire [255:0] sbuf_wdat_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:413" *)
  wire [255:0] sbuf_wdat_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:414" *)
  wire [255:0] sbuf_wdat_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:415" *)
  wire [255:0] sbuf_wdat_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:416" *)
  wire [255:0] sbuf_wdat_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:417" *)
  wire [255:0] sbuf_wdat_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:418" *)
  wire [255:0] sbuf_wdat_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:419" *)
  wire [255:0] sbuf_wdat_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:420" *)
  wire [255:0] sbuf_wdat_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:421" *)
  wire [255:0] sbuf_wdat_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:422" *)
  wire [255:0] sbuf_wdat_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:423" *)
  wire [255:0] sbuf_wdat_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:424" *)
  wire sbuf_we_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:425" *)
  wire sbuf_we_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:426" *)
  wire sbuf_we_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:427" *)
  wire sbuf_we_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:428" *)
  wire sbuf_we_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:429" *)
  wire sbuf_we_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:430" *)
  wire sbuf_we_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:431" *)
  wire sbuf_we_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:432" *)
  wire sbuf_we_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:433" *)
  wire sbuf_we_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:434" *)
  wire sbuf_we_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:435" *)
  wire sbuf_we_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:436" *)
  wire sbuf_we_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:437" *)
  wire sbuf_we_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:438" *)
  wire sbuf_we_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:439" *)
  wire sbuf_we_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:81" *)
  input [7:0] wg2sbuf_p0_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:120" *)
  wire [1:0] wg2sbuf_p0_rd_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:82" *)
  output [255:0] wg2sbuf_p0_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:80" *)
  input wg2sbuf_p0_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:121" *)
  wire [3:0] wg2sbuf_p0_rd_esel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:440" *)
  wire wg2sbuf_p0_rd_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:441" *)
  wire wg2sbuf_p0_rd_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:442" *)
  wire wg2sbuf_p0_rd_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:443" *)
  wire wg2sbuf_p0_rd_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:444" *)
  wire wg2sbuf_p0_rd_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:445" *)
  wire wg2sbuf_p0_rd_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:446" *)
  wire wg2sbuf_p0_rd_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:447" *)
  wire wg2sbuf_p0_rd_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:448" *)
  wire wg2sbuf_p0_rd_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:449" *)
  wire wg2sbuf_p0_rd_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:450" *)
  wire wg2sbuf_p0_rd_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:451" *)
  wire wg2sbuf_p0_rd_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:452" *)
  wire wg2sbuf_p0_rd_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:453" *)
  wire wg2sbuf_p0_rd_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:454" *)
  wire wg2sbuf_p0_rd_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:455" *)
  wire wg2sbuf_p0_rd_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:63" *)
  input [7:0] wg2sbuf_p0_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:122" *)
  wire [3:0] wg2sbuf_p0_wr_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:64" *)
  input [255:0] wg2sbuf_p0_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:62" *)
  input wg2sbuf_p0_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:456" *)
  wire wg2sbuf_p0_wr_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:457" *)
  wire wg2sbuf_p0_wr_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:458" *)
  wire wg2sbuf_p0_wr_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:459" *)
  wire wg2sbuf_p0_wr_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:460" *)
  wire wg2sbuf_p0_wr_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:461" *)
  wire wg2sbuf_p0_wr_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:462" *)
  wire wg2sbuf_p0_wr_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:463" *)
  wire wg2sbuf_p0_wr_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:464" *)
  wire wg2sbuf_p0_wr_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:465" *)
  wire wg2sbuf_p0_wr_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:466" *)
  wire wg2sbuf_p0_wr_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:467" *)
  wire wg2sbuf_p0_wr_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:468" *)
  wire wg2sbuf_p0_wr_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:469" *)
  wire wg2sbuf_p0_wr_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:470" *)
  wire wg2sbuf_p0_wr_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:471" *)
  wire wg2sbuf_p0_wr_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:84" *)
  input [7:0] wg2sbuf_p1_rd_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:123" *)
  wire [1:0] wg2sbuf_p1_rd_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:85" *)
  output [255:0] wg2sbuf_p1_rd_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:83" *)
  input wg2sbuf_p1_rd_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:124" *)
  wire [3:0] wg2sbuf_p1_rd_esel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:472" *)
  wire wg2sbuf_p1_rd_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:473" *)
  wire wg2sbuf_p1_rd_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:474" *)
  wire wg2sbuf_p1_rd_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:475" *)
  wire wg2sbuf_p1_rd_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:476" *)
  wire wg2sbuf_p1_rd_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:477" *)
  wire wg2sbuf_p1_rd_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:478" *)
  wire wg2sbuf_p1_rd_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:479" *)
  wire wg2sbuf_p1_rd_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:480" *)
  wire wg2sbuf_p1_rd_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:481" *)
  wire wg2sbuf_p1_rd_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:482" *)
  wire wg2sbuf_p1_rd_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:483" *)
  wire wg2sbuf_p1_rd_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:484" *)
  wire wg2sbuf_p1_rd_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:485" *)
  wire wg2sbuf_p1_rd_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:486" *)
  wire wg2sbuf_p1_rd_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:487" *)
  wire wg2sbuf_p1_rd_sel_15;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:66" *)
  input [7:0] wg2sbuf_p1_wr_addr;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:125" *)
  wire [3:0] wg2sbuf_p1_wr_bsel;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:67" *)
  input [255:0] wg2sbuf_p1_wr_data;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:65" *)
  input wg2sbuf_p1_wr_en;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:488" *)
  wire wg2sbuf_p1_wr_sel_00;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:489" *)
  wire wg2sbuf_p1_wr_sel_01;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:490" *)
  wire wg2sbuf_p1_wr_sel_02;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:491" *)
  wire wg2sbuf_p1_wr_sel_03;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:492" *)
  wire wg2sbuf_p1_wr_sel_04;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:493" *)
  wire wg2sbuf_p1_wr_sel_05;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:494" *)
  wire wg2sbuf_p1_wr_sel_06;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:495" *)
  wire wg2sbuf_p1_wr_sel_07;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:496" *)
  wire wg2sbuf_p1_wr_sel_08;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:497" *)
  wire wg2sbuf_p1_wr_sel_09;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:498" *)
  wire wg2sbuf_p1_wr_sel_10;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:499" *)
  wire wg2sbuf_p1_wr_sel_11;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:500" *)
  wire wg2sbuf_p1_wr_sel_12;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:501" *)
  wire wg2sbuf_p1_wr_sel_13;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:502" *)
  wire wg2sbuf_p1_wr_sel_14;
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:503" *)
  wire wg2sbuf_p1_wr_sel_15;
  assign wg2sbuf_p1_wr_sel_13 = _0380_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1003" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_13 = _0381_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1009" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_13 = _0382_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1015" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_14 = _0383_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1021" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_14 = _0384_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1027" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_14 = _0385_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1033" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_14 = _0386_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1039" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_14 = _0387_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1045" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_14 = _0388_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1051" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_15 = _0389_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1057" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_15 = _0390_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1063" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_15 = _0391_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1069" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_15 = _0392_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1075" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_15 = _0393_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1081" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_15 = _0394_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1087" *) img2sbuf_p1_wr_en;
  assign _0044_ = { dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1343" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0045_ = { dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1344" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0046_ = { wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1345" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0047_ = { wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1346" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0048_ = { img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1347" *) img2sbuf_p0_wr_addr[3:0];
  assign _0049_ = { img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1348" *) img2sbuf_p1_wr_addr[3:0];
  assign _0050_ = { dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1364" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0051_ = { dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1365" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0052_ = { wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1366" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0053_ = { wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1367" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0054_ = { img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1368" *) img2sbuf_p0_wr_addr[3:0];
  assign _0055_ = { img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1369" *) img2sbuf_p1_wr_addr[3:0];
  assign _0056_ = { dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1385" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0057_ = { dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1386" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0058_ = { wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1387" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0059_ = { wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1388" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0060_ = { img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1389" *) img2sbuf_p0_wr_addr[3:0];
  assign _0061_ = { img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1390" *) img2sbuf_p1_wr_addr[3:0];
  assign _0062_ = { dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1406" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0063_ = { dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1407" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0064_ = { wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1408" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0065_ = { wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1409" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0066_ = { img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1410" *) img2sbuf_p0_wr_addr[3:0];
  assign _0067_ = { img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1411" *) img2sbuf_p1_wr_addr[3:0];
  assign _0068_ = { dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1427" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0069_ = { dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1428" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0070_ = { wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1429" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0071_ = { wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1430" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0072_ = { img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1431" *) img2sbuf_p0_wr_addr[3:0];
  assign _0073_ = { img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1432" *) img2sbuf_p1_wr_addr[3:0];
  assign _0074_ = { dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1448" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0075_ = { dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1449" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0076_ = { wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1450" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0077_ = { wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1451" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0078_ = { img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1452" *) img2sbuf_p0_wr_addr[3:0];
  assign _0079_ = { img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1453" *) img2sbuf_p1_wr_addr[3:0];
  assign _0080_ = { dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1469" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0081_ = { dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1470" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0082_ = { wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1471" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0083_ = { wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1472" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0084_ = { img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1473" *) img2sbuf_p0_wr_addr[3:0];
  assign _0085_ = { img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1474" *) img2sbuf_p1_wr_addr[3:0];
  assign _0086_ = { dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1490" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0087_ = { dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1491" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0088_ = { wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1492" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0089_ = { wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1493" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0090_ = { img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1494" *) img2sbuf_p0_wr_addr[3:0];
  assign _0091_ = { img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1495" *) img2sbuf_p1_wr_addr[3:0];
  assign _0092_ = { dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1511" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0093_ = { dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1512" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0094_ = { wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1513" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0095_ = { wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1514" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0096_ = { img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1515" *) img2sbuf_p0_wr_addr[3:0];
  assign _0097_ = { img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1516" *) img2sbuf_p1_wr_addr[3:0];
  assign _0098_ = { dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1532" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0099_ = { dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1533" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0100_ = { wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1534" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0101_ = { wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1535" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0102_ = { img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1536" *) img2sbuf_p0_wr_addr[3:0];
  assign _0103_ = { img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1537" *) img2sbuf_p1_wr_addr[3:0];
  assign _0104_ = { dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1553" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0105_ = { dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1554" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0106_ = { wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1555" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0107_ = { wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1556" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0108_ = { img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1557" *) img2sbuf_p0_wr_addr[3:0];
  assign _0109_ = { img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1558" *) img2sbuf_p1_wr_addr[3:0];
  assign _0110_ = { dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1574" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0111_ = { dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1575" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0112_ = { wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1576" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0113_ = { wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1577" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0114_ = { img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1578" *) img2sbuf_p0_wr_addr[3:0];
  assign _0115_ = { img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1579" *) img2sbuf_p1_wr_addr[3:0];
  assign _0116_ = { dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1595" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0117_ = { dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1596" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0118_ = { wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1597" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0119_ = { wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1598" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0120_ = { img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1599" *) img2sbuf_p0_wr_addr[3:0];
  assign _0121_ = { img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1600" *) img2sbuf_p1_wr_addr[3:0];
  assign _0122_ = { dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1616" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0123_ = { dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1617" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0124_ = { wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1618" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0125_ = { wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1619" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0126_ = { img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1620" *) img2sbuf_p0_wr_addr[3:0];
  assign _0127_ = { img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1621" *) img2sbuf_p1_wr_addr[3:0];
  assign _0128_ = { dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1637" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0129_ = { dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1638" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0130_ = { wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1639" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0131_ = { wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1640" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0132_ = { img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1641" *) img2sbuf_p0_wr_addr[3:0];
  assign _0133_ = { img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1642" *) img2sbuf_p1_wr_addr[3:0];
  assign _0134_ = { dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1658" *) dc2sbuf_p0_wr_addr[3:0];
  assign _0135_ = { dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1659" *) dc2sbuf_p1_wr_addr[3:0];
  assign _0136_ = { wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1660" *) wg2sbuf_p0_wr_addr[3:0];
  assign _0137_ = { wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1661" *) wg2sbuf_p1_wr_addr[3:0];
  assign _0138_ = { img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1662" *) img2sbuf_p0_wr_addr[3:0];
  assign _0139_ = { img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1663" *) img2sbuf_p1_wr_addr[3:0];
  assign _0140_ = { dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00, dc2sbuf_p0_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1679" *) dc2sbuf_p0_wr_data;
  assign _0141_ = { dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00, dc2sbuf_p1_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1680" *) dc2sbuf_p1_wr_data;
  assign _0142_ = { wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00, wg2sbuf_p0_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1681" *) wg2sbuf_p0_wr_data;
  assign _0143_ = { wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00, wg2sbuf_p1_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1682" *) wg2sbuf_p1_wr_data;
  assign _0144_ = { img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00, img2sbuf_p0_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1683" *) img2sbuf_p0_wr_data;
  assign _0145_ = { img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00, img2sbuf_p1_wr_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1684" *) img2sbuf_p1_wr_data;
  assign _0146_ = { dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01, dc2sbuf_p0_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1700" *) dc2sbuf_p0_wr_data;
  assign _0147_ = { dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01, dc2sbuf_p1_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1701" *) dc2sbuf_p1_wr_data;
  assign _0148_ = { wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01, wg2sbuf_p0_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1702" *) wg2sbuf_p0_wr_data;
  assign _0149_ = { wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01, wg2sbuf_p1_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1703" *) wg2sbuf_p1_wr_data;
  assign _0150_ = { img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01, img2sbuf_p0_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1704" *) img2sbuf_p0_wr_data;
  assign _0151_ = { img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01, img2sbuf_p1_wr_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1705" *) img2sbuf_p1_wr_data;
  assign _0152_ = { dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02, dc2sbuf_p0_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1721" *) dc2sbuf_p0_wr_data;
  assign _0153_ = { dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02, dc2sbuf_p1_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1722" *) dc2sbuf_p1_wr_data;
  assign _0154_ = { wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02, wg2sbuf_p0_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1723" *) wg2sbuf_p0_wr_data;
  assign _0155_ = { wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02, wg2sbuf_p1_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1724" *) wg2sbuf_p1_wr_data;
  assign _0156_ = { img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02, img2sbuf_p0_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1725" *) img2sbuf_p0_wr_data;
  assign _0157_ = { img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02, img2sbuf_p1_wr_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1726" *) img2sbuf_p1_wr_data;
  assign _0158_ = { dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03, dc2sbuf_p0_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1742" *) dc2sbuf_p0_wr_data;
  assign _0159_ = { dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03, dc2sbuf_p1_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1743" *) dc2sbuf_p1_wr_data;
  assign _0160_ = { wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03, wg2sbuf_p0_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1744" *) wg2sbuf_p0_wr_data;
  assign _0161_ = { wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03, wg2sbuf_p1_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1745" *) wg2sbuf_p1_wr_data;
  assign _0162_ = { img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03, img2sbuf_p0_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1746" *) img2sbuf_p0_wr_data;
  assign _0163_ = { img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03, img2sbuf_p1_wr_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1747" *) img2sbuf_p1_wr_data;
  assign _0164_ = { dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04, dc2sbuf_p0_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1763" *) dc2sbuf_p0_wr_data;
  assign _0165_ = { dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04, dc2sbuf_p1_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1764" *) dc2sbuf_p1_wr_data;
  assign _0166_ = { wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04, wg2sbuf_p0_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1765" *) wg2sbuf_p0_wr_data;
  assign _0167_ = { wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04, wg2sbuf_p1_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1766" *) wg2sbuf_p1_wr_data;
  assign _0168_ = { img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04, img2sbuf_p0_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1767" *) img2sbuf_p0_wr_data;
  assign _0169_ = { img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04, img2sbuf_p1_wr_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1768" *) img2sbuf_p1_wr_data;
  assign _0170_ = { dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05, dc2sbuf_p0_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1784" *) dc2sbuf_p0_wr_data;
  assign _0171_ = { dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05, dc2sbuf_p1_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1785" *) dc2sbuf_p1_wr_data;
  assign _0172_ = { wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05, wg2sbuf_p0_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1786" *) wg2sbuf_p0_wr_data;
  assign _0173_ = { wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05, wg2sbuf_p1_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1787" *) wg2sbuf_p1_wr_data;
  assign _0174_ = { img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05, img2sbuf_p0_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1788" *) img2sbuf_p0_wr_data;
  assign _0175_ = { img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05, img2sbuf_p1_wr_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1789" *) img2sbuf_p1_wr_data;
  assign _0176_ = { dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06, dc2sbuf_p0_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1805" *) dc2sbuf_p0_wr_data;
  assign _0177_ = { dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06, dc2sbuf_p1_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1806" *) dc2sbuf_p1_wr_data;
  assign _0178_ = { wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06, wg2sbuf_p0_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1807" *) wg2sbuf_p0_wr_data;
  assign _0179_ = { wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06, wg2sbuf_p1_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1808" *) wg2sbuf_p1_wr_data;
  assign _0180_ = { img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06, img2sbuf_p0_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1809" *) img2sbuf_p0_wr_data;
  assign _0181_ = { img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06, img2sbuf_p1_wr_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1810" *) img2sbuf_p1_wr_data;
  assign _0182_ = { dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07, dc2sbuf_p0_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1826" *) dc2sbuf_p0_wr_data;
  assign _0183_ = { dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07, dc2sbuf_p1_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1827" *) dc2sbuf_p1_wr_data;
  assign _0184_ = { wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07, wg2sbuf_p0_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1828" *) wg2sbuf_p0_wr_data;
  assign _0185_ = { wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07, wg2sbuf_p1_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1829" *) wg2sbuf_p1_wr_data;
  assign _0186_ = { img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07, img2sbuf_p0_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1830" *) img2sbuf_p0_wr_data;
  assign _0187_ = { img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07, img2sbuf_p1_wr_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1831" *) img2sbuf_p1_wr_data;
  assign _0188_ = { dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08, dc2sbuf_p0_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1847" *) dc2sbuf_p0_wr_data;
  assign _0189_ = { dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08, dc2sbuf_p1_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1848" *) dc2sbuf_p1_wr_data;
  assign _0190_ = { wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08, wg2sbuf_p0_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1849" *) wg2sbuf_p0_wr_data;
  assign _0191_ = { wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08, wg2sbuf_p1_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1850" *) wg2sbuf_p1_wr_data;
  assign _0192_ = { img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08, img2sbuf_p0_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1851" *) img2sbuf_p0_wr_data;
  assign _0193_ = { img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08, img2sbuf_p1_wr_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1852" *) img2sbuf_p1_wr_data;
  assign _0194_ = { dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09, dc2sbuf_p0_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1868" *) dc2sbuf_p0_wr_data;
  assign _0195_ = { dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09, dc2sbuf_p1_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1869" *) dc2sbuf_p1_wr_data;
  assign _0196_ = { wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09, wg2sbuf_p0_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1870" *) wg2sbuf_p0_wr_data;
  assign _0197_ = { wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09, wg2sbuf_p1_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1871" *) wg2sbuf_p1_wr_data;
  assign _0198_ = { img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09, img2sbuf_p0_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1872" *) img2sbuf_p0_wr_data;
  assign _0199_ = { img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09, img2sbuf_p1_wr_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1873" *) img2sbuf_p1_wr_data;
  assign _0200_ = { dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10, dc2sbuf_p0_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1889" *) dc2sbuf_p0_wr_data;
  assign _0201_ = { dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10, dc2sbuf_p1_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1890" *) dc2sbuf_p1_wr_data;
  assign _0202_ = { wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10, wg2sbuf_p0_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1891" *) wg2sbuf_p0_wr_data;
  assign _0203_ = { wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10, wg2sbuf_p1_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1892" *) wg2sbuf_p1_wr_data;
  assign _0204_ = { img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10, img2sbuf_p0_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1893" *) img2sbuf_p0_wr_data;
  assign _0205_ = { img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10, img2sbuf_p1_wr_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1894" *) img2sbuf_p1_wr_data;
  assign _0206_ = { dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11, dc2sbuf_p0_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1910" *) dc2sbuf_p0_wr_data;
  assign _0207_ = { dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11, dc2sbuf_p1_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1911" *) dc2sbuf_p1_wr_data;
  assign _0208_ = { wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11, wg2sbuf_p0_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1912" *) wg2sbuf_p0_wr_data;
  assign _0209_ = { wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11, wg2sbuf_p1_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1913" *) wg2sbuf_p1_wr_data;
  assign _0210_ = { img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11, img2sbuf_p0_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1914" *) img2sbuf_p0_wr_data;
  assign _0211_ = { img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11, img2sbuf_p1_wr_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1915" *) img2sbuf_p1_wr_data;
  assign _0212_ = { dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12, dc2sbuf_p0_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1931" *) dc2sbuf_p0_wr_data;
  assign _0213_ = { dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12, dc2sbuf_p1_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1932" *) dc2sbuf_p1_wr_data;
  assign _0214_ = { wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12, wg2sbuf_p0_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1933" *) wg2sbuf_p0_wr_data;
  assign _0215_ = { wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12, wg2sbuf_p1_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1934" *) wg2sbuf_p1_wr_data;
  assign _0216_ = { img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12, img2sbuf_p0_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1935" *) img2sbuf_p0_wr_data;
  assign _0217_ = { img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12, img2sbuf_p1_wr_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1936" *) img2sbuf_p1_wr_data;
  assign _0218_ = { dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13, dc2sbuf_p0_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1952" *) dc2sbuf_p0_wr_data;
  assign _0219_ = { dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13, dc2sbuf_p1_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1953" *) dc2sbuf_p1_wr_data;
  assign _0220_ = { wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13, wg2sbuf_p0_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1954" *) wg2sbuf_p0_wr_data;
  assign _0221_ = { wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13, wg2sbuf_p1_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1955" *) wg2sbuf_p1_wr_data;
  assign _0222_ = { img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13, img2sbuf_p0_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1956" *) img2sbuf_p0_wr_data;
  assign _0223_ = { img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13, img2sbuf_p1_wr_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1957" *) img2sbuf_p1_wr_data;
  assign _0224_ = { dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14, dc2sbuf_p0_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1973" *) dc2sbuf_p0_wr_data;
  assign _0225_ = { dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14, dc2sbuf_p1_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1974" *) dc2sbuf_p1_wr_data;
  assign _0226_ = { wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14, wg2sbuf_p0_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1975" *) wg2sbuf_p0_wr_data;
  assign _0227_ = { wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14, wg2sbuf_p1_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1976" *) wg2sbuf_p1_wr_data;
  assign _0228_ = { img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14, img2sbuf_p0_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1977" *) img2sbuf_p0_wr_data;
  assign _0229_ = { img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14, img2sbuf_p1_wr_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1978" *) img2sbuf_p1_wr_data;
  assign _0230_ = { dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15, dc2sbuf_p0_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1994" *) dc2sbuf_p0_wr_data;
  assign _0231_ = { dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15, dc2sbuf_p1_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1995" *) dc2sbuf_p1_wr_data;
  assign _0232_ = { wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15, wg2sbuf_p0_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1996" *) wg2sbuf_p0_wr_data;
  assign _0233_ = { wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15, wg2sbuf_p1_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1997" *) wg2sbuf_p1_wr_data;
  assign _0234_ = { img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15, img2sbuf_p0_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1998" *) img2sbuf_p0_wr_data;
  assign _0235_ = { img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15, img2sbuf_p1_wr_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1999" *) img2sbuf_p1_wr_data;
  assign dc2sbuf_p0_rd_sel_00 = _0395_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2177" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_00 = _0396_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2183" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_00 = _0397_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2189" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_00 = _0398_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2195" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_01 = _0399_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2201" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_01 = _0400_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2207" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_01 = _0401_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2213" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_01 = _0402_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2219" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_02 = _0403_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2225" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_02 = _0404_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2231" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_02 = _0405_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2237" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_02 = _0406_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2243" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_03 = _0407_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2249" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_03 = _0408_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2255" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_03 = _0409_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2261" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_03 = _0410_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2267" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_04 = _0411_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2273" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_04 = _0412_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2279" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_04 = _0413_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2285" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_04 = _0414_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2291" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_05 = _0415_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2297" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_05 = _0416_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2303" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_05 = _0417_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2309" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_05 = _0418_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2315" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_06 = _0419_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2321" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_06 = _0420_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2327" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_06 = _0421_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2333" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_06 = _0422_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2339" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_07 = _0423_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2345" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_07 = _0424_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2351" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_07 = _0425_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2357" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_07 = _0426_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2363" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_08 = _0427_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2369" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_08 = _0428_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2375" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_08 = _0429_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2381" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_08 = _0430_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2387" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_09 = _0431_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2393" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_09 = _0432_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2399" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_09 = _0433_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2405" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_09 = _0434_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2411" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_10 = _0435_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2417" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_10 = _0436_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2423" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_10 = _0437_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2429" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_10 = _0438_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2435" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_11 = _0439_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2441" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_11 = _0440_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2447" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_11 = _0441_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2453" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_11 = _0442_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2459" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_12 = _0443_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2465" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_12 = _0444_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2471" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_12 = _0445_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2477" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_12 = _0446_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2483" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_13 = _0447_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2489" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_13 = _0448_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2495" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_13 = _0449_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2501" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_13 = _0450_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2507" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_14 = _0451_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2513" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_14 = _0452_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2519" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_14 = _0453_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2525" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_14 = _0454_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2531" *) img2sbuf_p1_rd_en;
  assign dc2sbuf_p0_rd_sel_15 = _0455_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2537" *) dc2sbuf_p0_rd_en;
  assign dc2sbuf_p1_rd_sel_15 = _0456_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2543" *) dc2sbuf_p1_rd_en;
  assign img2sbuf_p0_rd_sel_15 = _0457_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2549" *) img2sbuf_p0_rd_en;
  assign img2sbuf_p1_rd_sel_15 = _0458_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2555" *) img2sbuf_p1_rd_en;
  assign wg2sbuf_p0_rd_sel_00 = _0459_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2561" *) wg2sbuf_p0_rd_en;
  assign wg2sbuf_p1_rd_sel_00 = _0460_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2567" *) wg2sbuf_p1_rd_en;
  assign wg2sbuf_p0_rd_sel_04 = _0461_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2609" *) wg2sbuf_p0_rd_en;
  assign wg2sbuf_p1_rd_sel_04 = _0462_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2615" *) wg2sbuf_p1_rd_en;
  assign wg2sbuf_p0_rd_sel_08 = _0463_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2657" *) wg2sbuf_p0_rd_en;
  assign wg2sbuf_p1_rd_sel_08 = _0464_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2663" *) wg2sbuf_p1_rd_en;
  assign wg2sbuf_p0_rd_sel_12 = _0465_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2705" *) wg2sbuf_p0_rd_en;
  assign wg2sbuf_p1_rd_sel_12 = _0466_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2711" *) wg2sbuf_p1_rd_en;
  assign _0236_ = { dc2sbuf_p0_rd_sel_00, dc2sbuf_p0_rd_sel_00, dc2sbuf_p0_rd_sel_00, dc2sbuf_p0_rd_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3089" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0237_ = { dc2sbuf_p1_rd_sel_00, dc2sbuf_p1_rd_sel_00, dc2sbuf_p1_rd_sel_00, dc2sbuf_p1_rd_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3090" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0238_ = { wg2sbuf_p0_rd_sel_00, wg2sbuf_p0_rd_sel_00, wg2sbuf_p0_rd_sel_00, wg2sbuf_p0_rd_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3091" *) wg2sbuf_p0_rd_addr[5:2];
  assign _0239_ = { wg2sbuf_p1_rd_sel_00, wg2sbuf_p1_rd_sel_00, wg2sbuf_p1_rd_sel_00, wg2sbuf_p1_rd_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3092" *) wg2sbuf_p1_rd_addr[5:2];
  assign _0240_ = { img2sbuf_p0_rd_sel_00, img2sbuf_p0_rd_sel_00, img2sbuf_p0_rd_sel_00, img2sbuf_p0_rd_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3093" *) img2sbuf_p0_rd_addr[3:0];
  assign _0241_ = { img2sbuf_p1_rd_sel_00, img2sbuf_p1_rd_sel_00, img2sbuf_p1_rd_sel_00, img2sbuf_p1_rd_sel_00 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3094" *) img2sbuf_p1_rd_addr[3:0];
  assign _0242_ = { dc2sbuf_p0_rd_sel_01, dc2sbuf_p0_rd_sel_01, dc2sbuf_p0_rd_sel_01, dc2sbuf_p0_rd_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3110" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0243_ = { dc2sbuf_p1_rd_sel_01, dc2sbuf_p1_rd_sel_01, dc2sbuf_p1_rd_sel_01, dc2sbuf_p1_rd_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3111" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0244_ = { img2sbuf_p0_rd_sel_01, img2sbuf_p0_rd_sel_01, img2sbuf_p0_rd_sel_01, img2sbuf_p0_rd_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3114" *) img2sbuf_p0_rd_addr[3:0];
  assign _0245_ = { img2sbuf_p1_rd_sel_01, img2sbuf_p1_rd_sel_01, img2sbuf_p1_rd_sel_01, img2sbuf_p1_rd_sel_01 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3115" *) img2sbuf_p1_rd_addr[3:0];
  assign _0246_ = { dc2sbuf_p0_rd_sel_02, dc2sbuf_p0_rd_sel_02, dc2sbuf_p0_rd_sel_02, dc2sbuf_p0_rd_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3131" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0247_ = { dc2sbuf_p1_rd_sel_02, dc2sbuf_p1_rd_sel_02, dc2sbuf_p1_rd_sel_02, dc2sbuf_p1_rd_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3132" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0248_ = { img2sbuf_p0_rd_sel_02, img2sbuf_p0_rd_sel_02, img2sbuf_p0_rd_sel_02, img2sbuf_p0_rd_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3135" *) img2sbuf_p0_rd_addr[3:0];
  assign _0249_ = { img2sbuf_p1_rd_sel_02, img2sbuf_p1_rd_sel_02, img2sbuf_p1_rd_sel_02, img2sbuf_p1_rd_sel_02 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3136" *) img2sbuf_p1_rd_addr[3:0];
  assign _0250_ = { dc2sbuf_p0_rd_sel_03, dc2sbuf_p0_rd_sel_03, dc2sbuf_p0_rd_sel_03, dc2sbuf_p0_rd_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3152" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0251_ = { dc2sbuf_p1_rd_sel_03, dc2sbuf_p1_rd_sel_03, dc2sbuf_p1_rd_sel_03, dc2sbuf_p1_rd_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3153" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0252_ = { img2sbuf_p0_rd_sel_03, img2sbuf_p0_rd_sel_03, img2sbuf_p0_rd_sel_03, img2sbuf_p0_rd_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3156" *) img2sbuf_p0_rd_addr[3:0];
  assign _0253_ = { img2sbuf_p1_rd_sel_03, img2sbuf_p1_rd_sel_03, img2sbuf_p1_rd_sel_03, img2sbuf_p1_rd_sel_03 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3157" *) img2sbuf_p1_rd_addr[3:0];
  assign _0254_ = { dc2sbuf_p0_rd_sel_04, dc2sbuf_p0_rd_sel_04, dc2sbuf_p0_rd_sel_04, dc2sbuf_p0_rd_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3173" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0255_ = { dc2sbuf_p1_rd_sel_04, dc2sbuf_p1_rd_sel_04, dc2sbuf_p1_rd_sel_04, dc2sbuf_p1_rd_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3174" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0256_ = { wg2sbuf_p0_rd_sel_04, wg2sbuf_p0_rd_sel_04, wg2sbuf_p0_rd_sel_04, wg2sbuf_p0_rd_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3175" *) wg2sbuf_p0_rd_addr[5:2];
  assign _0257_ = { wg2sbuf_p1_rd_sel_04, wg2sbuf_p1_rd_sel_04, wg2sbuf_p1_rd_sel_04, wg2sbuf_p1_rd_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3176" *) wg2sbuf_p1_rd_addr[5:2];
  assign _0258_ = { img2sbuf_p0_rd_sel_04, img2sbuf_p0_rd_sel_04, img2sbuf_p0_rd_sel_04, img2sbuf_p0_rd_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3177" *) img2sbuf_p0_rd_addr[3:0];
  assign _0259_ = { img2sbuf_p1_rd_sel_04, img2sbuf_p1_rd_sel_04, img2sbuf_p1_rd_sel_04, img2sbuf_p1_rd_sel_04 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3178" *) img2sbuf_p1_rd_addr[3:0];
  assign _0260_ = { dc2sbuf_p0_rd_sel_05, dc2sbuf_p0_rd_sel_05, dc2sbuf_p0_rd_sel_05, dc2sbuf_p0_rd_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3194" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0261_ = { dc2sbuf_p1_rd_sel_05, dc2sbuf_p1_rd_sel_05, dc2sbuf_p1_rd_sel_05, dc2sbuf_p1_rd_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3195" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0262_ = { img2sbuf_p0_rd_sel_05, img2sbuf_p0_rd_sel_05, img2sbuf_p0_rd_sel_05, img2sbuf_p0_rd_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3198" *) img2sbuf_p0_rd_addr[3:0];
  assign _0263_ = { img2sbuf_p1_rd_sel_05, img2sbuf_p1_rd_sel_05, img2sbuf_p1_rd_sel_05, img2sbuf_p1_rd_sel_05 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3199" *) img2sbuf_p1_rd_addr[3:0];
  assign _0264_ = { dc2sbuf_p0_rd_sel_06, dc2sbuf_p0_rd_sel_06, dc2sbuf_p0_rd_sel_06, dc2sbuf_p0_rd_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3215" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0265_ = { dc2sbuf_p1_rd_sel_06, dc2sbuf_p1_rd_sel_06, dc2sbuf_p1_rd_sel_06, dc2sbuf_p1_rd_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3216" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0266_ = { img2sbuf_p0_rd_sel_06, img2sbuf_p0_rd_sel_06, img2sbuf_p0_rd_sel_06, img2sbuf_p0_rd_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3219" *) img2sbuf_p0_rd_addr[3:0];
  assign _0267_ = { img2sbuf_p1_rd_sel_06, img2sbuf_p1_rd_sel_06, img2sbuf_p1_rd_sel_06, img2sbuf_p1_rd_sel_06 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3220" *) img2sbuf_p1_rd_addr[3:0];
  assign _0268_ = { dc2sbuf_p0_rd_sel_07, dc2sbuf_p0_rd_sel_07, dc2sbuf_p0_rd_sel_07, dc2sbuf_p0_rd_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3236" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0269_ = { dc2sbuf_p1_rd_sel_07, dc2sbuf_p1_rd_sel_07, dc2sbuf_p1_rd_sel_07, dc2sbuf_p1_rd_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3237" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0270_ = { img2sbuf_p0_rd_sel_07, img2sbuf_p0_rd_sel_07, img2sbuf_p0_rd_sel_07, img2sbuf_p0_rd_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3240" *) img2sbuf_p0_rd_addr[3:0];
  assign _0271_ = { img2sbuf_p1_rd_sel_07, img2sbuf_p1_rd_sel_07, img2sbuf_p1_rd_sel_07, img2sbuf_p1_rd_sel_07 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3241" *) img2sbuf_p1_rd_addr[3:0];
  assign _0272_ = { dc2sbuf_p0_rd_sel_08, dc2sbuf_p0_rd_sel_08, dc2sbuf_p0_rd_sel_08, dc2sbuf_p0_rd_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3257" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0273_ = { dc2sbuf_p1_rd_sel_08, dc2sbuf_p1_rd_sel_08, dc2sbuf_p1_rd_sel_08, dc2sbuf_p1_rd_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3258" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0274_ = { wg2sbuf_p0_rd_sel_08, wg2sbuf_p0_rd_sel_08, wg2sbuf_p0_rd_sel_08, wg2sbuf_p0_rd_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3259" *) wg2sbuf_p0_rd_addr[5:2];
  assign _0275_ = { wg2sbuf_p1_rd_sel_08, wg2sbuf_p1_rd_sel_08, wg2sbuf_p1_rd_sel_08, wg2sbuf_p1_rd_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3260" *) wg2sbuf_p1_rd_addr[5:2];
  assign _0276_ = { img2sbuf_p0_rd_sel_08, img2sbuf_p0_rd_sel_08, img2sbuf_p0_rd_sel_08, img2sbuf_p0_rd_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3261" *) img2sbuf_p0_rd_addr[3:0];
  assign _0277_ = { img2sbuf_p1_rd_sel_08, img2sbuf_p1_rd_sel_08, img2sbuf_p1_rd_sel_08, img2sbuf_p1_rd_sel_08 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3262" *) img2sbuf_p1_rd_addr[3:0];
  assign _0278_ = { dc2sbuf_p0_rd_sel_09, dc2sbuf_p0_rd_sel_09, dc2sbuf_p0_rd_sel_09, dc2sbuf_p0_rd_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3278" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0279_ = { dc2sbuf_p1_rd_sel_09, dc2sbuf_p1_rd_sel_09, dc2sbuf_p1_rd_sel_09, dc2sbuf_p1_rd_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3279" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0280_ = { img2sbuf_p0_rd_sel_09, img2sbuf_p0_rd_sel_09, img2sbuf_p0_rd_sel_09, img2sbuf_p0_rd_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3282" *) img2sbuf_p0_rd_addr[3:0];
  assign _0281_ = { img2sbuf_p1_rd_sel_09, img2sbuf_p1_rd_sel_09, img2sbuf_p1_rd_sel_09, img2sbuf_p1_rd_sel_09 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3283" *) img2sbuf_p1_rd_addr[3:0];
  assign _0282_ = { dc2sbuf_p0_rd_sel_10, dc2sbuf_p0_rd_sel_10, dc2sbuf_p0_rd_sel_10, dc2sbuf_p0_rd_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3299" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0283_ = { dc2sbuf_p1_rd_sel_10, dc2sbuf_p1_rd_sel_10, dc2sbuf_p1_rd_sel_10, dc2sbuf_p1_rd_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3300" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0284_ = { img2sbuf_p0_rd_sel_10, img2sbuf_p0_rd_sel_10, img2sbuf_p0_rd_sel_10, img2sbuf_p0_rd_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3303" *) img2sbuf_p0_rd_addr[3:0];
  assign _0285_ = { img2sbuf_p1_rd_sel_10, img2sbuf_p1_rd_sel_10, img2sbuf_p1_rd_sel_10, img2sbuf_p1_rd_sel_10 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3304" *) img2sbuf_p1_rd_addr[3:0];
  assign _0286_ = { dc2sbuf_p0_rd_sel_11, dc2sbuf_p0_rd_sel_11, dc2sbuf_p0_rd_sel_11, dc2sbuf_p0_rd_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3320" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0287_ = { dc2sbuf_p1_rd_sel_11, dc2sbuf_p1_rd_sel_11, dc2sbuf_p1_rd_sel_11, dc2sbuf_p1_rd_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3321" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0288_ = { img2sbuf_p0_rd_sel_11, img2sbuf_p0_rd_sel_11, img2sbuf_p0_rd_sel_11, img2sbuf_p0_rd_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3324" *) img2sbuf_p0_rd_addr[3:0];
  assign _0289_ = { img2sbuf_p1_rd_sel_11, img2sbuf_p1_rd_sel_11, img2sbuf_p1_rd_sel_11, img2sbuf_p1_rd_sel_11 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3325" *) img2sbuf_p1_rd_addr[3:0];
  assign _0290_ = { dc2sbuf_p0_rd_sel_12, dc2sbuf_p0_rd_sel_12, dc2sbuf_p0_rd_sel_12, dc2sbuf_p0_rd_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3341" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0291_ = { dc2sbuf_p1_rd_sel_12, dc2sbuf_p1_rd_sel_12, dc2sbuf_p1_rd_sel_12, dc2sbuf_p1_rd_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3342" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0292_ = { wg2sbuf_p0_rd_sel_12, wg2sbuf_p0_rd_sel_12, wg2sbuf_p0_rd_sel_12, wg2sbuf_p0_rd_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3343" *) wg2sbuf_p0_rd_addr[5:2];
  assign _0293_ = { wg2sbuf_p1_rd_sel_12, wg2sbuf_p1_rd_sel_12, wg2sbuf_p1_rd_sel_12, wg2sbuf_p1_rd_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3344" *) wg2sbuf_p1_rd_addr[5:2];
  assign _0294_ = { img2sbuf_p0_rd_sel_12, img2sbuf_p0_rd_sel_12, img2sbuf_p0_rd_sel_12, img2sbuf_p0_rd_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3345" *) img2sbuf_p0_rd_addr[3:0];
  assign _0295_ = { img2sbuf_p1_rd_sel_12, img2sbuf_p1_rd_sel_12, img2sbuf_p1_rd_sel_12, img2sbuf_p1_rd_sel_12 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3346" *) img2sbuf_p1_rd_addr[3:0];
  assign _0296_ = { dc2sbuf_p0_rd_sel_13, dc2sbuf_p0_rd_sel_13, dc2sbuf_p0_rd_sel_13, dc2sbuf_p0_rd_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3362" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0297_ = { dc2sbuf_p1_rd_sel_13, dc2sbuf_p1_rd_sel_13, dc2sbuf_p1_rd_sel_13, dc2sbuf_p1_rd_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3363" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0298_ = { img2sbuf_p0_rd_sel_13, img2sbuf_p0_rd_sel_13, img2sbuf_p0_rd_sel_13, img2sbuf_p0_rd_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3366" *) img2sbuf_p0_rd_addr[3:0];
  assign _0299_ = { img2sbuf_p1_rd_sel_13, img2sbuf_p1_rd_sel_13, img2sbuf_p1_rd_sel_13, img2sbuf_p1_rd_sel_13 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3367" *) img2sbuf_p1_rd_addr[3:0];
  assign _0300_ = { dc2sbuf_p0_rd_sel_14, dc2sbuf_p0_rd_sel_14, dc2sbuf_p0_rd_sel_14, dc2sbuf_p0_rd_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3383" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0301_ = { dc2sbuf_p1_rd_sel_14, dc2sbuf_p1_rd_sel_14, dc2sbuf_p1_rd_sel_14, dc2sbuf_p1_rd_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3384" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0302_ = { img2sbuf_p0_rd_sel_14, img2sbuf_p0_rd_sel_14, img2sbuf_p0_rd_sel_14, img2sbuf_p0_rd_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3387" *) img2sbuf_p0_rd_addr[3:0];
  assign _0303_ = { img2sbuf_p1_rd_sel_14, img2sbuf_p1_rd_sel_14, img2sbuf_p1_rd_sel_14, img2sbuf_p1_rd_sel_14 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3388" *) img2sbuf_p1_rd_addr[3:0];
  assign _0304_ = { dc2sbuf_p0_rd_sel_15, dc2sbuf_p0_rd_sel_15, dc2sbuf_p0_rd_sel_15, dc2sbuf_p0_rd_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3404" *) dc2sbuf_p0_rd_addr[3:0];
  assign _0305_ = { dc2sbuf_p1_rd_sel_15, dc2sbuf_p1_rd_sel_15, dc2sbuf_p1_rd_sel_15, dc2sbuf_p1_rd_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3405" *) dc2sbuf_p1_rd_addr[3:0];
  assign _0306_ = { img2sbuf_p0_rd_sel_15, img2sbuf_p0_rd_sel_15, img2sbuf_p0_rd_sel_15, img2sbuf_p0_rd_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3408" *) img2sbuf_p0_rd_addr[3:0];
  assign _0307_ = { img2sbuf_p1_rd_sel_15, img2sbuf_p1_rd_sel_15, img2sbuf_p1_rd_sel_15, img2sbuf_p1_rd_sel_15 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3409" *) img2sbuf_p1_rd_addr[3:0];
  assign sbuf_p0_wg_sel_q0 = _0467_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3415" *) wg2sbuf_p0_rd_en;
  assign sbuf_p0_wg_sel_q1 = _0468_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3421" *) wg2sbuf_p0_rd_en;
  assign sbuf_p0_wg_sel_q2 = _0469_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3427" *) wg2sbuf_p0_rd_en;
  assign sbuf_p0_wg_sel_q3 = _0470_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3433" *) wg2sbuf_p0_rd_en;
  assign sbuf_p1_wg_sel_q0 = _0471_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3439" *) wg2sbuf_p1_rd_en;
  assign sbuf_p1_wg_sel_q1 = _0472_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3445" *) wg2sbuf_p1_rd_en;
  assign sbuf_p1_wg_sel_q2 = _0473_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3451" *) wg2sbuf_p1_rd_en;
  assign sbuf_p1_wg_sel_q3 = _0474_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3457" *) wg2sbuf_p1_rd_en;
  assign _0002_ = sbuf_p0_re_00 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3466" *) _0556_;
  assign _0024_ = sbuf_p1_re_00 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3473" *) _0557_;
  assign _0004_ = sbuf_p0_re_01 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3480" *) _0556_;
  assign _0026_ = sbuf_p1_re_01 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3487" *) _0557_;
  assign _0006_ = sbuf_p0_re_02 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3494" *) _0556_;
  assign _0028_ = sbuf_p1_re_02 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3501" *) _0557_;
  assign _0008_ = sbuf_p0_re_03 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3508" *) _0556_;
  assign _0030_ = sbuf_p1_re_03 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3515" *) _0557_;
  assign _0010_ = sbuf_p0_re_04 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3522" *) _0556_;
  assign _0032_ = sbuf_p1_re_04 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3529" *) _0557_;
  assign _0011_ = sbuf_p0_re_05 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3536" *) _0556_;
  assign _0033_ = sbuf_p1_re_05 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3543" *) _0557_;
  assign _0012_ = sbuf_p0_re_06 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3550" *) _0556_;
  assign _0034_ = sbuf_p1_re_06 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3557" *) _0557_;
  assign _0013_ = sbuf_p0_re_07 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3564" *) _0556_;
  assign _0035_ = sbuf_p1_re_07 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3571" *) _0557_;
  assign _0014_ = sbuf_p0_re_08 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3578" *) _0556_;
  assign _0036_ = sbuf_p1_re_08 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3585" *) _0557_;
  assign _0015_ = sbuf_p0_re_09 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3592" *) _0556_;
  assign _0037_ = sbuf_p1_re_09 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3599" *) _0557_;
  assign _0016_ = sbuf_p0_re_10 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3606" *) _0556_;
  assign _0038_ = sbuf_p1_re_10 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3613" *) _0557_;
  assign _0017_ = sbuf_p0_re_11 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3620" *) _0556_;
  assign _0039_ = sbuf_p1_re_11 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3627" *) _0557_;
  assign _0018_ = sbuf_p0_re_12 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3634" *) _0556_;
  assign _0040_ = sbuf_p1_re_12 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3641" *) _0557_;
  assign _0019_ = sbuf_p0_re_13 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3648" *) _0556_;
  assign _0041_ = sbuf_p1_re_13 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3655" *) _0557_;
  assign _0020_ = sbuf_p0_re_14 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3662" *) _0556_;
  assign _0042_ = sbuf_p1_re_14 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3669" *) _0557_;
  assign _0021_ = sbuf_p0_re_15 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3676" *) _0556_;
  assign _0043_ = sbuf_p1_re_15 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3683" *) _0557_;
  assign _0003_ = sbuf_p0_re_00 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3690" *) wg2sbuf_p0_rd_en;
  assign _0025_ = sbuf_p1_re_00 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3697" *) wg2sbuf_p1_rd_en;
  assign _0005_ = sbuf_p0_re_04 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3704" *) wg2sbuf_p0_rd_en;
  assign _0027_ = sbuf_p1_re_04 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3711" *) wg2sbuf_p1_rd_en;
  assign _0007_ = sbuf_p0_re_08 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3718" *) wg2sbuf_p0_rd_en;
  assign _0029_ = sbuf_p1_re_08 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3725" *) wg2sbuf_p1_rd_en;
  assign _0009_ = sbuf_p0_re_12 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3732" *) wg2sbuf_p0_rd_en;
  assign _0031_ = sbuf_p1_re_12 & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3739" *) wg2sbuf_p1_rd_en;
  assign _0308_ = { sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1, sbuf_p0_re_00_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3849" *) sbuf_rdat_00;
  assign _0309_ = { sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1, sbuf_p0_re_01_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3850" *) sbuf_rdat_01;
  assign _0310_ = { sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1, sbuf_p0_re_02_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3851" *) sbuf_rdat_02;
  assign _0311_ = { sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1, sbuf_p0_re_03_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3852" *) sbuf_rdat_03;
  assign _0312_ = { sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1, sbuf_p0_re_04_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3853" *) sbuf_rdat_04;
  assign _0313_ = { sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1, sbuf_p0_re_05_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3854" *) sbuf_rdat_05;
  assign _0314_ = { sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1, sbuf_p0_re_06_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3855" *) sbuf_rdat_06;
  assign _0315_ = { sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1, sbuf_p0_re_07_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3856" *) sbuf_rdat_07;
  assign _0316_ = { sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1, sbuf_p0_re_08_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3857" *) sbuf_rdat_08;
  assign _0317_ = { sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1, sbuf_p0_re_09_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3858" *) sbuf_rdat_09;
  assign _0318_ = { sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1, sbuf_p0_re_10_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3859" *) sbuf_rdat_10;
  assign _0319_ = { sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1, sbuf_p0_re_11_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3860" *) sbuf_rdat_11;
  assign _0320_ = { sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1, sbuf_p0_re_12_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3861" *) sbuf_rdat_12;
  assign _0321_ = { sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1, sbuf_p0_re_13_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3862" *) sbuf_rdat_13;
  assign _0322_ = { sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1, sbuf_p0_re_14_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3863" *) sbuf_rdat_14;
  assign _0323_ = { sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1, sbuf_p0_re_15_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3864" *) sbuf_rdat_15;
  assign _0324_ = { sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1, sbuf_p1_re_00_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3900" *) sbuf_rdat_00;
  assign _0325_ = { sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1, sbuf_p1_re_01_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3901" *) sbuf_rdat_01;
  assign _0326_ = { sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1, sbuf_p1_re_02_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3902" *) sbuf_rdat_02;
  assign _0327_ = { sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1, sbuf_p1_re_03_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3903" *) sbuf_rdat_03;
  assign _0328_ = { sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1, sbuf_p1_re_04_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3904" *) sbuf_rdat_04;
  assign _0329_ = { sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1, sbuf_p1_re_05_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3905" *) sbuf_rdat_05;
  assign _0330_ = { sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1, sbuf_p1_re_06_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3906" *) sbuf_rdat_06;
  assign _0331_ = { sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1, sbuf_p1_re_07_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3907" *) sbuf_rdat_07;
  assign _0332_ = { sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1, sbuf_p1_re_08_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3908" *) sbuf_rdat_08;
  assign _0333_ = { sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1, sbuf_p1_re_09_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3909" *) sbuf_rdat_09;
  assign _0334_ = { sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1, sbuf_p1_re_10_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3910" *) sbuf_rdat_10;
  assign _0335_ = { sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1, sbuf_p1_re_11_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3911" *) sbuf_rdat_11;
  assign _0336_ = { sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1, sbuf_p1_re_12_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3912" *) sbuf_rdat_12;
  assign _0337_ = { sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1, sbuf_p1_re_13_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3913" *) sbuf_rdat_13;
  assign _0338_ = { sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1, sbuf_p1_re_14_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3914" *) sbuf_rdat_14;
  assign _0339_ = { sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1, sbuf_p1_re_15_norm_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3915" *) sbuf_rdat_15;
  assign _0340_ = { sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3927" *) sbuf_rdat_00;
  assign _0341_ = { sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3928" *) sbuf_rdat_04;
  assign _0342_ = { sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3929" *) sbuf_rdat_08;
  assign _0343_ = { sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3930" *) sbuf_rdat_12;
  assign _0344_ = { sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3942" *) sbuf_rdat_01;
  assign _0345_ = { sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3943" *) sbuf_rdat_05;
  assign _0346_ = { sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3944" *) sbuf_rdat_09;
  assign _0347_ = { sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3945" *) sbuf_rdat_13;
  assign _0348_ = { sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3957" *) sbuf_rdat_02;
  assign _0349_ = { sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3958" *) sbuf_rdat_06;
  assign _0350_ = { sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3959" *) sbuf_rdat_10;
  assign _0351_ = { sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3960" *) sbuf_rdat_14;
  assign _0352_ = { sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1, sbuf_p0_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3972" *) sbuf_rdat_03;
  assign _0353_ = { sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1, sbuf_p0_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3973" *) sbuf_rdat_07;
  assign _0354_ = { sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1, sbuf_p0_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3974" *) sbuf_rdat_11;
  assign _0355_ = { sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1, sbuf_p0_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3975" *) sbuf_rdat_15;
  assign _0356_ = { sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3987" *) sbuf_rdat_00;
  assign _0357_ = { sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3988" *) sbuf_rdat_04;
  assign _0358_ = { sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3989" *) sbuf_rdat_08;
  assign _0359_ = { sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3990" *) sbuf_rdat_12;
  assign _0360_ = { sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4002" *) sbuf_rdat_01;
  assign _0361_ = { sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4003" *) sbuf_rdat_05;
  assign _0362_ = { sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4004" *) sbuf_rdat_09;
  assign _0363_ = { sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4005" *) sbuf_rdat_13;
  assign _0364_ = { sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4017" *) sbuf_rdat_02;
  assign _0365_ = { sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4018" *) sbuf_rdat_06;
  assign _0366_ = { sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4019" *) sbuf_rdat_10;
  assign _0367_ = { sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4020" *) sbuf_rdat_14;
  assign _0368_ = { sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1, sbuf_p1_re_00_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4032" *) sbuf_rdat_03;
  assign _0369_ = { sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1, sbuf_p1_re_01_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4033" *) sbuf_rdat_07;
  assign _0370_ = { sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1, sbuf_p1_re_02_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4034" *) sbuf_rdat_11;
  assign _0371_ = { sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1, sbuf_p1_re_03_wg_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4035" *) sbuf_rdat_15;
  assign _0372_ = { sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1, sbuf_p0_wg_sel_q0_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4047" *) { sbuf_p0_wg_rdat_src_3[63:0], sbuf_p0_wg_rdat_src_2[63:0], sbuf_p0_wg_rdat_src_1[63:0], sbuf_p0_wg_rdat_src_0[63:0] };
  assign _0373_ = { sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1, sbuf_p0_wg_sel_q1_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4048" *) { sbuf_p0_wg_rdat_src_3[127:64], sbuf_p0_wg_rdat_src_2[127:64], sbuf_p0_wg_rdat_src_1[127:64], sbuf_p0_wg_rdat_src_0[127:64] };
  assign _0374_ = { sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1, sbuf_p0_wg_sel_q2_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4049" *) { sbuf_p0_wg_rdat_src_3[191:128], sbuf_p0_wg_rdat_src_2[191:128], sbuf_p0_wg_rdat_src_1[191:128], sbuf_p0_wg_rdat_src_0[191:128] };
  assign _0375_ = { sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1, sbuf_p0_wg_sel_q3_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4050" *) { sbuf_p0_wg_rdat_src_3[255:192], sbuf_p0_wg_rdat_src_2[255:192], sbuf_p0_wg_rdat_src_1[255:192], sbuf_p0_wg_rdat_src_0[255:192] };
  assign _0376_ = { sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1, sbuf_p1_wg_sel_q0_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4062" *) { sbuf_p1_wg_rdat_src_3[63:0], sbuf_p1_wg_rdat_src_2[63:0], sbuf_p1_wg_rdat_src_1[63:0], sbuf_p1_wg_rdat_src_0[63:0] };
  assign _0377_ = { sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1, sbuf_p1_wg_sel_q1_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4063" *) { sbuf_p1_wg_rdat_src_3[127:64], sbuf_p1_wg_rdat_src_2[127:64], sbuf_p1_wg_rdat_src_1[127:64], sbuf_p1_wg_rdat_src_0[127:64] };
  assign _0378_ = { sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1, sbuf_p1_wg_sel_q2_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4064" *) { sbuf_p1_wg_rdat_src_3[191:128], sbuf_p1_wg_rdat_src_2[191:128], sbuf_p1_wg_rdat_src_1[191:128], sbuf_p1_wg_rdat_src_0[191:128] };
  assign _0379_ = { sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1, sbuf_p1_wg_sel_q3_d1 } & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4065" *) { sbuf_p1_wg_rdat_src_3[255:192], sbuf_p1_wg_rdat_src_2[255:192], sbuf_p1_wg_rdat_src_1[255:192], sbuf_p1_wg_rdat_src_0[255:192] };
  assign dc2sbuf_p0_wr_sel_00 = _0475_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:517" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_00 = _0476_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:523" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_00 = _0477_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:529" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_00 = _0478_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:535" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_00 = _0479_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:541" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_00 = _0480_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:547" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_01 = _0481_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:553" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_01 = _0482_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:559" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_01 = _0483_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:565" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_01 = _0484_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:571" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_01 = _0485_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:577" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_01 = _0486_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:583" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_02 = _0487_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:589" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_02 = _0488_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:595" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_02 = _0489_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:601" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_02 = _0490_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:607" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_02 = _0491_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:613" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_02 = _0492_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:619" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_03 = _0493_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:625" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_03 = _0494_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:631" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_03 = _0495_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:637" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_03 = _0496_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:643" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_03 = _0497_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:649" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_03 = _0498_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:655" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_04 = _0499_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:661" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_04 = _0500_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:667" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_04 = _0501_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:673" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_04 = _0502_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:679" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_04 = _0503_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:685" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_04 = _0504_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:691" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_05 = _0505_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:697" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_05 = _0506_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:703" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_05 = _0507_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:709" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_05 = _0508_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:715" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_05 = _0509_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:721" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_05 = _0510_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:727" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_06 = _0511_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:733" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_06 = _0512_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:739" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_06 = _0513_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:745" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_06 = _0514_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:751" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_06 = _0515_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:757" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_06 = _0516_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:763" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_07 = _0517_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:769" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_07 = _0518_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:775" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_07 = _0519_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:781" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_07 = _0520_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:787" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_07 = _0521_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:793" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_07 = _0522_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:799" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_08 = _0523_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:805" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_08 = _0524_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:811" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_08 = _0525_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:817" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_08 = _0526_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:823" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_08 = _0527_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:829" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_08 = _0528_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:835" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_09 = _0529_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:841" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_09 = _0530_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:847" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_09 = _0531_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:853" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_09 = _0532_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:859" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_09 = _0533_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:865" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_09 = _0534_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:871" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_10 = _0535_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:877" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_10 = _0536_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:883" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_10 = _0537_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:889" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_10 = _0538_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:895" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_10 = _0539_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:901" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_10 = _0540_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:907" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_11 = _0541_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:913" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_11 = _0542_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:919" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_11 = _0543_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:925" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_11 = _0544_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:931" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_11 = _0545_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:937" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_11 = _0546_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:943" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_12 = _0547_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:949" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_12 = _0548_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:955" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_12 = _0549_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:961" *) wg2sbuf_p0_wr_en;
  assign wg2sbuf_p1_wr_sel_12 = _0550_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:967" *) wg2sbuf_p1_wr_en;
  assign img2sbuf_p0_wr_sel_12 = _0551_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:973" *) img2sbuf_p0_wr_en;
  assign img2sbuf_p1_wr_sel_12 = _0552_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:979" *) img2sbuf_p1_wr_en;
  assign dc2sbuf_p0_wr_sel_13 = _0553_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:985" *) dc2sbuf_p0_wr_en;
  assign dc2sbuf_p1_wr_sel_13 = _0554_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:991" *) dc2sbuf_p1_wr_en;
  assign wg2sbuf_p0_wr_sel_13 = _0555_ & (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:997" *) wg2sbuf_p0_wr_en;
  assign _0380_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1003" *) 4'b1101;
  assign _0381_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1009" *) 4'b1101;
  assign _0382_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1015" *) 4'b1101;
  assign _0383_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1021" *) 4'b1110;
  assign _0384_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1027" *) 4'b1110;
  assign _0385_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1033" *) 4'b1110;
  assign _0386_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1039" *) 4'b1110;
  assign _0387_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1045" *) 4'b1110;
  assign _0388_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1051" *) 4'b1110;
  assign _0389_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1057" *) 4'b1111;
  assign _0390_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1063" *) 4'b1111;
  assign _0391_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1069" *) 4'b1111;
  assign _0392_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1075" *) 4'b1111;
  assign _0393_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1081" *) 4'b1111;
  assign _0394_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1087" *) 4'b1111;
  assign _0395_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2177" *) dc2sbuf_p0_rd_addr[7:4];
  assign _0396_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2183" *) dc2sbuf_p1_rd_addr[7:4];
  assign _0397_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2189" *) img2sbuf_p0_rd_addr[7:4];
  assign _0398_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2195" *) img2sbuf_p1_rd_addr[7:4];
  assign _0399_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2201" *) 1'b1;
  assign _0400_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2207" *) 1'b1;
  assign _0401_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2213" *) 1'b1;
  assign _0402_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2219" *) 1'b1;
  assign _0403_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2225" *) 2'b10;
  assign _0404_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2231" *) 2'b10;
  assign _0405_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2237" *) 2'b10;
  assign _0406_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2243" *) 2'b10;
  assign _0407_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2249" *) 2'b11;
  assign _0408_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2255" *) 2'b11;
  assign _0409_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2261" *) 2'b11;
  assign _0410_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2267" *) 2'b11;
  assign _0411_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2273" *) 3'b100;
  assign _0412_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2279" *) 3'b100;
  assign _0413_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2285" *) 3'b100;
  assign _0414_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2291" *) 3'b100;
  assign _0415_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2297" *) 3'b101;
  assign _0416_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2303" *) 3'b101;
  assign _0417_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2309" *) 3'b101;
  assign _0418_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2315" *) 3'b101;
  assign _0419_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2321" *) 3'b110;
  assign _0420_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2327" *) 3'b110;
  assign _0421_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2333" *) 3'b110;
  assign _0422_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2339" *) 3'b110;
  assign _0423_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2345" *) 3'b111;
  assign _0424_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2351" *) 3'b111;
  assign _0425_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2357" *) 3'b111;
  assign _0426_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2363" *) 3'b111;
  assign _0427_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2369" *) 4'b1000;
  assign _0428_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2375" *) 4'b1000;
  assign _0429_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2381" *) 4'b1000;
  assign _0430_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2387" *) 4'b1000;
  assign _0431_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2393" *) 4'b1001;
  assign _0432_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2399" *) 4'b1001;
  assign _0433_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2405" *) 4'b1001;
  assign _0434_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2411" *) 4'b1001;
  assign _0435_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2417" *) 4'b1010;
  assign _0436_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2423" *) 4'b1010;
  assign _0437_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2429" *) 4'b1010;
  assign _0438_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2435" *) 4'b1010;
  assign _0439_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2441" *) 4'b1011;
  assign _0440_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2447" *) 4'b1011;
  assign _0441_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2453" *) 4'b1011;
  assign _0442_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2459" *) 4'b1011;
  assign _0443_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2465" *) 4'b1100;
  assign _0444_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2471" *) 4'b1100;
  assign _0445_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2477" *) 4'b1100;
  assign _0446_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2483" *) 4'b1100;
  assign _0447_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2489" *) 4'b1101;
  assign _0448_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2495" *) 4'b1101;
  assign _0449_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2501" *) 4'b1101;
  assign _0450_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2507" *) 4'b1101;
  assign _0451_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2513" *) 4'b1110;
  assign _0452_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2519" *) 4'b1110;
  assign _0453_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2525" *) 4'b1110;
  assign _0454_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2531" *) 4'b1110;
  assign _0455_ = dc2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2537" *) 4'b1111;
  assign _0456_ = dc2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2543" *) 4'b1111;
  assign _0457_ = img2sbuf_p0_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2549" *) 4'b1111;
  assign _0458_ = img2sbuf_p1_rd_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2555" *) 4'b1111;
  assign _0459_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2561" *) wg2sbuf_p0_rd_addr[7:6];
  assign _0460_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2567" *) wg2sbuf_p1_rd_addr[7:6];
  assign _0461_ = wg2sbuf_p0_rd_addr[7:6] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2609" *) 1'b1;
  assign _0462_ = wg2sbuf_p1_rd_addr[7:6] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2615" *) 1'b1;
  assign _0463_ = wg2sbuf_p0_rd_addr[7:6] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2657" *) 2'b10;
  assign _0464_ = wg2sbuf_p1_rd_addr[7:6] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2663" *) 2'b10;
  assign _0465_ = wg2sbuf_p0_rd_addr[7:6] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2705" *) 2'b11;
  assign _0466_ = wg2sbuf_p1_rd_addr[7:6] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2711" *) 2'b11;
  assign _0467_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3415" *) wg2sbuf_p0_rd_addr[1:0];
  assign _0468_ = wg2sbuf_p0_rd_addr[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3421" *) 1'b1;
  assign _0469_ = wg2sbuf_p0_rd_addr[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3427" *) 2'b10;
  assign _0470_ = wg2sbuf_p0_rd_addr[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3433" *) 2'b11;
  assign _0471_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3439" *) wg2sbuf_p1_rd_addr[1:0];
  assign _0472_ = wg2sbuf_p1_rd_addr[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3445" *) 1'b1;
  assign _0473_ = wg2sbuf_p1_rd_addr[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3451" *) 2'b10;
  assign _0474_ = wg2sbuf_p1_rd_addr[1:0] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3457" *) 2'b11;
  assign _0475_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:517" *) dc2sbuf_p0_wr_addr[7:4];
  assign _0476_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:523" *) dc2sbuf_p1_wr_addr[7:4];
  assign _0477_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:529" *) wg2sbuf_p0_wr_addr[7:4];
  assign _0478_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:535" *) wg2sbuf_p1_wr_addr[7:4];
  assign _0479_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:541" *) img2sbuf_p0_wr_addr[7:4];
  assign _0480_ = ! (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:547" *) img2sbuf_p1_wr_addr[7:4];
  assign _0481_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:553" *) 1'b1;
  assign _0482_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:559" *) 1'b1;
  assign _0483_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:565" *) 1'b1;
  assign _0484_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:571" *) 1'b1;
  assign _0485_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:577" *) 1'b1;
  assign _0486_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:583" *) 1'b1;
  assign _0487_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:589" *) 2'b10;
  assign _0488_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:595" *) 2'b10;
  assign _0489_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:601" *) 2'b10;
  assign _0490_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:607" *) 2'b10;
  assign _0491_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:613" *) 2'b10;
  assign _0492_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:619" *) 2'b10;
  assign _0493_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:625" *) 2'b11;
  assign _0494_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:631" *) 2'b11;
  assign _0495_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:637" *) 2'b11;
  assign _0496_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:643" *) 2'b11;
  assign _0497_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:649" *) 2'b11;
  assign _0498_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:655" *) 2'b11;
  assign _0499_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:661" *) 3'b100;
  assign _0500_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:667" *) 3'b100;
  assign _0501_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:673" *) 3'b100;
  assign _0502_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:679" *) 3'b100;
  assign _0503_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:685" *) 3'b100;
  assign _0504_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:691" *) 3'b100;
  assign _0505_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:697" *) 3'b101;
  assign _0506_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:703" *) 3'b101;
  assign _0507_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:709" *) 3'b101;
  assign _0508_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:715" *) 3'b101;
  assign _0509_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:721" *) 3'b101;
  assign _0510_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:727" *) 3'b101;
  assign _0511_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:733" *) 3'b110;
  assign _0512_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:739" *) 3'b110;
  assign _0513_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:745" *) 3'b110;
  assign _0514_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:751" *) 3'b110;
  assign _0515_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:757" *) 3'b110;
  assign _0516_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:763" *) 3'b110;
  assign _0517_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:769" *) 3'b111;
  assign _0518_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:775" *) 3'b111;
  assign _0519_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:781" *) 3'b111;
  assign _0520_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:787" *) 3'b111;
  assign _0521_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:793" *) 3'b111;
  assign _0522_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:799" *) 3'b111;
  assign _0523_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:805" *) 4'b1000;
  assign _0524_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:811" *) 4'b1000;
  assign _0525_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:817" *) 4'b1000;
  assign _0526_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:823" *) 4'b1000;
  assign _0527_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:829" *) 4'b1000;
  assign _0528_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:835" *) 4'b1000;
  assign _0529_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:841" *) 4'b1001;
  assign _0530_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:847" *) 4'b1001;
  assign _0531_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:853" *) 4'b1001;
  assign _0532_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:859" *) 4'b1001;
  assign _0533_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:865" *) 4'b1001;
  assign _0534_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:871" *) 4'b1001;
  assign _0535_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:877" *) 4'b1010;
  assign _0536_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:883" *) 4'b1010;
  assign _0537_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:889" *) 4'b1010;
  assign _0538_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:895" *) 4'b1010;
  assign _0539_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:901" *) 4'b1010;
  assign _0540_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:907" *) 4'b1010;
  assign _0541_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:913" *) 4'b1011;
  assign _0542_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:919" *) 4'b1011;
  assign _0543_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:925" *) 4'b1011;
  assign _0544_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:931" *) 4'b1011;
  assign _0545_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:937" *) 4'b1011;
  assign _0546_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:943" *) 4'b1011;
  assign _0547_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:949" *) 4'b1100;
  assign _0548_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:955" *) 4'b1100;
  assign _0549_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:961" *) 4'b1100;
  assign _0550_ = wg2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:967" *) 4'b1100;
  assign _0551_ = img2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:973" *) 4'b1100;
  assign _0552_ = img2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:979" *) 4'b1100;
  assign _0553_ = dc2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:985" *) 4'b1101;
  assign _0554_ = dc2sbuf_p1_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:991" *) 4'b1101;
  assign _0555_ = wg2sbuf_p0_wr_addr[7:4] == (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:997" *) 4'b1101;
  assign _0556_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3466" *) wg2sbuf_p0_rd_en;
  assign _0557_ = ~ (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3473" *) wg2sbuf_p1_rd_en;
  assign _0558_ = dc2sbuf_p0_wr_sel_00 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1098" *) dc2sbuf_p1_wr_sel_00;
  assign _0559_ = _0558_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1099" *) wg2sbuf_p0_wr_sel_00;
  assign _0560_ = _0559_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1100" *) wg2sbuf_p1_wr_sel_00;
  assign _0561_ = _0560_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1101" *) img2sbuf_p0_wr_sel_00;
  assign sbuf_we_00 = _0561_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1102" *) img2sbuf_p1_wr_sel_00;
  assign _0562_ = dc2sbuf_p0_wr_sel_01 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1113" *) dc2sbuf_p1_wr_sel_01;
  assign _0563_ = _0562_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1114" *) wg2sbuf_p0_wr_sel_01;
  assign _0564_ = _0563_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1115" *) wg2sbuf_p1_wr_sel_01;
  assign _0565_ = _0564_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1116" *) img2sbuf_p0_wr_sel_01;
  assign sbuf_we_01 = _0565_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1117" *) img2sbuf_p1_wr_sel_01;
  assign _0566_ = dc2sbuf_p0_wr_sel_02 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1128" *) dc2sbuf_p1_wr_sel_02;
  assign _0567_ = _0566_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1129" *) wg2sbuf_p0_wr_sel_02;
  assign _0568_ = _0567_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1130" *) wg2sbuf_p1_wr_sel_02;
  assign _0569_ = _0568_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1131" *) img2sbuf_p0_wr_sel_02;
  assign sbuf_we_02 = _0569_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1132" *) img2sbuf_p1_wr_sel_02;
  assign _0570_ = dc2sbuf_p0_wr_sel_03 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1143" *) dc2sbuf_p1_wr_sel_03;
  assign _0571_ = _0570_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1144" *) wg2sbuf_p0_wr_sel_03;
  assign _0572_ = _0571_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1145" *) wg2sbuf_p1_wr_sel_03;
  assign _0573_ = _0572_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1146" *) img2sbuf_p0_wr_sel_03;
  assign sbuf_we_03 = _0573_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1147" *) img2sbuf_p1_wr_sel_03;
  assign _0574_ = dc2sbuf_p0_wr_sel_04 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1158" *) dc2sbuf_p1_wr_sel_04;
  assign _0575_ = _0574_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1159" *) wg2sbuf_p0_wr_sel_04;
  assign _0576_ = _0575_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1160" *) wg2sbuf_p1_wr_sel_04;
  assign _0577_ = _0576_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1161" *) img2sbuf_p0_wr_sel_04;
  assign sbuf_we_04 = _0577_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1162" *) img2sbuf_p1_wr_sel_04;
  assign _0578_ = dc2sbuf_p0_wr_sel_05 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1173" *) dc2sbuf_p1_wr_sel_05;
  assign _0579_ = _0578_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1174" *) wg2sbuf_p0_wr_sel_05;
  assign _0580_ = _0579_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1175" *) wg2sbuf_p1_wr_sel_05;
  assign _0581_ = _0580_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1176" *) img2sbuf_p0_wr_sel_05;
  assign sbuf_we_05 = _0581_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1177" *) img2sbuf_p1_wr_sel_05;
  assign _0582_ = dc2sbuf_p0_wr_sel_06 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1188" *) dc2sbuf_p1_wr_sel_06;
  assign _0583_ = _0582_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1189" *) wg2sbuf_p0_wr_sel_06;
  assign _0584_ = _0583_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1190" *) wg2sbuf_p1_wr_sel_06;
  assign _0585_ = _0584_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1191" *) img2sbuf_p0_wr_sel_06;
  assign sbuf_we_06 = _0585_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1192" *) img2sbuf_p1_wr_sel_06;
  assign _0586_ = dc2sbuf_p0_wr_sel_07 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1203" *) dc2sbuf_p1_wr_sel_07;
  assign _0587_ = _0586_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1204" *) wg2sbuf_p0_wr_sel_07;
  assign _0588_ = _0587_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1205" *) wg2sbuf_p1_wr_sel_07;
  assign _0589_ = _0588_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1206" *) img2sbuf_p0_wr_sel_07;
  assign sbuf_we_07 = _0589_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1207" *) img2sbuf_p1_wr_sel_07;
  assign _0590_ = dc2sbuf_p0_wr_sel_08 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1218" *) dc2sbuf_p1_wr_sel_08;
  assign _0591_ = _0590_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1219" *) wg2sbuf_p0_wr_sel_08;
  assign _0592_ = _0591_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1220" *) wg2sbuf_p1_wr_sel_08;
  assign _0593_ = _0592_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1221" *) img2sbuf_p0_wr_sel_08;
  assign sbuf_we_08 = _0593_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1222" *) img2sbuf_p1_wr_sel_08;
  assign _0594_ = dc2sbuf_p0_wr_sel_09 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1233" *) dc2sbuf_p1_wr_sel_09;
  assign _0595_ = _0594_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1234" *) wg2sbuf_p0_wr_sel_09;
  assign _0596_ = _0595_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1235" *) wg2sbuf_p1_wr_sel_09;
  assign _0597_ = _0596_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1236" *) img2sbuf_p0_wr_sel_09;
  assign sbuf_we_09 = _0597_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1237" *) img2sbuf_p1_wr_sel_09;
  assign _0598_ = dc2sbuf_p0_wr_sel_10 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1248" *) dc2sbuf_p1_wr_sel_10;
  assign _0599_ = _0598_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1249" *) wg2sbuf_p0_wr_sel_10;
  assign _0600_ = _0599_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1250" *) wg2sbuf_p1_wr_sel_10;
  assign _0601_ = _0600_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1251" *) img2sbuf_p0_wr_sel_10;
  assign sbuf_we_10 = _0601_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1252" *) img2sbuf_p1_wr_sel_10;
  assign _0602_ = dc2sbuf_p0_wr_sel_11 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1263" *) dc2sbuf_p1_wr_sel_11;
  assign _0603_ = _0602_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1264" *) wg2sbuf_p0_wr_sel_11;
  assign _0604_ = _0603_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1265" *) wg2sbuf_p1_wr_sel_11;
  assign _0605_ = _0604_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1266" *) img2sbuf_p0_wr_sel_11;
  assign sbuf_we_11 = _0605_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1267" *) img2sbuf_p1_wr_sel_11;
  assign _0606_ = dc2sbuf_p0_wr_sel_12 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1278" *) dc2sbuf_p1_wr_sel_12;
  assign _0607_ = _0606_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1279" *) wg2sbuf_p0_wr_sel_12;
  assign _0608_ = _0607_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1280" *) wg2sbuf_p1_wr_sel_12;
  assign _0609_ = _0608_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1281" *) img2sbuf_p0_wr_sel_12;
  assign sbuf_we_12 = _0609_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1282" *) img2sbuf_p1_wr_sel_12;
  assign _0610_ = dc2sbuf_p0_wr_sel_13 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1293" *) dc2sbuf_p1_wr_sel_13;
  assign _0611_ = _0610_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1294" *) wg2sbuf_p0_wr_sel_13;
  assign _0612_ = _0611_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1295" *) wg2sbuf_p1_wr_sel_13;
  assign _0613_ = _0612_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1296" *) img2sbuf_p0_wr_sel_13;
  assign sbuf_we_13 = _0613_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1297" *) img2sbuf_p1_wr_sel_13;
  assign _0614_ = dc2sbuf_p0_wr_sel_14 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1308" *) dc2sbuf_p1_wr_sel_14;
  assign _0615_ = _0614_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1309" *) wg2sbuf_p0_wr_sel_14;
  assign _0616_ = _0615_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1310" *) wg2sbuf_p1_wr_sel_14;
  assign _0617_ = _0616_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1311" *) img2sbuf_p0_wr_sel_14;
  assign sbuf_we_14 = _0617_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1312" *) img2sbuf_p1_wr_sel_14;
  assign _0618_ = dc2sbuf_p0_wr_sel_15 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1323" *) dc2sbuf_p1_wr_sel_15;
  assign _0619_ = _0618_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1324" *) wg2sbuf_p0_wr_sel_15;
  assign _0620_ = _0619_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1325" *) wg2sbuf_p1_wr_sel_15;
  assign _0621_ = _0620_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1326" *) img2sbuf_p0_wr_sel_15;
  assign sbuf_we_15 = _0621_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1327" *) img2sbuf_p1_wr_sel_15;
  assign _0622_ = _0044_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1344" *) _0045_;
  assign _0623_ = _0622_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1345" *) _0046_;
  assign _0624_ = _0623_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1346" *) _0047_;
  assign _0625_ = _0624_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1347" *) _0048_;
  assign sbuf_wa_00 = _0625_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1348" *) _0049_;
  assign _0626_ = _0050_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1365" *) _0051_;
  assign _0627_ = _0626_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1366" *) _0052_;
  assign _0628_ = _0627_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1367" *) _0053_;
  assign _0629_ = _0628_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1368" *) _0054_;
  assign sbuf_wa_01 = _0629_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1369" *) _0055_;
  assign _0630_ = _0056_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1386" *) _0057_;
  assign _0631_ = _0630_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1387" *) _0058_;
  assign _0632_ = _0631_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1388" *) _0059_;
  assign _0633_ = _0632_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1389" *) _0060_;
  assign sbuf_wa_02 = _0633_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1390" *) _0061_;
  assign _0634_ = _0062_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1407" *) _0063_;
  assign _0635_ = _0634_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1408" *) _0064_;
  assign _0636_ = _0635_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1409" *) _0065_;
  assign _0637_ = _0636_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1410" *) _0066_;
  assign sbuf_wa_03 = _0637_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1411" *) _0067_;
  assign _0638_ = _0068_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1428" *) _0069_;
  assign _0639_ = _0638_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1429" *) _0070_;
  assign _0640_ = _0639_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1430" *) _0071_;
  assign _0641_ = _0640_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1431" *) _0072_;
  assign sbuf_wa_04 = _0641_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1432" *) _0073_;
  assign _0642_ = _0074_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1449" *) _0075_;
  assign _0643_ = _0642_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1450" *) _0076_;
  assign _0644_ = _0643_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1451" *) _0077_;
  assign _0645_ = _0644_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1452" *) _0078_;
  assign sbuf_wa_05 = _0645_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1453" *) _0079_;
  assign _0646_ = _0080_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1470" *) _0081_;
  assign _0647_ = _0646_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1471" *) _0082_;
  assign _0648_ = _0647_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1472" *) _0083_;
  assign _0649_ = _0648_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1473" *) _0084_;
  assign sbuf_wa_06 = _0649_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1474" *) _0085_;
  assign _0650_ = _0086_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1491" *) _0087_;
  assign _0651_ = _0650_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1492" *) _0088_;
  assign _0652_ = _0651_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1493" *) _0089_;
  assign _0653_ = _0652_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1494" *) _0090_;
  assign sbuf_wa_07 = _0653_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1495" *) _0091_;
  assign _0654_ = _0092_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1512" *) _0093_;
  assign _0655_ = _0654_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1513" *) _0094_;
  assign _0656_ = _0655_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1514" *) _0095_;
  assign _0657_ = _0656_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1515" *) _0096_;
  assign sbuf_wa_08 = _0657_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1516" *) _0097_;
  assign _0658_ = _0098_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1533" *) _0099_;
  assign _0659_ = _0658_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1534" *) _0100_;
  assign _0660_ = _0659_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1535" *) _0101_;
  assign _0661_ = _0660_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1536" *) _0102_;
  assign sbuf_wa_09 = _0661_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1537" *) _0103_;
  assign _0662_ = _0104_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1554" *) _0105_;
  assign _0663_ = _0662_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1555" *) _0106_;
  assign _0664_ = _0663_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1556" *) _0107_;
  assign _0665_ = _0664_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1557" *) _0108_;
  assign sbuf_wa_10 = _0665_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1558" *) _0109_;
  assign _0666_ = _0110_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1575" *) _0111_;
  assign _0667_ = _0666_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1576" *) _0112_;
  assign _0668_ = _0667_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1577" *) _0113_;
  assign _0669_ = _0668_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1578" *) _0114_;
  assign sbuf_wa_11 = _0669_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1579" *) _0115_;
  assign _0670_ = _0116_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1596" *) _0117_;
  assign _0671_ = _0670_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1597" *) _0118_;
  assign _0672_ = _0671_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1598" *) _0119_;
  assign _0673_ = _0672_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1599" *) _0120_;
  assign sbuf_wa_12 = _0673_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1600" *) _0121_;
  assign _0674_ = _0122_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1617" *) _0123_;
  assign _0675_ = _0674_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1618" *) _0124_;
  assign _0676_ = _0675_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1619" *) _0125_;
  assign _0677_ = _0676_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1620" *) _0126_;
  assign sbuf_wa_13 = _0677_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1621" *) _0127_;
  assign _0678_ = _0128_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1638" *) _0129_;
  assign _0679_ = _0678_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1639" *) _0130_;
  assign _0680_ = _0679_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1640" *) _0131_;
  assign _0681_ = _0680_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1641" *) _0132_;
  assign sbuf_wa_14 = _0681_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1642" *) _0133_;
  assign _0682_ = _0134_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1659" *) _0135_;
  assign _0683_ = _0682_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1660" *) _0136_;
  assign _0684_ = _0683_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1661" *) _0137_;
  assign _0685_ = _0684_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1662" *) _0138_;
  assign sbuf_wa_15 = _0685_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1663" *) _0139_;
  assign _0686_ = _0140_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1680" *) _0141_;
  assign _0687_ = _0686_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1681" *) _0142_;
  assign _0688_ = _0687_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1682" *) _0143_;
  assign _0689_ = _0688_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1683" *) _0144_;
  assign sbuf_wdat_00 = _0689_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1684" *) _0145_;
  assign _0690_ = _0146_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1701" *) _0147_;
  assign _0691_ = _0690_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1702" *) _0148_;
  assign _0692_ = _0691_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1703" *) _0149_;
  assign _0693_ = _0692_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1704" *) _0150_;
  assign sbuf_wdat_01 = _0693_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1705" *) _0151_;
  assign _0694_ = _0152_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1722" *) _0153_;
  assign _0695_ = _0694_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1723" *) _0154_;
  assign _0696_ = _0695_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1724" *) _0155_;
  assign _0697_ = _0696_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1725" *) _0156_;
  assign sbuf_wdat_02 = _0697_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1726" *) _0157_;
  assign _0698_ = _0158_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1743" *) _0159_;
  assign _0699_ = _0698_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1744" *) _0160_;
  assign _0700_ = _0699_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1745" *) _0161_;
  assign _0701_ = _0700_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1746" *) _0162_;
  assign sbuf_wdat_03 = _0701_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1747" *) _0163_;
  assign _0702_ = _0164_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1764" *) _0165_;
  assign _0703_ = _0702_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1765" *) _0166_;
  assign _0704_ = _0703_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1766" *) _0167_;
  assign _0705_ = _0704_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1767" *) _0168_;
  assign sbuf_wdat_04 = _0705_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1768" *) _0169_;
  assign _0706_ = _0170_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1785" *) _0171_;
  assign _0707_ = _0706_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1786" *) _0172_;
  assign _0708_ = _0707_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1787" *) _0173_;
  assign _0709_ = _0708_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1788" *) _0174_;
  assign sbuf_wdat_05 = _0709_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1789" *) _0175_;
  assign _0710_ = _0176_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1806" *) _0177_;
  assign _0711_ = _0710_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1807" *) _0178_;
  assign _0712_ = _0711_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1808" *) _0179_;
  assign _0713_ = _0712_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1809" *) _0180_;
  assign sbuf_wdat_06 = _0713_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1810" *) _0181_;
  assign _0714_ = _0182_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1827" *) _0183_;
  assign _0715_ = _0714_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1828" *) _0184_;
  assign _0716_ = _0715_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1829" *) _0185_;
  assign _0717_ = _0716_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1830" *) _0186_;
  assign sbuf_wdat_07 = _0717_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1831" *) _0187_;
  assign _0718_ = _0188_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1848" *) _0189_;
  assign _0719_ = _0718_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1849" *) _0190_;
  assign _0720_ = _0719_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1850" *) _0191_;
  assign _0721_ = _0720_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1851" *) _0192_;
  assign sbuf_wdat_08 = _0721_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1852" *) _0193_;
  assign _0722_ = _0194_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1869" *) _0195_;
  assign _0723_ = _0722_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1870" *) _0196_;
  assign _0724_ = _0723_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1871" *) _0197_;
  assign _0725_ = _0724_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1872" *) _0198_;
  assign sbuf_wdat_09 = _0725_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1873" *) _0199_;
  assign _0726_ = _0200_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1890" *) _0201_;
  assign _0727_ = _0726_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1891" *) _0202_;
  assign _0728_ = _0727_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1892" *) _0203_;
  assign _0729_ = _0728_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1893" *) _0204_;
  assign sbuf_wdat_10 = _0729_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1894" *) _0205_;
  assign _0730_ = _0206_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1911" *) _0207_;
  assign _0731_ = _0730_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1912" *) _0208_;
  assign _0732_ = _0731_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1913" *) _0209_;
  assign _0733_ = _0732_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1914" *) _0210_;
  assign sbuf_wdat_11 = _0733_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1915" *) _0211_;
  assign _0734_ = _0212_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1932" *) _0213_;
  assign _0735_ = _0734_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1933" *) _0214_;
  assign _0736_ = _0735_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1934" *) _0215_;
  assign _0737_ = _0736_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1935" *) _0216_;
  assign sbuf_wdat_12 = _0737_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1936" *) _0217_;
  assign _0738_ = _0218_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1953" *) _0219_;
  assign _0739_ = _0738_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1954" *) _0220_;
  assign _0740_ = _0739_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1955" *) _0221_;
  assign _0741_ = _0740_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1956" *) _0222_;
  assign sbuf_wdat_13 = _0741_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1957" *) _0223_;
  assign _0742_ = _0224_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1974" *) _0225_;
  assign _0743_ = _0742_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1975" *) _0226_;
  assign _0744_ = _0743_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1976" *) _0227_;
  assign _0745_ = _0744_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1977" *) _0228_;
  assign sbuf_wdat_14 = _0745_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1978" *) _0229_;
  assign _0746_ = _0230_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1995" *) _0231_;
  assign _0747_ = _0746_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1996" *) _0232_;
  assign _0748_ = _0747_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1997" *) _0233_;
  assign _0749_ = _0748_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1998" *) _0234_;
  assign sbuf_wdat_15 = _0749_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:1999" *) _0235_;
  assign _0750_ = dc2sbuf_p0_rd_sel_00 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2754" *) wg2sbuf_p0_rd_sel_00;
  assign sbuf_p0_re_00 = _0750_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2754" *) img2sbuf_p0_rd_sel_00;
  assign _0751_ = dc2sbuf_p1_rd_sel_00 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2761" *) wg2sbuf_p1_rd_sel_00;
  assign sbuf_p1_re_00 = _0751_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2761" *) img2sbuf_p1_rd_sel_00;
  assign _0752_ = dc2sbuf_p0_rd_sel_01 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2768" *) wg2sbuf_p0_rd_sel_00;
  assign sbuf_p0_re_01 = _0752_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2768" *) img2sbuf_p0_rd_sel_01;
  assign _0753_ = dc2sbuf_p1_rd_sel_01 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2775" *) wg2sbuf_p1_rd_sel_00;
  assign sbuf_p1_re_01 = _0753_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2775" *) img2sbuf_p1_rd_sel_01;
  assign _0754_ = dc2sbuf_p0_rd_sel_02 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2782" *) wg2sbuf_p0_rd_sel_00;
  assign sbuf_p0_re_02 = _0754_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2782" *) img2sbuf_p0_rd_sel_02;
  assign _0755_ = dc2sbuf_p1_rd_sel_02 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2789" *) wg2sbuf_p1_rd_sel_00;
  assign sbuf_p1_re_02 = _0755_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2789" *) img2sbuf_p1_rd_sel_02;
  assign _0756_ = dc2sbuf_p0_rd_sel_03 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2796" *) wg2sbuf_p0_rd_sel_00;
  assign sbuf_p0_re_03 = _0756_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2796" *) img2sbuf_p0_rd_sel_03;
  assign _0757_ = dc2sbuf_p1_rd_sel_03 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2803" *) wg2sbuf_p1_rd_sel_00;
  assign sbuf_p1_re_03 = _0757_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2803" *) img2sbuf_p1_rd_sel_03;
  assign _0758_ = dc2sbuf_p0_rd_sel_04 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2810" *) wg2sbuf_p0_rd_sel_04;
  assign sbuf_p0_re_04 = _0758_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2810" *) img2sbuf_p0_rd_sel_04;
  assign _0759_ = dc2sbuf_p1_rd_sel_04 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2817" *) wg2sbuf_p1_rd_sel_04;
  assign sbuf_p1_re_04 = _0759_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2817" *) img2sbuf_p1_rd_sel_04;
  assign _0760_ = dc2sbuf_p0_rd_sel_05 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2824" *) wg2sbuf_p0_rd_sel_04;
  assign sbuf_p0_re_05 = _0760_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2824" *) img2sbuf_p0_rd_sel_05;
  assign _0761_ = dc2sbuf_p1_rd_sel_05 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2831" *) wg2sbuf_p1_rd_sel_04;
  assign sbuf_p1_re_05 = _0761_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2831" *) img2sbuf_p1_rd_sel_05;
  assign _0762_ = dc2sbuf_p0_rd_sel_06 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2838" *) wg2sbuf_p0_rd_sel_04;
  assign sbuf_p0_re_06 = _0762_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2838" *) img2sbuf_p0_rd_sel_06;
  assign _0763_ = dc2sbuf_p1_rd_sel_06 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2845" *) wg2sbuf_p1_rd_sel_04;
  assign sbuf_p1_re_06 = _0763_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2845" *) img2sbuf_p1_rd_sel_06;
  assign _0764_ = dc2sbuf_p0_rd_sel_07 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2852" *) wg2sbuf_p0_rd_sel_04;
  assign sbuf_p0_re_07 = _0764_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2852" *) img2sbuf_p0_rd_sel_07;
  assign _0765_ = dc2sbuf_p1_rd_sel_07 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2859" *) wg2sbuf_p1_rd_sel_04;
  assign sbuf_p1_re_07 = _0765_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2859" *) img2sbuf_p1_rd_sel_07;
  assign _0766_ = dc2sbuf_p0_rd_sel_08 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2866" *) wg2sbuf_p0_rd_sel_08;
  assign sbuf_p0_re_08 = _0766_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2866" *) img2sbuf_p0_rd_sel_08;
  assign _0767_ = dc2sbuf_p1_rd_sel_08 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2873" *) wg2sbuf_p1_rd_sel_08;
  assign sbuf_p1_re_08 = _0767_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2873" *) img2sbuf_p1_rd_sel_08;
  assign _0768_ = dc2sbuf_p0_rd_sel_09 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2880" *) wg2sbuf_p0_rd_sel_08;
  assign sbuf_p0_re_09 = _0768_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2880" *) img2sbuf_p0_rd_sel_09;
  assign _0769_ = dc2sbuf_p1_rd_sel_09 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2887" *) wg2sbuf_p1_rd_sel_08;
  assign sbuf_p1_re_09 = _0769_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2887" *) img2sbuf_p1_rd_sel_09;
  assign _0770_ = dc2sbuf_p0_rd_sel_10 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2894" *) wg2sbuf_p0_rd_sel_08;
  assign sbuf_p0_re_10 = _0770_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2894" *) img2sbuf_p0_rd_sel_10;
  assign _0771_ = dc2sbuf_p1_rd_sel_10 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2901" *) wg2sbuf_p1_rd_sel_08;
  assign sbuf_p1_re_10 = _0771_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2901" *) img2sbuf_p1_rd_sel_10;
  assign _0772_ = dc2sbuf_p0_rd_sel_11 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2908" *) wg2sbuf_p0_rd_sel_08;
  assign sbuf_p0_re_11 = _0772_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2908" *) img2sbuf_p0_rd_sel_11;
  assign _0773_ = dc2sbuf_p1_rd_sel_11 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2915" *) wg2sbuf_p1_rd_sel_08;
  assign sbuf_p1_re_11 = _0773_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2915" *) img2sbuf_p1_rd_sel_11;
  assign _0774_ = dc2sbuf_p0_rd_sel_12 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2922" *) wg2sbuf_p0_rd_sel_12;
  assign sbuf_p0_re_12 = _0774_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2922" *) img2sbuf_p0_rd_sel_12;
  assign _0775_ = dc2sbuf_p1_rd_sel_12 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2929" *) wg2sbuf_p1_rd_sel_12;
  assign sbuf_p1_re_12 = _0775_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2929" *) img2sbuf_p1_rd_sel_12;
  assign _0776_ = dc2sbuf_p0_rd_sel_13 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2936" *) wg2sbuf_p0_rd_sel_12;
  assign sbuf_p0_re_13 = _0776_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2936" *) img2sbuf_p0_rd_sel_13;
  assign _0777_ = dc2sbuf_p1_rd_sel_13 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2943" *) wg2sbuf_p1_rd_sel_12;
  assign sbuf_p1_re_13 = _0777_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2943" *) img2sbuf_p1_rd_sel_13;
  assign _0778_ = dc2sbuf_p0_rd_sel_14 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2950" *) wg2sbuf_p0_rd_sel_12;
  assign sbuf_p0_re_14 = _0778_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2950" *) img2sbuf_p0_rd_sel_14;
  assign _0779_ = dc2sbuf_p1_rd_sel_14 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2957" *) wg2sbuf_p1_rd_sel_12;
  assign sbuf_p1_re_14 = _0779_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2957" *) img2sbuf_p1_rd_sel_14;
  assign _0780_ = dc2sbuf_p0_rd_sel_15 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2964" *) wg2sbuf_p0_rd_sel_12;
  assign sbuf_p0_re_15 = _0780_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2964" *) img2sbuf_p0_rd_sel_15;
  assign _0781_ = dc2sbuf_p1_rd_sel_15 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2971" *) wg2sbuf_p1_rd_sel_12;
  assign sbuf_p1_re_15 = _0781_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2971" *) img2sbuf_p1_rd_sel_15;
  assign sbuf_re_00 = sbuf_p0_re_00 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2977" *) sbuf_p1_re_00;
  assign sbuf_re_01 = sbuf_p0_re_01 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2983" *) sbuf_p1_re_01;
  assign sbuf_re_02 = sbuf_p0_re_02 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2989" *) sbuf_p1_re_02;
  assign sbuf_re_03 = sbuf_p0_re_03 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2995" *) sbuf_p1_re_03;
  assign sbuf_re_04 = sbuf_p0_re_04 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3001" *) sbuf_p1_re_04;
  assign sbuf_re_05 = sbuf_p0_re_05 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3007" *) sbuf_p1_re_05;
  assign sbuf_re_06 = sbuf_p0_re_06 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3013" *) sbuf_p1_re_06;
  assign sbuf_re_07 = sbuf_p0_re_07 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3019" *) sbuf_p1_re_07;
  assign sbuf_re_08 = sbuf_p0_re_08 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3025" *) sbuf_p1_re_08;
  assign sbuf_re_09 = sbuf_p0_re_09 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3031" *) sbuf_p1_re_09;
  assign sbuf_re_10 = sbuf_p0_re_10 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3037" *) sbuf_p1_re_10;
  assign sbuf_re_11 = sbuf_p0_re_11 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3043" *) sbuf_p1_re_11;
  assign sbuf_re_12 = sbuf_p0_re_12 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3049" *) sbuf_p1_re_12;
  assign sbuf_re_13 = sbuf_p0_re_13 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3055" *) sbuf_p1_re_13;
  assign sbuf_re_14 = sbuf_p0_re_14 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3061" *) sbuf_p1_re_14;
  assign sbuf_re_15 = sbuf_p0_re_15 | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3067" *) sbuf_p1_re_15;
  assign _0782_ = _0236_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3090" *) _0237_;
  assign _0783_ = _0782_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3091" *) _0238_;
  assign _0784_ = _0783_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3092" *) _0239_;
  assign _0785_ = _0784_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3093" *) _0240_;
  assign sbuf_ra_00 = _0785_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3094" *) _0241_;
  assign _0786_ = _0242_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3111" *) _0243_;
  assign _0787_ = _0786_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3112" *) _0238_;
  assign _0788_ = _0787_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3113" *) _0239_;
  assign _0789_ = _0788_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3114" *) _0244_;
  assign sbuf_ra_01 = _0789_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3115" *) _0245_;
  assign _0790_ = _0246_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3132" *) _0247_;
  assign _0791_ = _0790_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3133" *) _0238_;
  assign _0792_ = _0791_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3134" *) _0239_;
  assign _0793_ = _0792_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3135" *) _0248_;
  assign sbuf_ra_02 = _0793_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3136" *) _0249_;
  assign _0794_ = _0250_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3153" *) _0251_;
  assign _0795_ = _0794_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3154" *) _0238_;
  assign _0796_ = _0795_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3155" *) _0239_;
  assign _0797_ = _0796_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3156" *) _0252_;
  assign sbuf_ra_03 = _0797_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3157" *) _0253_;
  assign _0798_ = _0254_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3174" *) _0255_;
  assign _0799_ = _0798_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3175" *) _0256_;
  assign _0800_ = _0799_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3176" *) _0257_;
  assign _0801_ = _0800_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3177" *) _0258_;
  assign sbuf_ra_04 = _0801_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3178" *) _0259_;
  assign _0802_ = _0260_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3195" *) _0261_;
  assign _0803_ = _0802_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3196" *) _0256_;
  assign _0804_ = _0803_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3197" *) _0257_;
  assign _0805_ = _0804_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3198" *) _0262_;
  assign sbuf_ra_05 = _0805_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3199" *) _0263_;
  assign _0806_ = _0264_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3216" *) _0265_;
  assign _0807_ = _0806_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3217" *) _0256_;
  assign _0808_ = _0807_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3218" *) _0257_;
  assign _0809_ = _0808_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3219" *) _0266_;
  assign sbuf_ra_06 = _0809_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3220" *) _0267_;
  assign _0810_ = _0268_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3237" *) _0269_;
  assign _0811_ = _0810_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3238" *) _0256_;
  assign _0812_ = _0811_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3239" *) _0257_;
  assign _0813_ = _0812_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3240" *) _0270_;
  assign sbuf_ra_07 = _0813_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3241" *) _0271_;
  assign _0814_ = _0272_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3258" *) _0273_;
  assign _0815_ = _0814_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3259" *) _0274_;
  assign _0816_ = _0815_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3260" *) _0275_;
  assign _0817_ = _0816_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3261" *) _0276_;
  assign sbuf_ra_08 = _0817_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3262" *) _0277_;
  assign _0818_ = _0278_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3279" *) _0279_;
  assign _0819_ = _0818_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3280" *) _0274_;
  assign _0820_ = _0819_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3281" *) _0275_;
  assign _0821_ = _0820_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3282" *) _0280_;
  assign sbuf_ra_09 = _0821_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3283" *) _0281_;
  assign _0822_ = _0282_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3300" *) _0283_;
  assign _0823_ = _0822_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3301" *) _0274_;
  assign _0824_ = _0823_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3302" *) _0275_;
  assign _0825_ = _0824_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3303" *) _0284_;
  assign sbuf_ra_10 = _0825_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3304" *) _0285_;
  assign _0826_ = _0286_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3321" *) _0287_;
  assign _0827_ = _0826_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3322" *) _0274_;
  assign _0828_ = _0827_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3323" *) _0275_;
  assign _0829_ = _0828_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3324" *) _0288_;
  assign sbuf_ra_11 = _0829_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3325" *) _0289_;
  assign _0830_ = _0290_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3342" *) _0291_;
  assign _0831_ = _0830_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3343" *) _0292_;
  assign _0832_ = _0831_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3344" *) _0293_;
  assign _0833_ = _0832_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3345" *) _0294_;
  assign sbuf_ra_12 = _0833_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3346" *) _0295_;
  assign _0834_ = _0296_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3363" *) _0297_;
  assign _0835_ = _0834_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3364" *) _0292_;
  assign _0836_ = _0835_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3365" *) _0293_;
  assign _0837_ = _0836_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3366" *) _0298_;
  assign sbuf_ra_13 = _0837_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3367" *) _0299_;
  assign _0838_ = _0300_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3384" *) _0301_;
  assign _0839_ = _0838_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3385" *) _0292_;
  assign _0840_ = _0839_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3386" *) _0293_;
  assign _0841_ = _0840_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3387" *) _0302_;
  assign sbuf_ra_14 = _0841_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3388" *) _0303_;
  assign _0842_ = _0304_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3405" *) _0305_;
  assign _0843_ = _0842_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3406" *) _0292_;
  assign _0844_ = _0843_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3407" *) _0293_;
  assign _0845_ = _0844_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3408" *) _0306_;
  assign sbuf_ra_15 = _0845_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3409" *) _0307_;
  assign _0846_ = dc2sbuf_p0_rd_en | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3802" *) wg2sbuf_p0_rd_en;
  assign _0000_ = _0846_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3802" *) img2sbuf_p0_rd_en;
  assign _0847_ = dc2sbuf_p1_rd_en | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3809" *) wg2sbuf_p1_rd_en;
  assign _0022_ = _0847_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3809" *) img2sbuf_p1_rd_en;
  assign _0848_ = _0308_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3850" *) _0309_;
  assign _0849_ = _0848_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3851" *) _0310_;
  assign _0850_ = _0849_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3852" *) _0311_;
  assign _0851_ = _0850_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3853" *) _0312_;
  assign _0852_ = _0851_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3854" *) _0313_;
  assign _0853_ = _0852_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3855" *) _0314_;
  assign _0854_ = _0853_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3856" *) _0315_;
  assign _0855_ = _0854_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3857" *) _0316_;
  assign _0856_ = _0855_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3858" *) _0317_;
  assign _0857_ = _0856_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3859" *) _0318_;
  assign _0858_ = _0857_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3860" *) _0319_;
  assign _0859_ = _0858_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3861" *) _0320_;
  assign _0860_ = _0859_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3862" *) _0321_;
  assign _0861_ = _0860_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3863" *) _0322_;
  assign sbuf_p0_norm_rdat = _0861_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3864" *) _0323_;
  assign _0862_ = _0324_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3901" *) _0325_;
  assign _0863_ = _0862_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3902" *) _0326_;
  assign _0864_ = _0863_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3903" *) _0327_;
  assign _0865_ = _0864_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3904" *) _0328_;
  assign _0866_ = _0865_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3905" *) _0329_;
  assign _0867_ = _0866_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3906" *) _0330_;
  assign _0868_ = _0867_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3907" *) _0331_;
  assign _0869_ = _0868_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3908" *) _0332_;
  assign _0870_ = _0869_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3909" *) _0333_;
  assign _0871_ = _0870_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3910" *) _0334_;
  assign _0872_ = _0871_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3911" *) _0335_;
  assign _0873_ = _0872_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3912" *) _0336_;
  assign _0874_ = _0873_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3913" *) _0337_;
  assign _0875_ = _0874_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3914" *) _0338_;
  assign sbuf_p1_norm_rdat = _0875_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3915" *) _0339_;
  assign _0876_ = _0340_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3928" *) _0341_;
  assign _0877_ = _0876_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3929" *) _0342_;
  assign sbuf_p0_wg_rdat_src_0 = _0877_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3930" *) _0343_;
  assign _0878_ = _0344_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3943" *) _0345_;
  assign _0879_ = _0878_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3944" *) _0346_;
  assign sbuf_p0_wg_rdat_src_1 = _0879_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3945" *) _0347_;
  assign _0880_ = _0348_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3958" *) _0349_;
  assign _0881_ = _0880_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3959" *) _0350_;
  assign sbuf_p0_wg_rdat_src_2 = _0881_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3960" *) _0351_;
  assign _0882_ = _0352_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3973" *) _0353_;
  assign _0883_ = _0882_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3974" *) _0354_;
  assign sbuf_p0_wg_rdat_src_3 = _0883_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3975" *) _0355_;
  assign _0884_ = _0356_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3988" *) _0357_;
  assign _0885_ = _0884_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3989" *) _0358_;
  assign sbuf_p1_wg_rdat_src_0 = _0885_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:3990" *) _0359_;
  assign _0886_ = _0360_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4003" *) _0361_;
  assign _0887_ = _0886_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4004" *) _0362_;
  assign sbuf_p1_wg_rdat_src_1 = _0887_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4005" *) _0363_;
  assign _0888_ = _0364_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4018" *) _0365_;
  assign _0889_ = _0888_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4019" *) _0366_;
  assign sbuf_p1_wg_rdat_src_2 = _0889_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4020" *) _0367_;
  assign _0890_ = _0368_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4033" *) _0369_;
  assign _0891_ = _0890_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4034" *) _0370_;
  assign sbuf_p1_wg_rdat_src_3 = _0891_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4035" *) _0371_;
  assign _0892_ = _0372_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4048" *) _0373_;
  assign _0893_ = _0892_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4049" *) _0374_;
  assign sbuf_p0_wg_rdat = _0893_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4050" *) _0375_;
  assign _0894_ = _0376_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4063" *) _0377_;
  assign _0895_ = _0894_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4064" *) _0378_;
  assign sbuf_p1_wg_rdat = _0895_ | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4065" *) _0379_;
  assign sbuf_p0_rdat = sbuf_p0_norm_rdat | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4071" *) sbuf_p0_wg_rdat;
  assign sbuf_p1_rdat = sbuf_p1_norm_rdat | (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4077" *) sbuf_p1_wg_rdat;
  always @(posedge nvdla_core_clk)
      sbuf_p1_rdat_d2 <= _0023_;
  always @(posedge nvdla_core_clk)
      sbuf_p0_rdat_d2 <= _0001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_rd_en_d1 <= 1'b0;
    else
      sbuf_p1_rd_en_d1 <= _0022_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_rd_en_d1 <= 1'b0;
    else
      sbuf_p0_rd_en_d1 <= _0000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_wg_sel_q3_d1 <= 1'b0;
    else
      sbuf_p1_wg_sel_q3_d1 <= sbuf_p1_wg_sel_q3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_wg_sel_q2_d1 <= 1'b0;
    else
      sbuf_p1_wg_sel_q2_d1 <= sbuf_p1_wg_sel_q2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_wg_sel_q1_d1 <= 1'b0;
    else
      sbuf_p1_wg_sel_q1_d1 <= sbuf_p1_wg_sel_q1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_wg_sel_q0_d1 <= 1'b0;
    else
      sbuf_p1_wg_sel_q0_d1 <= sbuf_p1_wg_sel_q0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_wg_sel_q3_d1 <= 1'b0;
    else
      sbuf_p0_wg_sel_q3_d1 <= sbuf_p0_wg_sel_q3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_wg_sel_q2_d1 <= 1'b0;
    else
      sbuf_p0_wg_sel_q2_d1 <= sbuf_p0_wg_sel_q2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_wg_sel_q1_d1 <= 1'b0;
    else
      sbuf_p0_wg_sel_q1_d1 <= sbuf_p0_wg_sel_q1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_wg_sel_q0_d1 <= 1'b0;
    else
      sbuf_p0_wg_sel_q0_d1 <= sbuf_p0_wg_sel_q0;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_03_wg_d1 <= 1'b0;
    else
      sbuf_p1_re_03_wg_d1 <= _0031_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_03_wg_d1 <= 1'b0;
    else
      sbuf_p0_re_03_wg_d1 <= _0009_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_02_wg_d1 <= 1'b0;
    else
      sbuf_p1_re_02_wg_d1 <= _0029_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_02_wg_d1 <= 1'b0;
    else
      sbuf_p0_re_02_wg_d1 <= _0007_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_01_wg_d1 <= 1'b0;
    else
      sbuf_p1_re_01_wg_d1 <= _0027_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_01_wg_d1 <= 1'b0;
    else
      sbuf_p0_re_01_wg_d1 <= _0005_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_00_wg_d1 <= 1'b0;
    else
      sbuf_p1_re_00_wg_d1 <= _0025_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_00_wg_d1 <= 1'b0;
    else
      sbuf_p0_re_00_wg_d1 <= _0003_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_15_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_15_norm_d1 <= _0043_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_15_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_15_norm_d1 <= _0021_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_14_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_14_norm_d1 <= _0042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_14_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_14_norm_d1 <= _0020_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_13_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_13_norm_d1 <= _0041_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_13_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_13_norm_d1 <= _0019_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_12_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_12_norm_d1 <= _0040_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_12_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_12_norm_d1 <= _0018_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_11_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_11_norm_d1 <= _0039_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_11_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_11_norm_d1 <= _0017_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_10_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_10_norm_d1 <= _0038_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_10_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_10_norm_d1 <= _0016_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_09_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_09_norm_d1 <= _0037_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_09_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_09_norm_d1 <= _0015_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_08_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_08_norm_d1 <= _0036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_08_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_08_norm_d1 <= _0014_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_07_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_07_norm_d1 <= _0035_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_07_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_07_norm_d1 <= _0013_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_06_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_06_norm_d1 <= _0034_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_06_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_06_norm_d1 <= _0012_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_05_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_05_norm_d1 <= _0033_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_05_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_05_norm_d1 <= _0011_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_04_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_04_norm_d1 <= _0032_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_04_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_04_norm_d1 <= _0010_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_03_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_03_norm_d1 <= _0030_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_03_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_03_norm_d1 <= _0008_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_02_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_02_norm_d1 <= _0028_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_02_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_02_norm_d1 <= _0006_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_01_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_01_norm_d1 <= _0026_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_01_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_01_norm_d1 <= _0004_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p1_re_00_norm_d1 <= 1'b0;
    else
      sbuf_p1_re_00_norm_d1 <= _0024_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sbuf_p0_re_00_norm_d1 <= 1'b0;
    else
      sbuf_p0_re_00_norm_d1 <= _0002_;
  assign _0023_ = sbuf_p1_rd_en_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4093" *) sbuf_p1_rdat : sbuf_p1_rdat_d2;
  assign _0001_ = sbuf_p0_rd_en_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:4083" *) sbuf_p0_rdat : sbuf_p0_rdat_d2;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2004" *)
  nv_ram_rws_16x256 u_shared_buffer_00 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_00),
    .dout(sbuf_rdat_00),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_00),
    .re(sbuf_re_00),
    .wa(sbuf_wa_00),
    .we(sbuf_we_00)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2014" *)
  nv_ram_rws_16x256 u_shared_buffer_01 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_01),
    .dout(sbuf_rdat_01),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_01),
    .re(sbuf_re_01),
    .wa(sbuf_wa_01),
    .we(sbuf_we_01)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2024" *)
  nv_ram_rws_16x256 u_shared_buffer_02 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_02),
    .dout(sbuf_rdat_02),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_02),
    .re(sbuf_re_02),
    .wa(sbuf_wa_02),
    .we(sbuf_we_02)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2034" *)
  nv_ram_rws_16x256 u_shared_buffer_03 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_03),
    .dout(sbuf_rdat_03),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_03),
    .re(sbuf_re_03),
    .wa(sbuf_wa_03),
    .we(sbuf_we_03)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2044" *)
  nv_ram_rws_16x256 u_shared_buffer_04 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_04),
    .dout(sbuf_rdat_04),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_04),
    .re(sbuf_re_04),
    .wa(sbuf_wa_04),
    .we(sbuf_we_04)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2054" *)
  nv_ram_rws_16x256 u_shared_buffer_05 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_05),
    .dout(sbuf_rdat_05),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_05),
    .re(sbuf_re_05),
    .wa(sbuf_wa_05),
    .we(sbuf_we_05)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2064" *)
  nv_ram_rws_16x256 u_shared_buffer_06 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_06),
    .dout(sbuf_rdat_06),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_06),
    .re(sbuf_re_06),
    .wa(sbuf_wa_06),
    .we(sbuf_we_06)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2074" *)
  nv_ram_rws_16x256 u_shared_buffer_07 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_07),
    .dout(sbuf_rdat_07),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_07),
    .re(sbuf_re_07),
    .wa(sbuf_wa_07),
    .we(sbuf_we_07)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2084" *)
  nv_ram_rws_16x256 u_shared_buffer_08 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_08),
    .dout(sbuf_rdat_08),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_08),
    .re(sbuf_re_08),
    .wa(sbuf_wa_08),
    .we(sbuf_we_08)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2094" *)
  nv_ram_rws_16x256 u_shared_buffer_09 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_09),
    .dout(sbuf_rdat_09),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_09),
    .re(sbuf_re_09),
    .wa(sbuf_wa_09),
    .we(sbuf_we_09)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2104" *)
  nv_ram_rws_16x256 u_shared_buffer_10 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_10),
    .dout(sbuf_rdat_10),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_10),
    .re(sbuf_re_10),
    .wa(sbuf_wa_10),
    .we(sbuf_we_10)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2114" *)
  nv_ram_rws_16x256 u_shared_buffer_11 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_11),
    .dout(sbuf_rdat_11),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_11),
    .re(sbuf_re_11),
    .wa(sbuf_wa_11),
    .we(sbuf_we_11)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2124" *)
  nv_ram_rws_16x256 u_shared_buffer_12 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_12),
    .dout(sbuf_rdat_12),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_12),
    .re(sbuf_re_12),
    .wa(sbuf_wa_12),
    .we(sbuf_we_12)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2134" *)
  nv_ram_rws_16x256 u_shared_buffer_13 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_13),
    .dout(sbuf_rdat_13),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_13),
    .re(sbuf_re_13),
    .wa(sbuf_wa_13),
    .we(sbuf_we_13)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2144" *)
  nv_ram_rws_16x256 u_shared_buffer_14 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_14),
    .dout(sbuf_rdat_14),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_14),
    .re(sbuf_re_14),
    .wa(sbuf_wa_14),
    .we(sbuf_we_14)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cdma/NV_NVDLA_CDMA_shared_buffer.v:2154" *)
  nv_ram_rws_16x256 u_shared_buffer_15 (
    .clk(nvdla_core_clk),
    .di(sbuf_wdat_15),
    .dout(sbuf_rdat_15),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(sbuf_ra_15),
    .re(sbuf_re_15),
    .wa(sbuf_wa_15),
    .we(sbuf_we_15)
  );
  assign dc2sbuf_p0_rd_bsel = dc2sbuf_p0_rd_addr[7:4];
  assign dc2sbuf_p0_rd_data = sbuf_p0_rdat_d2;
  assign dc2sbuf_p0_rd_esel = dc2sbuf_p0_rd_addr[3:0];
  assign dc2sbuf_p0_wr_bsel = dc2sbuf_p0_wr_addr[7:4];
  assign dc2sbuf_p1_rd_bsel = dc2sbuf_p1_rd_addr[7:4];
  assign dc2sbuf_p1_rd_data = sbuf_p1_rdat_d2;
  assign dc2sbuf_p1_rd_esel = dc2sbuf_p1_rd_addr[3:0];
  assign dc2sbuf_p1_wr_bsel = dc2sbuf_p1_wr_addr[7:4];
  assign img2sbuf_p0_rd_bsel = img2sbuf_p0_rd_addr[7:4];
  assign img2sbuf_p0_rd_data = sbuf_p0_rdat_d2;
  assign img2sbuf_p0_rd_esel = img2sbuf_p0_rd_addr[3:0];
  assign img2sbuf_p0_wr_bsel = img2sbuf_p0_wr_addr[7:4];
  assign img2sbuf_p1_rd_bsel = img2sbuf_p1_rd_addr[7:4];
  assign img2sbuf_p1_rd_data = sbuf_p1_rdat_d2;
  assign img2sbuf_p1_rd_esel = img2sbuf_p1_rd_addr[3:0];
  assign img2sbuf_p1_wr_bsel = img2sbuf_p1_wr_addr[7:4];
  assign wg2sbuf_p0_rd_bsel = wg2sbuf_p0_rd_addr[7:6];
  assign wg2sbuf_p0_rd_data = sbuf_p0_rdat_d2;
  assign wg2sbuf_p0_rd_esel = wg2sbuf_p0_rd_addr[5:2];
  assign wg2sbuf_p0_rd_sel_01 = wg2sbuf_p0_rd_sel_00;
  assign wg2sbuf_p0_rd_sel_02 = wg2sbuf_p0_rd_sel_00;
  assign wg2sbuf_p0_rd_sel_03 = wg2sbuf_p0_rd_sel_00;
  assign wg2sbuf_p0_rd_sel_05 = wg2sbuf_p0_rd_sel_04;
  assign wg2sbuf_p0_rd_sel_06 = wg2sbuf_p0_rd_sel_04;
  assign wg2sbuf_p0_rd_sel_07 = wg2sbuf_p0_rd_sel_04;
  assign wg2sbuf_p0_rd_sel_09 = wg2sbuf_p0_rd_sel_08;
  assign wg2sbuf_p0_rd_sel_10 = wg2sbuf_p0_rd_sel_08;
  assign wg2sbuf_p0_rd_sel_11 = wg2sbuf_p0_rd_sel_08;
  assign wg2sbuf_p0_rd_sel_13 = wg2sbuf_p0_rd_sel_12;
  assign wg2sbuf_p0_rd_sel_14 = wg2sbuf_p0_rd_sel_12;
  assign wg2sbuf_p0_rd_sel_15 = wg2sbuf_p0_rd_sel_12;
  assign wg2sbuf_p0_wr_bsel = wg2sbuf_p0_wr_addr[7:4];
  assign wg2sbuf_p1_rd_bsel = wg2sbuf_p1_rd_addr[7:6];
  assign wg2sbuf_p1_rd_data = sbuf_p1_rdat_d2;
  assign wg2sbuf_p1_rd_esel = wg2sbuf_p1_rd_addr[5:2];
  assign wg2sbuf_p1_rd_sel_01 = wg2sbuf_p1_rd_sel_00;
  assign wg2sbuf_p1_rd_sel_02 = wg2sbuf_p1_rd_sel_00;
  assign wg2sbuf_p1_rd_sel_03 = wg2sbuf_p1_rd_sel_00;
  assign wg2sbuf_p1_rd_sel_05 = wg2sbuf_p1_rd_sel_04;
  assign wg2sbuf_p1_rd_sel_06 = wg2sbuf_p1_rd_sel_04;
  assign wg2sbuf_p1_rd_sel_07 = wg2sbuf_p1_rd_sel_04;
  assign wg2sbuf_p1_rd_sel_09 = wg2sbuf_p1_rd_sel_08;
  assign wg2sbuf_p1_rd_sel_10 = wg2sbuf_p1_rd_sel_08;
  assign wg2sbuf_p1_rd_sel_11 = wg2sbuf_p1_rd_sel_08;
  assign wg2sbuf_p1_rd_sel_13 = wg2sbuf_p1_rd_sel_12;
  assign wg2sbuf_p1_rd_sel_14 = wg2sbuf_p1_rd_sel_12;
  assign wg2sbuf_p1_rd_sel_15 = wg2sbuf_p1_rd_sel_12;
  assign wg2sbuf_p1_wr_bsel = wg2sbuf_p1_wr_addr[7:4];
endmodule
