module \$paramod\CDP_OCVT_mgc_in_wire_v1\rscid=4\width=6 (d, z);
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:78" *)
  output [5:0] d;
  (* src = "./vmod/vlibs/HLS_cdp_ocvt.v:79" *)
  input [5:0] z;
  assign d = z;
endmodule
