module \$paramod\SDP_X_mgc_in_wire_v1\rscid=28\width=6 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:109" *)
  output [5:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:110" *)
  input [5:0] z;
  assign d = z;
endmodule
