module FP16_TO_FP17_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp16_to_fp17.v:179" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp16_to_fp17.v:180" *)
  output outsig;
  assign outsig = in_0;
endmodule
