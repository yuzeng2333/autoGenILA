module FP32_ADD_chn_o_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp32_add.v:341" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp32_add.v:342" *)
  output outsig;
  assign outsig = in_0;
endmodule
