module SDP_C_leading_sign_17_0(mantissa, rtn);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:282" *)
  wire _000_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *)
  wire _001_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:290" *)
  wire _002_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:291" *)
  wire _003_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *)
  wire _004_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *)
  wire _005_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _006_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _007_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _008_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _009_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _010_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _011_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *)
  wire _012_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:274" *)
  wire _013_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:281" *)
  wire _014_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:270" *)
  wire _015_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:271" *)
  wire _016_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:272" *)
  wire _017_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:276" *)
  wire _018_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:277" *)
  wire _019_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:278" *)
  wire _020_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *)
  wire _021_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _022_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _023_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _024_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:284" *)
  wire _025_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *)
  wire _026_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *)
  wire _027_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:291" *)
  wire _028_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *)
  wire _029_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *)
  wire _030_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *)
  wire _031_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *)
  wire _032_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _033_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _034_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _035_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _036_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _037_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _038_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _039_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _040_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _041_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *)
  wire _042_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *)
  wire _043_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *)
  wire _044_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:287" *)
  wire _045_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:290" *)
  wire _046_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:291" *)
  wire _047_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *)
  wire _048_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *)
  wire _049_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _050_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *)
  wire _051_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *)
  wire _052_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *)
  wire _053_;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:267" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:266" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:268" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:265" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:258" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:254" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:259" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:255" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:260" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:256" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:257" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:253" *)
  wire IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:261" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:262" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:263" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:264" *)
  wire c_h_1_7;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:250" *)
  input [16:0] mantissa;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:251" *)
  output [4:0] rtn;
  assign c_h_1_2 = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:273" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3 = _013_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:275" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:279" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:280" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _014_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:282" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:282" *) c_h_1_5;
  assign c_h_1_7 = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:283" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl = c_h_1_6 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:284" *) _025_;
  assign _001_ = c_h_1_2 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *) _044_;
  assign _002_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:290" *) _046_;
  assign _003_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:291" *) _047_;
  assign _004_ = _028_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *) c_h_1_6;
  assign _005_ = _002_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *) _029_;
  assign _006_ = _050_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) c_h_1_2;
  assign _007_ = _032_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _034_;
  assign _008_ = _052_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) c_h_1_5;
  assign _009_ = _036_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _038_;
  assign _010_ = _039_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) c_h_1_6;
  assign _011_ = _007_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _040_;
  assign _012_ = _043_ & (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *) c_h_1_7;
  assign _013_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:274" *) mantissa[10:9];
  assign _014_ = ! (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:281" *) mantissa[2:1];
  assign _015_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:270" *) mantissa[14:13];
  assign _016_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:271" *) mantissa[16:15];
  assign _017_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:272" *) mantissa[12:11];
  assign _018_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:276" *) mantissa[6:5];
  assign _019_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:277" *) mantissa[8:7];
  assign _020_ = | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:278" *) mantissa[4:3];
  assign _021_ = mantissa[15:14] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *) 1'b1;
  assign _022_ = mantissa[11:10] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) 1'b1;
  assign _023_ = mantissa[7:6] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) 1'b1;
  assign _024_ = mantissa[3:2] != (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) 1'b1;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:270" *) _015_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:271" *) _016_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:272" *) _017_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:276" *) _018_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:277" *) _019_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:278" *) _020_;
  assign _025_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:284" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_42_4_sdt_4;
  assign _026_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *) IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_18_3_sdt_3;
  assign _027_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *) _001_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:287" *) _045_;
  assign _028_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:291" *) _003_;
  assign _029_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *) _004_;
  assign _030_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *) _005_;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *) _048_;
  assign _031_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *) _021_;
  assign _032_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *) _049_;
  assign _033_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _022_;
  assign _034_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _006_;
  assign _035_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _023_;
  assign _036_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _051_;
  assign _037_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _024_;
  assign _038_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _008_;
  assign _039_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _009_;
  assign _040_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _010_;
  assign _041_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _011_;
  assign _042_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *) _053_;
  assign _043_ = ~ (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *) mantissa[0];
  assign _044_ = c_h_1_5 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:286" *) _026_;
  assign _045_ = _027_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:287" *) c_h_1_7;
  assign _046_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:290" *) _015_;
  assign _047_ = IntLeadZero_17U_leading_sign_17_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:291" *) _018_;
  assign _048_ = _030_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:292" *) c_h_1_7;
  assign _049_ = mantissa[16] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:294" *) _031_;
  assign _050_ = mantissa[12] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _033_;
  assign _051_ = mantissa[8] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:295" *) _035_;
  assign _052_ = mantissa[4] | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:296" *) _037_;
  assign _053_ = _041_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *) c_h_1_7;
  assign IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl = _042_ | (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:297" *) _012_;
  assign rtn = { c_h_1_7, IntLeadZero_17U_leading_sign_17_0_rtn_and_63_nl, IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_nl, IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_nor_10_nl, IntLeadZero_17U_leading_sign_17_0_rtn_IntLeadZero_17U_leading_sign_17_0_rtn_or_nl };
endmodule
