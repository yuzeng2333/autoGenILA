module one_round(clk, state_in, key, state_out);
  logic [7:0] _0000_;
  logic _0001_;
  logic _0002_;
  logic _0003_;
  logic _0004_;
  logic _0005_;
  logic _0006_;
  logic _0007_;
  logic _0008_;
  logic _0009_;
  logic _0010_;
  logic _0011_;
  logic _0012_;
  logic _0013_;
  logic _0014_;
  logic _0015_;
  logic _0016_;
  logic _0017_;
  logic _0018_;
  logic _0019_;
  logic _0020_;
  logic _0021_;
  logic _0022_;
  logic _0023_;
  logic _0024_;
  logic _0025_;
  logic _0026_;
  logic _0027_;
  logic _0028_;
  logic _0029_;
  logic _0030_;
  logic _0031_;
  logic _0032_;
  logic _0033_;
  logic _0034_;
  logic _0035_;
  logic _0036_;
  logic _0037_;
  logic _0038_;
  logic _0039_;
  logic _0040_;
  logic _0041_;
  logic _0042_;
  logic _0043_;
  logic _0044_;
  logic _0045_;
  logic _0046_;
  logic _0047_;
  logic _0048_;
  logic _0049_;
  logic _0050_;
  logic _0051_;
  logic _0052_;
  logic _0053_;
  logic _0054_;
  logic _0055_;
  logic _0056_;
  logic _0057_;
  logic _0058_;
  logic _0059_;
  logic _0060_;
  logic _0061_;
  logic _0062_;
  logic _0063_;
  logic _0064_;
  logic _0065_;
  logic _0066_;
  logic _0067_;
  logic _0068_;
  logic _0069_;
  logic _0070_;
  logic _0071_;
  logic _0072_;
  logic _0073_;
  logic _0074_;
  logic _0075_;
  logic _0076_;
  logic _0077_;
  logic _0078_;
  logic _0079_;
  logic _0080_;
  logic _0081_;
  logic _0082_;
  logic _0083_;
  logic _0084_;
  logic _0085_;
  logic _0086_;
  logic _0087_;
  logic _0088_;
  logic _0089_;
  logic _0090_;
  logic _0091_;
  logic _0092_;
  logic _0093_;
  logic _0094_;
  logic _0095_;
  logic _0096_;
  logic _0097_;
  logic _0098_;
  logic _0099_;
  logic _0100_;
  logic _0101_;
  logic _0102_;
  logic _0103_;
  logic _0104_;
  logic _0105_;
  logic _0106_;
  logic _0107_;
  logic _0108_;
  logic _0109_;
  logic _0110_;
  logic _0111_;
  logic _0112_;
  logic _0113_;
  logic _0114_;
  logic _0115_;
  logic _0116_;
  logic _0117_;
  logic _0118_;
  logic _0119_;
  logic _0120_;
  logic _0121_;
  logic _0122_;
  logic _0123_;
  logic _0124_;
  logic _0125_;
  logic _0126_;
  logic _0127_;
  logic _0128_;
  logic _0129_;
  logic _0130_;
  logic _0131_;
  logic _0132_;
  logic _0133_;
  logic _0134_;
  logic _0135_;
  logic _0136_;
  logic _0137_;
  logic _0138_;
  logic _0139_;
  logic _0140_;
  logic _0141_;
  logic _0142_;
  logic _0143_;
  logic _0144_;
  logic _0145_;
  logic _0146_;
  logic _0147_;
  logic _0148_;
  logic _0149_;
  logic _0150_;
  logic _0151_;
  logic _0152_;
  logic _0153_;
  logic _0154_;
  logic _0155_;
  logic _0156_;
  logic _0157_;
  logic _0158_;
  logic _0159_;
  logic _0160_;
  logic _0161_;
  logic _0162_;
  logic _0163_;
  logic _0164_;
  logic _0165_;
  logic _0166_;
  logic _0167_;
  logic _0168_;
  logic _0169_;
  logic _0170_;
  logic _0171_;
  logic _0172_;
  logic _0173_;
  logic _0174_;
  logic _0175_;
  logic _0176_;
  logic _0177_;
  logic _0178_;
  logic _0179_;
  logic _0180_;
  logic _0181_;
  logic _0182_;
  logic _0183_;
  logic _0184_;
  logic _0185_;
  logic _0186_;
  logic _0187_;
  logic _0188_;
  logic _0189_;
  logic _0190_;
  logic _0191_;
  logic _0192_;
  logic _0193_;
  logic _0194_;
  logic _0195_;
  logic _0196_;
  logic _0197_;
  logic _0198_;
  logic _0199_;
  logic _0200_;
  logic _0201_;
  logic _0202_;
  logic _0203_;
  logic _0204_;
  logic _0205_;
  logic _0206_;
  logic _0207_;
  logic _0208_;
  logic _0209_;
  logic _0210_;
  logic _0211_;
  logic _0212_;
  logic _0213_;
  logic _0214_;
  logic _0215_;
  logic _0216_;
  logic _0217_;
  logic _0218_;
  logic _0219_;
  logic _0220_;
  logic _0221_;
  logic _0222_;
  logic _0223_;
  logic _0224_;
  logic _0225_;
  logic _0226_;
  logic _0227_;
  logic _0228_;
  logic _0229_;
  logic _0230_;
  logic _0231_;
  logic _0232_;
  logic _0233_;
  logic _0234_;
  logic _0235_;
  logic _0236_;
  logic _0237_;
  logic _0238_;
  logic _0239_;
  logic _0240_;
  logic _0241_;
  logic _0242_;
  logic _0243_;
  logic _0244_;
  logic _0245_;
  logic _0246_;
  logic _0247_;
  logic _0248_;
  logic _0249_;
  logic _0250_;
  logic _0251_;
  logic _0252_;
  logic _0253_;
  logic _0254_;
  logic _0255_;
  logic _0256_;
  logic [7:0] _0257_;
  logic [7:0] _0258_;
  logic _0259_;
  logic _0260_;
  logic _0261_;
  logic _0262_;
  logic _0263_;
  logic _0264_;
  logic _0265_;
  logic _0266_;
  logic _0267_;
  logic _0268_;
  logic _0269_;
  logic _0270_;
  logic _0271_;
  logic _0272_;
  logic _0273_;
  logic _0274_;
  logic _0275_;
  logic _0276_;
  logic _0277_;
  logic _0278_;
  logic _0279_;
  logic _0280_;
  logic _0281_;
  logic _0282_;
  logic _0283_;
  logic _0284_;
  logic _0285_;
  logic _0286_;
  logic _0287_;
  logic _0288_;
  logic _0289_;
  logic _0290_;
  logic _0291_;
  logic _0292_;
  logic _0293_;
  logic _0294_;
  logic _0295_;
  logic _0296_;
  logic _0297_;
  logic _0298_;
  logic _0299_;
  logic _0300_;
  logic _0301_;
  logic _0302_;
  logic _0303_;
  logic _0304_;
  logic _0305_;
  logic _0306_;
  logic _0307_;
  logic _0308_;
  logic _0309_;
  logic _0310_;
  logic _0311_;
  logic _0312_;
  logic _0313_;
  logic _0314_;
  logic _0315_;
  logic _0316_;
  logic _0317_;
  logic _0318_;
  logic _0319_;
  logic _0320_;
  logic _0321_;
  logic _0322_;
  logic _0323_;
  logic _0324_;
  logic _0325_;
  logic _0326_;
  logic _0327_;
  logic _0328_;
  logic _0329_;
  logic _0330_;
  logic _0331_;
  logic _0332_;
  logic _0333_;
  logic _0334_;
  logic _0335_;
  logic _0336_;
  logic _0337_;
  logic _0338_;
  logic _0339_;
  logic _0340_;
  logic _0341_;
  logic _0342_;
  logic _0343_;
  logic _0344_;
  logic _0345_;
  logic _0346_;
  logic _0347_;
  logic _0348_;
  logic _0349_;
  logic _0350_;
  logic _0351_;
  logic _0352_;
  logic _0353_;
  logic _0354_;
  logic _0355_;
  logic _0356_;
  logic _0357_;
  logic _0358_;
  logic _0359_;
  logic _0360_;
  logic _0361_;
  logic _0362_;
  logic _0363_;
  logic _0364_;
  logic _0365_;
  logic _0366_;
  logic _0367_;
  logic _0368_;
  logic _0369_;
  logic _0370_;
  logic _0371_;
  logic _0372_;
  logic _0373_;
  logic _0374_;
  logic _0375_;
  logic _0376_;
  logic _0377_;
  logic _0378_;
  logic _0379_;
  logic _0380_;
  logic _0381_;
  logic _0382_;
  logic _0383_;
  logic _0384_;
  logic _0385_;
  logic _0386_;
  logic _0387_;
  logic _0388_;
  logic _0389_;
  logic _0390_;
  logic _0391_;
  logic _0392_;
  logic _0393_;
  logic _0394_;
  logic _0395_;
  logic _0396_;
  logic _0397_;
  logic _0398_;
  logic _0399_;
  logic _0400_;
  logic _0401_;
  logic _0402_;
  logic _0403_;
  logic _0404_;
  logic _0405_;
  logic _0406_;
  logic _0407_;
  logic _0408_;
  logic _0409_;
  logic _0410_;
  logic _0411_;
  logic _0412_;
  logic _0413_;
  logic _0414_;
  logic _0415_;
  logic _0416_;
  logic _0417_;
  logic _0418_;
  logic _0419_;
  logic _0420_;
  logic _0421_;
  logic _0422_;
  logic _0423_;
  logic _0424_;
  logic _0425_;
  logic _0426_;
  logic _0427_;
  logic _0428_;
  logic _0429_;
  logic _0430_;
  logic _0431_;
  logic _0432_;
  logic _0433_;
  logic _0434_;
  logic _0435_;
  logic _0436_;
  logic _0437_;
  logic _0438_;
  logic _0439_;
  logic _0440_;
  logic _0441_;
  logic _0442_;
  logic _0443_;
  logic _0444_;
  logic _0445_;
  logic _0446_;
  logic _0447_;
  logic _0448_;
  logic _0449_;
  logic _0450_;
  logic _0451_;
  logic _0452_;
  logic _0453_;
  logic _0454_;
  logic _0455_;
  logic _0456_;
  logic _0457_;
  logic _0458_;
  logic _0459_;
  logic _0460_;
  logic _0461_;
  logic _0462_;
  logic _0463_;
  logic _0464_;
  logic _0465_;
  logic _0466_;
  logic _0467_;
  logic _0468_;
  logic _0469_;
  logic _0470_;
  logic _0471_;
  logic _0472_;
  logic _0473_;
  logic _0474_;
  logic _0475_;
  logic _0476_;
  logic _0477_;
  logic _0478_;
  logic _0479_;
  logic _0480_;
  logic _0481_;
  logic _0482_;
  logic _0483_;
  logic _0484_;
  logic _0485_;
  logic _0486_;
  logic _0487_;
  logic _0488_;
  logic _0489_;
  logic _0490_;
  logic _0491_;
  logic _0492_;
  logic _0493_;
  logic _0494_;
  logic _0495_;
  logic _0496_;
  logic _0497_;
  logic _0498_;
  logic _0499_;
  logic _0500_;
  logic _0501_;
  logic _0502_;
  logic _0503_;
  logic _0504_;
  logic _0505_;
  logic _0506_;
  logic _0507_;
  logic _0508_;
  logic _0509_;
  logic _0510_;
  logic _0511_;
  logic _0512_;
  logic _0513_;
  logic _0514_;
  logic [7:0] _0515_;
  logic [7:0] _0516_;
  logic _0517_;
  logic _0518_;
  logic _0519_;
  logic _0520_;
  logic _0521_;
  logic _0522_;
  logic _0523_;
  logic _0524_;
  logic _0525_;
  logic _0526_;
  logic _0527_;
  logic _0528_;
  logic _0529_;
  logic _0530_;
  logic _0531_;
  logic _0532_;
  logic _0533_;
  logic _0534_;
  logic _0535_;
  logic _0536_;
  logic _0537_;
  logic _0538_;
  logic _0539_;
  logic _0540_;
  logic _0541_;
  logic _0542_;
  logic _0543_;
  logic _0544_;
  logic _0545_;
  logic _0546_;
  logic _0547_;
  logic _0548_;
  logic _0549_;
  logic _0550_;
  logic _0551_;
  logic _0552_;
  logic _0553_;
  logic _0554_;
  logic _0555_;
  logic _0556_;
  logic _0557_;
  logic _0558_;
  logic _0559_;
  logic _0560_;
  logic _0561_;
  logic _0562_;
  logic _0563_;
  logic _0564_;
  logic _0565_;
  logic _0566_;
  logic _0567_;
  logic _0568_;
  logic _0569_;
  logic _0570_;
  logic _0571_;
  logic _0572_;
  logic _0573_;
  logic _0574_;
  logic _0575_;
  logic _0576_;
  logic _0577_;
  logic _0578_;
  logic _0579_;
  logic _0580_;
  logic _0581_;
  logic _0582_;
  logic _0583_;
  logic _0584_;
  logic _0585_;
  logic _0586_;
  logic _0587_;
  logic _0588_;
  logic _0589_;
  logic _0590_;
  logic _0591_;
  logic _0592_;
  logic _0593_;
  logic _0594_;
  logic _0595_;
  logic _0596_;
  logic _0597_;
  logic _0598_;
  logic _0599_;
  logic _0600_;
  logic _0601_;
  logic _0602_;
  logic _0603_;
  logic _0604_;
  logic _0605_;
  logic _0606_;
  logic _0607_;
  logic _0608_;
  logic _0609_;
  logic _0610_;
  logic _0611_;
  logic _0612_;
  logic _0613_;
  logic _0614_;
  logic _0615_;
  logic _0616_;
  logic _0617_;
  logic _0618_;
  logic _0619_;
  logic _0620_;
  logic _0621_;
  logic _0622_;
  logic _0623_;
  logic _0624_;
  logic _0625_;
  logic _0626_;
  logic _0627_;
  logic _0628_;
  logic _0629_;
  logic _0630_;
  logic _0631_;
  logic _0632_;
  logic _0633_;
  logic _0634_;
  logic _0635_;
  logic _0636_;
  logic _0637_;
  logic _0638_;
  logic _0639_;
  logic _0640_;
  logic _0641_;
  logic _0642_;
  logic _0643_;
  logic _0644_;
  logic _0645_;
  logic _0646_;
  logic _0647_;
  logic _0648_;
  logic _0649_;
  logic _0650_;
  logic _0651_;
  logic _0652_;
  logic _0653_;
  logic _0654_;
  logic _0655_;
  logic _0656_;
  logic _0657_;
  logic _0658_;
  logic _0659_;
  logic _0660_;
  logic _0661_;
  logic _0662_;
  logic _0663_;
  logic _0664_;
  logic _0665_;
  logic _0666_;
  logic _0667_;
  logic _0668_;
  logic _0669_;
  logic _0670_;
  logic _0671_;
  logic _0672_;
  logic _0673_;
  logic _0674_;
  logic _0675_;
  logic _0676_;
  logic _0677_;
  logic _0678_;
  logic _0679_;
  logic _0680_;
  logic _0681_;
  logic _0682_;
  logic _0683_;
  logic _0684_;
  logic _0685_;
  logic _0686_;
  logic _0687_;
  logic _0688_;
  logic _0689_;
  logic _0690_;
  logic _0691_;
  logic _0692_;
  logic _0693_;
  logic _0694_;
  logic _0695_;
  logic _0696_;
  logic _0697_;
  logic _0698_;
  logic _0699_;
  logic _0700_;
  logic _0701_;
  logic _0702_;
  logic _0703_;
  logic _0704_;
  logic _0705_;
  logic _0706_;
  logic _0707_;
  logic _0708_;
  logic _0709_;
  logic _0710_;
  logic _0711_;
  logic _0712_;
  logic _0713_;
  logic _0714_;
  logic _0715_;
  logic _0716_;
  logic _0717_;
  logic _0718_;
  logic _0719_;
  logic _0720_;
  logic _0721_;
  logic _0722_;
  logic _0723_;
  logic _0724_;
  logic _0725_;
  logic _0726_;
  logic _0727_;
  logic _0728_;
  logic _0729_;
  logic _0730_;
  logic _0731_;
  logic _0732_;
  logic _0733_;
  logic _0734_;
  logic _0735_;
  logic _0736_;
  logic _0737_;
  logic _0738_;
  logic _0739_;
  logic _0740_;
  logic _0741_;
  logic _0742_;
  logic _0743_;
  logic _0744_;
  logic _0745_;
  logic _0746_;
  logic _0747_;
  logic _0748_;
  logic _0749_;
  logic _0750_;
  logic _0751_;
  logic _0752_;
  logic _0753_;
  logic _0754_;
  logic _0755_;
  logic _0756_;
  logic _0757_;
  logic _0758_;
  logic _0759_;
  logic _0760_;
  logic _0761_;
  logic _0762_;
  logic _0763_;
  logic _0764_;
  logic _0765_;
  logic _0766_;
  logic _0767_;
  logic _0768_;
  logic _0769_;
  logic _0770_;
  logic _0771_;
  logic _0772_;
  logic [7:0] _0773_;
  logic [7:0] _0774_;
  logic _0775_;
  logic _0776_;
  logic _0777_;
  logic _0778_;
  logic _0779_;
  logic _0780_;
  logic _0781_;
  logic _0782_;
  logic _0783_;
  logic _0784_;
  logic _0785_;
  logic _0786_;
  logic _0787_;
  logic _0788_;
  logic _0789_;
  logic _0790_;
  logic _0791_;
  logic _0792_;
  logic _0793_;
  logic _0794_;
  logic _0795_;
  logic _0796_;
  logic _0797_;
  logic _0798_;
  logic _0799_;
  logic _0800_;
  logic _0801_;
  logic _0802_;
  logic _0803_;
  logic _0804_;
  logic _0805_;
  logic _0806_;
  logic _0807_;
  logic _0808_;
  logic _0809_;
  logic _0810_;
  logic _0811_;
  logic _0812_;
  logic _0813_;
  logic _0814_;
  logic _0815_;
  logic _0816_;
  logic _0817_;
  logic _0818_;
  logic _0819_;
  logic _0820_;
  logic _0821_;
  logic _0822_;
  logic _0823_;
  logic _0824_;
  logic _0825_;
  logic _0826_;
  logic _0827_;
  logic _0828_;
  logic _0829_;
  logic _0830_;
  logic _0831_;
  logic _0832_;
  logic _0833_;
  logic _0834_;
  logic _0835_;
  logic _0836_;
  logic _0837_;
  logic _0838_;
  logic _0839_;
  logic _0840_;
  logic _0841_;
  logic _0842_;
  logic _0843_;
  logic _0844_;
  logic _0845_;
  logic _0846_;
  logic _0847_;
  logic _0848_;
  logic _0849_;
  logic _0850_;
  logic _0851_;
  logic _0852_;
  logic _0853_;
  logic _0854_;
  logic _0855_;
  logic _0856_;
  logic _0857_;
  logic _0858_;
  logic _0859_;
  logic _0860_;
  logic _0861_;
  logic _0862_;
  logic _0863_;
  logic _0864_;
  logic _0865_;
  logic _0866_;
  logic _0867_;
  logic _0868_;
  logic _0869_;
  logic _0870_;
  logic _0871_;
  logic _0872_;
  logic _0873_;
  logic _0874_;
  logic _0875_;
  logic _0876_;
  logic _0877_;
  logic _0878_;
  logic _0879_;
  logic _0880_;
  logic _0881_;
  logic _0882_;
  logic _0883_;
  logic _0884_;
  logic _0885_;
  logic _0886_;
  logic _0887_;
  logic _0888_;
  logic _0889_;
  logic _0890_;
  logic _0891_;
  logic _0892_;
  logic _0893_;
  logic _0894_;
  logic _0895_;
  logic _0896_;
  logic _0897_;
  logic _0898_;
  logic _0899_;
  logic _0900_;
  logic _0901_;
  logic _0902_;
  logic _0903_;
  logic _0904_;
  logic _0905_;
  logic _0906_;
  logic _0907_;
  logic _0908_;
  logic _0909_;
  logic _0910_;
  logic _0911_;
  logic _0912_;
  logic _0913_;
  logic _0914_;
  logic _0915_;
  logic _0916_;
  logic _0917_;
  logic _0918_;
  logic _0919_;
  logic _0920_;
  logic _0921_;
  logic _0922_;
  logic _0923_;
  logic _0924_;
  logic _0925_;
  logic _0926_;
  logic _0927_;
  logic _0928_;
  logic _0929_;
  logic _0930_;
  logic _0931_;
  logic _0932_;
  logic _0933_;
  logic _0934_;
  logic _0935_;
  logic _0936_;
  logic _0937_;
  logic _0938_;
  logic _0939_;
  logic _0940_;
  logic _0941_;
  logic _0942_;
  logic _0943_;
  logic _0944_;
  logic _0945_;
  logic _0946_;
  logic _0947_;
  logic _0948_;
  logic _0949_;
  logic _0950_;
  logic _0951_;
  logic _0952_;
  logic _0953_;
  logic _0954_;
  logic _0955_;
  logic _0956_;
  logic _0957_;
  logic _0958_;
  logic _0959_;
  logic _0960_;
  logic _0961_;
  logic _0962_;
  logic _0963_;
  logic _0964_;
  logic _0965_;
  logic _0966_;
  logic _0967_;
  logic _0968_;
  logic _0969_;
  logic _0970_;
  logic _0971_;
  logic _0972_;
  logic _0973_;
  logic _0974_;
  logic _0975_;
  logic _0976_;
  logic _0977_;
  logic _0978_;
  logic _0979_;
  logic _0980_;
  logic _0981_;
  logic _0982_;
  logic _0983_;
  logic _0984_;
  logic _0985_;
  logic _0986_;
  logic _0987_;
  logic _0988_;
  logic _0989_;
  logic _0990_;
  logic _0991_;
  logic _0992_;
  logic _0993_;
  logic _0994_;
  logic _0995_;
  logic _0996_;
  logic _0997_;
  logic _0998_;
  logic _0999_;
  logic _1000_;
  logic _1001_;
  logic _1002_;
  logic _1003_;
  logic _1004_;
  logic _1005_;
  logic _1006_;
  logic _1007_;
  logic _1008_;
  logic _1009_;
  logic _1010_;
  logic _1011_;
  logic _1012_;
  logic _1013_;
  logic _1014_;
  logic _1015_;
  logic _1016_;
  logic _1017_;
  logic _1018_;
  logic _1019_;
  logic _1020_;
  logic _1021_;
  logic _1022_;
  logic _1023_;
  logic _1024_;
  logic _1025_;
  logic _1026_;
  logic _1027_;
  logic _1028_;
  logic _1029_;
  logic _1030_;
  logic [7:0] _1031_;
  logic [7:0] _1032_;
  logic _1033_;
  logic _1034_;
  logic _1035_;
  logic _1036_;
  logic _1037_;
  logic _1038_;
  logic _1039_;
  logic _1040_;
  logic _1041_;
  logic _1042_;
  logic _1043_;
  logic _1044_;
  logic _1045_;
  logic _1046_;
  logic _1047_;
  logic _1048_;
  logic _1049_;
  logic _1050_;
  logic _1051_;
  logic _1052_;
  logic _1053_;
  logic _1054_;
  logic _1055_;
  logic _1056_;
  logic _1057_;
  logic _1058_;
  logic _1059_;
  logic _1060_;
  logic _1061_;
  logic _1062_;
  logic _1063_;
  logic _1064_;
  logic _1065_;
  logic _1066_;
  logic _1067_;
  logic _1068_;
  logic _1069_;
  logic _1070_;
  logic _1071_;
  logic _1072_;
  logic _1073_;
  logic _1074_;
  logic _1075_;
  logic _1076_;
  logic _1077_;
  logic _1078_;
  logic _1079_;
  logic _1080_;
  logic _1081_;
  logic _1082_;
  logic _1083_;
  logic _1084_;
  logic _1085_;
  logic _1086_;
  logic _1087_;
  logic _1088_;
  logic _1089_;
  logic _1090_;
  logic _1091_;
  logic _1092_;
  logic _1093_;
  logic _1094_;
  logic _1095_;
  logic _1096_;
  logic _1097_;
  logic _1098_;
  logic _1099_;
  logic _1100_;
  logic _1101_;
  logic _1102_;
  logic _1103_;
  logic _1104_;
  logic _1105_;
  logic _1106_;
  logic _1107_;
  logic _1108_;
  logic _1109_;
  logic _1110_;
  logic _1111_;
  logic _1112_;
  logic _1113_;
  logic _1114_;
  logic _1115_;
  logic _1116_;
  logic _1117_;
  logic _1118_;
  logic _1119_;
  logic _1120_;
  logic _1121_;
  logic _1122_;
  logic _1123_;
  logic _1124_;
  logic _1125_;
  logic _1126_;
  logic _1127_;
  logic _1128_;
  logic _1129_;
  logic _1130_;
  logic _1131_;
  logic _1132_;
  logic _1133_;
  logic _1134_;
  logic _1135_;
  logic _1136_;
  logic _1137_;
  logic _1138_;
  logic _1139_;
  logic _1140_;
  logic _1141_;
  logic _1142_;
  logic _1143_;
  logic _1144_;
  logic _1145_;
  logic _1146_;
  logic _1147_;
  logic _1148_;
  logic _1149_;
  logic _1150_;
  logic _1151_;
  logic _1152_;
  logic _1153_;
  logic _1154_;
  logic _1155_;
  logic _1156_;
  logic _1157_;
  logic _1158_;
  logic _1159_;
  logic _1160_;
  logic _1161_;
  logic _1162_;
  logic _1163_;
  logic _1164_;
  logic _1165_;
  logic _1166_;
  logic _1167_;
  logic _1168_;
  logic _1169_;
  logic _1170_;
  logic _1171_;
  logic _1172_;
  logic _1173_;
  logic _1174_;
  logic _1175_;
  logic _1176_;
  logic _1177_;
  logic _1178_;
  logic _1179_;
  logic _1180_;
  logic _1181_;
  logic _1182_;
  logic _1183_;
  logic _1184_;
  logic _1185_;
  logic _1186_;
  logic _1187_;
  logic _1188_;
  logic _1189_;
  logic _1190_;
  logic _1191_;
  logic _1192_;
  logic _1193_;
  logic _1194_;
  logic _1195_;
  logic _1196_;
  logic _1197_;
  logic _1198_;
  logic _1199_;
  logic _1200_;
  logic _1201_;
  logic _1202_;
  logic _1203_;
  logic _1204_;
  logic _1205_;
  logic _1206_;
  logic _1207_;
  logic _1208_;
  logic _1209_;
  logic _1210_;
  logic _1211_;
  logic _1212_;
  logic _1213_;
  logic _1214_;
  logic _1215_;
  logic _1216_;
  logic _1217_;
  logic _1218_;
  logic _1219_;
  logic _1220_;
  logic _1221_;
  logic _1222_;
  logic _1223_;
  logic _1224_;
  logic _1225_;
  logic _1226_;
  logic _1227_;
  logic _1228_;
  logic _1229_;
  logic _1230_;
  logic _1231_;
  logic _1232_;
  logic _1233_;
  logic _1234_;
  logic _1235_;
  logic _1236_;
  logic _1237_;
  logic _1238_;
  logic _1239_;
  logic _1240_;
  logic _1241_;
  logic _1242_;
  logic _1243_;
  logic _1244_;
  logic _1245_;
  logic _1246_;
  logic _1247_;
  logic _1248_;
  logic _1249_;
  logic _1250_;
  logic _1251_;
  logic _1252_;
  logic _1253_;
  logic _1254_;
  logic _1255_;
  logic _1256_;
  logic _1257_;
  logic _1258_;
  logic _1259_;
  logic _1260_;
  logic _1261_;
  logic _1262_;
  logic _1263_;
  logic _1264_;
  logic _1265_;
  logic _1266_;
  logic _1267_;
  logic _1268_;
  logic _1269_;
  logic _1270_;
  logic _1271_;
  logic _1272_;
  logic _1273_;
  logic _1274_;
  logic _1275_;
  logic _1276_;
  logic _1277_;
  logic _1278_;
  logic _1279_;
  logic _1280_;
  logic _1281_;
  logic _1282_;
  logic _1283_;
  logic _1284_;
  logic _1285_;
  logic _1286_;
  logic _1287_;
  logic _1288_;
  logic [7:0] _1289_;
  logic [7:0] _1290_;
  logic _1291_;
  logic _1292_;
  logic _1293_;
  logic _1294_;
  logic _1295_;
  logic _1296_;
  logic _1297_;
  logic _1298_;
  logic _1299_;
  logic _1300_;
  logic _1301_;
  logic _1302_;
  logic _1303_;
  logic _1304_;
  logic _1305_;
  logic _1306_;
  logic _1307_;
  logic _1308_;
  logic _1309_;
  logic _1310_;
  logic _1311_;
  logic _1312_;
  logic _1313_;
  logic _1314_;
  logic _1315_;
  logic _1316_;
  logic _1317_;
  logic _1318_;
  logic _1319_;
  logic _1320_;
  logic _1321_;
  logic _1322_;
  logic _1323_;
  logic _1324_;
  logic _1325_;
  logic _1326_;
  logic _1327_;
  logic _1328_;
  logic _1329_;
  logic _1330_;
  logic _1331_;
  logic _1332_;
  logic _1333_;
  logic _1334_;
  logic _1335_;
  logic _1336_;
  logic _1337_;
  logic _1338_;
  logic _1339_;
  logic _1340_;
  logic _1341_;
  logic _1342_;
  logic _1343_;
  logic _1344_;
  logic _1345_;
  logic _1346_;
  logic _1347_;
  logic _1348_;
  logic _1349_;
  logic _1350_;
  logic _1351_;
  logic _1352_;
  logic _1353_;
  logic _1354_;
  logic _1355_;
  logic _1356_;
  logic _1357_;
  logic _1358_;
  logic _1359_;
  logic _1360_;
  logic _1361_;
  logic _1362_;
  logic _1363_;
  logic _1364_;
  logic _1365_;
  logic _1366_;
  logic _1367_;
  logic _1368_;
  logic _1369_;
  logic _1370_;
  logic _1371_;
  logic _1372_;
  logic _1373_;
  logic _1374_;
  logic _1375_;
  logic _1376_;
  logic _1377_;
  logic _1378_;
  logic _1379_;
  logic _1380_;
  logic _1381_;
  logic _1382_;
  logic _1383_;
  logic _1384_;
  logic _1385_;
  logic _1386_;
  logic _1387_;
  logic _1388_;
  logic _1389_;
  logic _1390_;
  logic _1391_;
  logic _1392_;
  logic _1393_;
  logic _1394_;
  logic _1395_;
  logic _1396_;
  logic _1397_;
  logic _1398_;
  logic _1399_;
  logic _1400_;
  logic _1401_;
  logic _1402_;
  logic _1403_;
  logic _1404_;
  logic _1405_;
  logic _1406_;
  logic _1407_;
  logic _1408_;
  logic _1409_;
  logic _1410_;
  logic _1411_;
  logic _1412_;
  logic _1413_;
  logic _1414_;
  logic _1415_;
  logic _1416_;
  logic _1417_;
  logic _1418_;
  logic _1419_;
  logic _1420_;
  logic _1421_;
  logic _1422_;
  logic _1423_;
  logic _1424_;
  logic _1425_;
  logic _1426_;
  logic _1427_;
  logic _1428_;
  logic _1429_;
  logic _1430_;
  logic _1431_;
  logic _1432_;
  logic _1433_;
  logic _1434_;
  logic _1435_;
  logic _1436_;
  logic _1437_;
  logic _1438_;
  logic _1439_;
  logic _1440_;
  logic _1441_;
  logic _1442_;
  logic _1443_;
  logic _1444_;
  logic _1445_;
  logic _1446_;
  logic _1447_;
  logic _1448_;
  logic _1449_;
  logic _1450_;
  logic _1451_;
  logic _1452_;
  logic _1453_;
  logic _1454_;
  logic _1455_;
  logic _1456_;
  logic _1457_;
  logic _1458_;
  logic _1459_;
  logic _1460_;
  logic _1461_;
  logic _1462_;
  logic _1463_;
  logic _1464_;
  logic _1465_;
  logic _1466_;
  logic _1467_;
  logic _1468_;
  logic _1469_;
  logic _1470_;
  logic _1471_;
  logic _1472_;
  logic _1473_;
  logic _1474_;
  logic _1475_;
  logic _1476_;
  logic _1477_;
  logic _1478_;
  logic _1479_;
  logic _1480_;
  logic _1481_;
  logic _1482_;
  logic _1483_;
  logic _1484_;
  logic _1485_;
  logic _1486_;
  logic _1487_;
  logic _1488_;
  logic _1489_;
  logic _1490_;
  logic _1491_;
  logic _1492_;
  logic _1493_;
  logic _1494_;
  logic _1495_;
  logic _1496_;
  logic _1497_;
  logic _1498_;
  logic _1499_;
  logic _1500_;
  logic _1501_;
  logic _1502_;
  logic _1503_;
  logic _1504_;
  logic _1505_;
  logic _1506_;
  logic _1507_;
  logic _1508_;
  logic _1509_;
  logic _1510_;
  logic _1511_;
  logic _1512_;
  logic _1513_;
  logic _1514_;
  logic _1515_;
  logic _1516_;
  logic _1517_;
  logic _1518_;
  logic _1519_;
  logic _1520_;
  logic _1521_;
  logic _1522_;
  logic _1523_;
  logic _1524_;
  logic _1525_;
  logic _1526_;
  logic _1527_;
  logic _1528_;
  logic _1529_;
  logic _1530_;
  logic _1531_;
  logic _1532_;
  logic _1533_;
  logic _1534_;
  logic _1535_;
  logic _1536_;
  logic _1537_;
  logic _1538_;
  logic _1539_;
  logic _1540_;
  logic _1541_;
  logic _1542_;
  logic _1543_;
  logic _1544_;
  logic _1545_;
  logic _1546_;
  logic [7:0] _1547_;
  logic [7:0] _1548_;
  logic _1549_;
  logic _1550_;
  logic _1551_;
  logic _1552_;
  logic _1553_;
  logic _1554_;
  logic _1555_;
  logic _1556_;
  logic _1557_;
  logic _1558_;
  logic _1559_;
  logic _1560_;
  logic _1561_;
  logic _1562_;
  logic _1563_;
  logic _1564_;
  logic _1565_;
  logic _1566_;
  logic _1567_;
  logic _1568_;
  logic _1569_;
  logic _1570_;
  logic _1571_;
  logic _1572_;
  logic _1573_;
  logic _1574_;
  logic _1575_;
  logic _1576_;
  logic _1577_;
  logic _1578_;
  logic _1579_;
  logic _1580_;
  logic _1581_;
  logic _1582_;
  logic _1583_;
  logic _1584_;
  logic _1585_;
  logic _1586_;
  logic _1587_;
  logic _1588_;
  logic _1589_;
  logic _1590_;
  logic _1591_;
  logic _1592_;
  logic _1593_;
  logic _1594_;
  logic _1595_;
  logic _1596_;
  logic _1597_;
  logic _1598_;
  logic _1599_;
  logic _1600_;
  logic _1601_;
  logic _1602_;
  logic _1603_;
  logic _1604_;
  logic _1605_;
  logic _1606_;
  logic _1607_;
  logic _1608_;
  logic _1609_;
  logic _1610_;
  logic _1611_;
  logic _1612_;
  logic _1613_;
  logic _1614_;
  logic _1615_;
  logic _1616_;
  logic _1617_;
  logic _1618_;
  logic _1619_;
  logic _1620_;
  logic _1621_;
  logic _1622_;
  logic _1623_;
  logic _1624_;
  logic _1625_;
  logic _1626_;
  logic _1627_;
  logic _1628_;
  logic _1629_;
  logic _1630_;
  logic _1631_;
  logic _1632_;
  logic _1633_;
  logic _1634_;
  logic _1635_;
  logic _1636_;
  logic _1637_;
  logic _1638_;
  logic _1639_;
  logic _1640_;
  logic _1641_;
  logic _1642_;
  logic _1643_;
  logic _1644_;
  logic _1645_;
  logic _1646_;
  logic _1647_;
  logic _1648_;
  logic _1649_;
  logic _1650_;
  logic _1651_;
  logic _1652_;
  logic _1653_;
  logic _1654_;
  logic _1655_;
  logic _1656_;
  logic _1657_;
  logic _1658_;
  logic _1659_;
  logic _1660_;
  logic _1661_;
  logic _1662_;
  logic _1663_;
  logic _1664_;
  logic _1665_;
  logic _1666_;
  logic _1667_;
  logic _1668_;
  logic _1669_;
  logic _1670_;
  logic _1671_;
  logic _1672_;
  logic _1673_;
  logic _1674_;
  logic _1675_;
  logic _1676_;
  logic _1677_;
  logic _1678_;
  logic _1679_;
  logic _1680_;
  logic _1681_;
  logic _1682_;
  logic _1683_;
  logic _1684_;
  logic _1685_;
  logic _1686_;
  logic _1687_;
  logic _1688_;
  logic _1689_;
  logic _1690_;
  logic _1691_;
  logic _1692_;
  logic _1693_;
  logic _1694_;
  logic _1695_;
  logic _1696_;
  logic _1697_;
  logic _1698_;
  logic _1699_;
  logic _1700_;
  logic _1701_;
  logic _1702_;
  logic _1703_;
  logic _1704_;
  logic _1705_;
  logic _1706_;
  logic _1707_;
  logic _1708_;
  logic _1709_;
  logic _1710_;
  logic _1711_;
  logic _1712_;
  logic _1713_;
  logic _1714_;
  logic _1715_;
  logic _1716_;
  logic _1717_;
  logic _1718_;
  logic _1719_;
  logic _1720_;
  logic _1721_;
  logic _1722_;
  logic _1723_;
  logic _1724_;
  logic _1725_;
  logic _1726_;
  logic _1727_;
  logic _1728_;
  logic _1729_;
  logic _1730_;
  logic _1731_;
  logic _1732_;
  logic _1733_;
  logic _1734_;
  logic _1735_;
  logic _1736_;
  logic _1737_;
  logic _1738_;
  logic _1739_;
  logic _1740_;
  logic _1741_;
  logic _1742_;
  logic _1743_;
  logic _1744_;
  logic _1745_;
  logic _1746_;
  logic _1747_;
  logic _1748_;
  logic _1749_;
  logic _1750_;
  logic _1751_;
  logic _1752_;
  logic _1753_;
  logic _1754_;
  logic _1755_;
  logic _1756_;
  logic _1757_;
  logic _1758_;
  logic _1759_;
  logic _1760_;
  logic _1761_;
  logic _1762_;
  logic _1763_;
  logic _1764_;
  logic _1765_;
  logic _1766_;
  logic _1767_;
  logic _1768_;
  logic _1769_;
  logic _1770_;
  logic _1771_;
  logic _1772_;
  logic _1773_;
  logic _1774_;
  logic _1775_;
  logic _1776_;
  logic _1777_;
  logic _1778_;
  logic _1779_;
  logic _1780_;
  logic _1781_;
  logic _1782_;
  logic _1783_;
  logic _1784_;
  logic _1785_;
  logic _1786_;
  logic _1787_;
  logic _1788_;
  logic _1789_;
  logic _1790_;
  logic _1791_;
  logic _1792_;
  logic _1793_;
  logic _1794_;
  logic _1795_;
  logic _1796_;
  logic _1797_;
  logic _1798_;
  logic _1799_;
  logic _1800_;
  logic _1801_;
  logic _1802_;
  logic _1803_;
  logic _1804_;
  logic [7:0] _1805_;
  logic [7:0] _1806_;
  logic _1807_;
  logic _1808_;
  logic _1809_;
  logic _1810_;
  logic _1811_;
  logic _1812_;
  logic _1813_;
  logic _1814_;
  logic _1815_;
  logic _1816_;
  logic _1817_;
  logic _1818_;
  logic _1819_;
  logic _1820_;
  logic _1821_;
  logic _1822_;
  logic _1823_;
  logic _1824_;
  logic _1825_;
  logic _1826_;
  logic _1827_;
  logic _1828_;
  logic _1829_;
  logic _1830_;
  logic _1831_;
  logic _1832_;
  logic _1833_;
  logic _1834_;
  logic _1835_;
  logic _1836_;
  logic _1837_;
  logic _1838_;
  logic _1839_;
  logic _1840_;
  logic _1841_;
  logic _1842_;
  logic _1843_;
  logic _1844_;
  logic _1845_;
  logic _1846_;
  logic _1847_;
  logic _1848_;
  logic _1849_;
  logic _1850_;
  logic _1851_;
  logic _1852_;
  logic _1853_;
  logic _1854_;
  logic _1855_;
  logic _1856_;
  logic _1857_;
  logic _1858_;
  logic _1859_;
  logic _1860_;
  logic _1861_;
  logic _1862_;
  logic _1863_;
  logic _1864_;
  logic _1865_;
  logic _1866_;
  logic _1867_;
  logic _1868_;
  logic _1869_;
  logic _1870_;
  logic _1871_;
  logic _1872_;
  logic _1873_;
  logic _1874_;
  logic _1875_;
  logic _1876_;
  logic _1877_;
  logic _1878_;
  logic _1879_;
  logic _1880_;
  logic _1881_;
  logic _1882_;
  logic _1883_;
  logic _1884_;
  logic _1885_;
  logic _1886_;
  logic _1887_;
  logic _1888_;
  logic _1889_;
  logic _1890_;
  logic _1891_;
  logic _1892_;
  logic _1893_;
  logic _1894_;
  logic _1895_;
  logic _1896_;
  logic _1897_;
  logic _1898_;
  logic _1899_;
  logic _1900_;
  logic _1901_;
  logic _1902_;
  logic _1903_;
  logic _1904_;
  logic _1905_;
  logic _1906_;
  logic _1907_;
  logic _1908_;
  logic _1909_;
  logic _1910_;
  logic _1911_;
  logic _1912_;
  logic _1913_;
  logic _1914_;
  logic _1915_;
  logic _1916_;
  logic _1917_;
  logic _1918_;
  logic _1919_;
  logic _1920_;
  logic _1921_;
  logic _1922_;
  logic _1923_;
  logic _1924_;
  logic _1925_;
  logic _1926_;
  logic _1927_;
  logic _1928_;
  logic _1929_;
  logic _1930_;
  logic _1931_;
  logic _1932_;
  logic _1933_;
  logic _1934_;
  logic _1935_;
  logic _1936_;
  logic _1937_;
  logic _1938_;
  logic _1939_;
  logic _1940_;
  logic _1941_;
  logic _1942_;
  logic _1943_;
  logic _1944_;
  logic _1945_;
  logic _1946_;
  logic _1947_;
  logic _1948_;
  logic _1949_;
  logic _1950_;
  logic _1951_;
  logic _1952_;
  logic _1953_;
  logic _1954_;
  logic _1955_;
  logic _1956_;
  logic _1957_;
  logic _1958_;
  logic _1959_;
  logic _1960_;
  logic _1961_;
  logic _1962_;
  logic _1963_;
  logic _1964_;
  logic _1965_;
  logic _1966_;
  logic _1967_;
  logic _1968_;
  logic _1969_;
  logic _1970_;
  logic _1971_;
  logic _1972_;
  logic _1973_;
  logic _1974_;
  logic _1975_;
  logic _1976_;
  logic _1977_;
  logic _1978_;
  logic _1979_;
  logic _1980_;
  logic _1981_;
  logic _1982_;
  logic _1983_;
  logic _1984_;
  logic _1985_;
  logic _1986_;
  logic _1987_;
  logic _1988_;
  logic _1989_;
  logic _1990_;
  logic _1991_;
  logic _1992_;
  logic _1993_;
  logic _1994_;
  logic _1995_;
  logic _1996_;
  logic _1997_;
  logic _1998_;
  logic _1999_;
  logic _2000_;
  logic _2001_;
  logic _2002_;
  logic _2003_;
  logic _2004_;
  logic _2005_;
  logic _2006_;
  logic _2007_;
  logic _2008_;
  logic _2009_;
  logic _2010_;
  logic _2011_;
  logic _2012_;
  logic _2013_;
  logic _2014_;
  logic _2015_;
  logic _2016_;
  logic _2017_;
  logic _2018_;
  logic _2019_;
  logic _2020_;
  logic _2021_;
  logic _2022_;
  logic _2023_;
  logic _2024_;
  logic _2025_;
  logic _2026_;
  logic _2027_;
  logic _2028_;
  logic _2029_;
  logic _2030_;
  logic _2031_;
  logic _2032_;
  logic _2033_;
  logic _2034_;
  logic _2035_;
  logic _2036_;
  logic _2037_;
  logic _2038_;
  logic _2039_;
  logic _2040_;
  logic _2041_;
  logic _2042_;
  logic _2043_;
  logic _2044_;
  logic _2045_;
  logic _2046_;
  logic _2047_;
  logic _2048_;
  logic _2049_;
  logic _2050_;
  logic _2051_;
  logic _2052_;
  logic _2053_;
  logic _2054_;
  logic _2055_;
  logic _2056_;
  logic _2057_;
  logic _2058_;
  logic _2059_;
  logic _2060_;
  logic _2061_;
  logic _2062_;
  logic [7:0] _2063_;
  logic [7:0] _2064_;
  logic _2065_;
  logic _2066_;
  logic _2067_;
  logic _2068_;
  logic _2069_;
  logic _2070_;
  logic _2071_;
  logic _2072_;
  logic _2073_;
  logic _2074_;
  logic _2075_;
  logic _2076_;
  logic _2077_;
  logic _2078_;
  logic _2079_;
  logic _2080_;
  logic _2081_;
  logic _2082_;
  logic _2083_;
  logic _2084_;
  logic _2085_;
  logic _2086_;
  logic _2087_;
  logic _2088_;
  logic _2089_;
  logic _2090_;
  logic _2091_;
  logic _2092_;
  logic _2093_;
  logic _2094_;
  logic _2095_;
  logic _2096_;
  logic _2097_;
  logic _2098_;
  logic _2099_;
  logic _2100_;
  logic _2101_;
  logic _2102_;
  logic _2103_;
  logic _2104_;
  logic _2105_;
  logic _2106_;
  logic _2107_;
  logic _2108_;
  logic _2109_;
  logic _2110_;
  logic _2111_;
  logic _2112_;
  logic _2113_;
  logic _2114_;
  logic _2115_;
  logic _2116_;
  logic _2117_;
  logic _2118_;
  logic _2119_;
  logic _2120_;
  logic _2121_;
  logic _2122_;
  logic _2123_;
  logic _2124_;
  logic _2125_;
  logic _2126_;
  logic _2127_;
  logic _2128_;
  logic _2129_;
  logic _2130_;
  logic _2131_;
  logic _2132_;
  logic _2133_;
  logic _2134_;
  logic _2135_;
  logic _2136_;
  logic _2137_;
  logic _2138_;
  logic _2139_;
  logic _2140_;
  logic _2141_;
  logic _2142_;
  logic _2143_;
  logic _2144_;
  logic _2145_;
  logic _2146_;
  logic _2147_;
  logic _2148_;
  logic _2149_;
  logic _2150_;
  logic _2151_;
  logic _2152_;
  logic _2153_;
  logic _2154_;
  logic _2155_;
  logic _2156_;
  logic _2157_;
  logic _2158_;
  logic _2159_;
  logic _2160_;
  logic _2161_;
  logic _2162_;
  logic _2163_;
  logic _2164_;
  logic _2165_;
  logic _2166_;
  logic _2167_;
  logic _2168_;
  logic _2169_;
  logic _2170_;
  logic _2171_;
  logic _2172_;
  logic _2173_;
  logic _2174_;
  logic _2175_;
  logic _2176_;
  logic _2177_;
  logic _2178_;
  logic _2179_;
  logic _2180_;
  logic _2181_;
  logic _2182_;
  logic _2183_;
  logic _2184_;
  logic _2185_;
  logic _2186_;
  logic _2187_;
  logic _2188_;
  logic _2189_;
  logic _2190_;
  logic _2191_;
  logic _2192_;
  logic _2193_;
  logic _2194_;
  logic _2195_;
  logic _2196_;
  logic _2197_;
  logic _2198_;
  logic _2199_;
  logic _2200_;
  logic _2201_;
  logic _2202_;
  logic _2203_;
  logic _2204_;
  logic _2205_;
  logic _2206_;
  logic _2207_;
  logic _2208_;
  logic _2209_;
  logic _2210_;
  logic _2211_;
  logic _2212_;
  logic _2213_;
  logic _2214_;
  logic _2215_;
  logic _2216_;
  logic _2217_;
  logic _2218_;
  logic _2219_;
  logic _2220_;
  logic _2221_;
  logic _2222_;
  logic _2223_;
  logic _2224_;
  logic _2225_;
  logic _2226_;
  logic _2227_;
  logic _2228_;
  logic _2229_;
  logic _2230_;
  logic _2231_;
  logic _2232_;
  logic _2233_;
  logic _2234_;
  logic _2235_;
  logic _2236_;
  logic _2237_;
  logic _2238_;
  logic _2239_;
  logic _2240_;
  logic _2241_;
  logic _2242_;
  logic _2243_;
  logic _2244_;
  logic _2245_;
  logic _2246_;
  logic _2247_;
  logic _2248_;
  logic _2249_;
  logic _2250_;
  logic _2251_;
  logic _2252_;
  logic _2253_;
  logic _2254_;
  logic _2255_;
  logic _2256_;
  logic _2257_;
  logic _2258_;
  logic _2259_;
  logic _2260_;
  logic _2261_;
  logic _2262_;
  logic _2263_;
  logic _2264_;
  logic _2265_;
  logic _2266_;
  logic _2267_;
  logic _2268_;
  logic _2269_;
  logic _2270_;
  logic _2271_;
  logic _2272_;
  logic _2273_;
  logic _2274_;
  logic _2275_;
  logic _2276_;
  logic _2277_;
  logic _2278_;
  logic _2279_;
  logic _2280_;
  logic _2281_;
  logic _2282_;
  logic _2283_;
  logic _2284_;
  logic _2285_;
  logic _2286_;
  logic _2287_;
  logic _2288_;
  logic _2289_;
  logic _2290_;
  logic _2291_;
  logic _2292_;
  logic _2293_;
  logic _2294_;
  logic _2295_;
  logic _2296_;
  logic _2297_;
  logic _2298_;
  logic _2299_;
  logic _2300_;
  logic _2301_;
  logic _2302_;
  logic _2303_;
  logic _2304_;
  logic _2305_;
  logic _2306_;
  logic _2307_;
  logic _2308_;
  logic _2309_;
  logic _2310_;
  logic _2311_;
  logic _2312_;
  logic _2313_;
  logic _2314_;
  logic _2315_;
  logic _2316_;
  logic _2317_;
  logic _2318_;
  logic _2319_;
  logic _2320_;
  logic [7:0] _2321_;
  logic [7:0] _2322_;
  logic _2323_;
  logic _2324_;
  logic _2325_;
  logic _2326_;
  logic _2327_;
  logic _2328_;
  logic _2329_;
  logic _2330_;
  logic _2331_;
  logic _2332_;
  logic _2333_;
  logic _2334_;
  logic _2335_;
  logic _2336_;
  logic _2337_;
  logic _2338_;
  logic _2339_;
  logic _2340_;
  logic _2341_;
  logic _2342_;
  logic _2343_;
  logic _2344_;
  logic _2345_;
  logic _2346_;
  logic _2347_;
  logic _2348_;
  logic _2349_;
  logic _2350_;
  logic _2351_;
  logic _2352_;
  logic _2353_;
  logic _2354_;
  logic _2355_;
  logic _2356_;
  logic _2357_;
  logic _2358_;
  logic _2359_;
  logic _2360_;
  logic _2361_;
  logic _2362_;
  logic _2363_;
  logic _2364_;
  logic _2365_;
  logic _2366_;
  logic _2367_;
  logic _2368_;
  logic _2369_;
  logic _2370_;
  logic _2371_;
  logic _2372_;
  logic _2373_;
  logic _2374_;
  logic _2375_;
  logic _2376_;
  logic _2377_;
  logic _2378_;
  logic _2379_;
  logic _2380_;
  logic _2381_;
  logic _2382_;
  logic _2383_;
  logic _2384_;
  logic _2385_;
  logic _2386_;
  logic _2387_;
  logic _2388_;
  logic _2389_;
  logic _2390_;
  logic _2391_;
  logic _2392_;
  logic _2393_;
  logic _2394_;
  logic _2395_;
  logic _2396_;
  logic _2397_;
  logic _2398_;
  logic _2399_;
  logic _2400_;
  logic _2401_;
  logic _2402_;
  logic _2403_;
  logic _2404_;
  logic _2405_;
  logic _2406_;
  logic _2407_;
  logic _2408_;
  logic _2409_;
  logic _2410_;
  logic _2411_;
  logic _2412_;
  logic _2413_;
  logic _2414_;
  logic _2415_;
  logic _2416_;
  logic _2417_;
  logic _2418_;
  logic _2419_;
  logic _2420_;
  logic _2421_;
  logic _2422_;
  logic _2423_;
  logic _2424_;
  logic _2425_;
  logic _2426_;
  logic _2427_;
  logic _2428_;
  logic _2429_;
  logic _2430_;
  logic _2431_;
  logic _2432_;
  logic _2433_;
  logic _2434_;
  logic _2435_;
  logic _2436_;
  logic _2437_;
  logic _2438_;
  logic _2439_;
  logic _2440_;
  logic _2441_;
  logic _2442_;
  logic _2443_;
  logic _2444_;
  logic _2445_;
  logic _2446_;
  logic _2447_;
  logic _2448_;
  logic _2449_;
  logic _2450_;
  logic _2451_;
  logic _2452_;
  logic _2453_;
  logic _2454_;
  logic _2455_;
  logic _2456_;
  logic _2457_;
  logic _2458_;
  logic _2459_;
  logic _2460_;
  logic _2461_;
  logic _2462_;
  logic _2463_;
  logic _2464_;
  logic _2465_;
  logic _2466_;
  logic _2467_;
  logic _2468_;
  logic _2469_;
  logic _2470_;
  logic _2471_;
  logic _2472_;
  logic _2473_;
  logic _2474_;
  logic _2475_;
  logic _2476_;
  logic _2477_;
  logic _2478_;
  logic _2479_;
  logic _2480_;
  logic _2481_;
  logic _2482_;
  logic _2483_;
  logic _2484_;
  logic _2485_;
  logic _2486_;
  logic _2487_;
  logic _2488_;
  logic _2489_;
  logic _2490_;
  logic _2491_;
  logic _2492_;
  logic _2493_;
  logic _2494_;
  logic _2495_;
  logic _2496_;
  logic _2497_;
  logic _2498_;
  logic _2499_;
  logic _2500_;
  logic _2501_;
  logic _2502_;
  logic _2503_;
  logic _2504_;
  logic _2505_;
  logic _2506_;
  logic _2507_;
  logic _2508_;
  logic _2509_;
  logic _2510_;
  logic _2511_;
  logic _2512_;
  logic _2513_;
  logic _2514_;
  logic _2515_;
  logic _2516_;
  logic _2517_;
  logic _2518_;
  logic _2519_;
  logic _2520_;
  logic _2521_;
  logic _2522_;
  logic _2523_;
  logic _2524_;
  logic _2525_;
  logic _2526_;
  logic _2527_;
  logic _2528_;
  logic _2529_;
  logic _2530_;
  logic _2531_;
  logic _2532_;
  logic _2533_;
  logic _2534_;
  logic _2535_;
  logic _2536_;
  logic _2537_;
  logic _2538_;
  logic _2539_;
  logic _2540_;
  logic _2541_;
  logic _2542_;
  logic _2543_;
  logic _2544_;
  logic _2545_;
  logic _2546_;
  logic _2547_;
  logic _2548_;
  logic _2549_;
  logic _2550_;
  logic _2551_;
  logic _2552_;
  logic _2553_;
  logic _2554_;
  logic _2555_;
  logic _2556_;
  logic _2557_;
  logic _2558_;
  logic _2559_;
  logic _2560_;
  logic _2561_;
  logic _2562_;
  logic _2563_;
  logic _2564_;
  logic _2565_;
  logic _2566_;
  logic _2567_;
  logic _2568_;
  logic _2569_;
  logic _2570_;
  logic _2571_;
  logic _2572_;
  logic _2573_;
  logic _2574_;
  logic _2575_;
  logic _2576_;
  logic _2577_;
  logic _2578_;
  logic [7:0] _2579_;
  logic [7:0] _2580_;
  logic _2581_;
  logic _2582_;
  logic _2583_;
  logic _2584_;
  logic _2585_;
  logic _2586_;
  logic _2587_;
  logic _2588_;
  logic _2589_;
  logic _2590_;
  logic _2591_;
  logic _2592_;
  logic _2593_;
  logic _2594_;
  logic _2595_;
  logic _2596_;
  logic _2597_;
  logic _2598_;
  logic _2599_;
  logic _2600_;
  logic _2601_;
  logic _2602_;
  logic _2603_;
  logic _2604_;
  logic _2605_;
  logic _2606_;
  logic _2607_;
  logic _2608_;
  logic _2609_;
  logic _2610_;
  logic _2611_;
  logic _2612_;
  logic _2613_;
  logic _2614_;
  logic _2615_;
  logic _2616_;
  logic _2617_;
  logic _2618_;
  logic _2619_;
  logic _2620_;
  logic _2621_;
  logic _2622_;
  logic _2623_;
  logic _2624_;
  logic _2625_;
  logic _2626_;
  logic _2627_;
  logic _2628_;
  logic _2629_;
  logic _2630_;
  logic _2631_;
  logic _2632_;
  logic _2633_;
  logic _2634_;
  logic _2635_;
  logic _2636_;
  logic _2637_;
  logic _2638_;
  logic _2639_;
  logic _2640_;
  logic _2641_;
  logic _2642_;
  logic _2643_;
  logic _2644_;
  logic _2645_;
  logic _2646_;
  logic _2647_;
  logic _2648_;
  logic _2649_;
  logic _2650_;
  logic _2651_;
  logic _2652_;
  logic _2653_;
  logic _2654_;
  logic _2655_;
  logic _2656_;
  logic _2657_;
  logic _2658_;
  logic _2659_;
  logic _2660_;
  logic _2661_;
  logic _2662_;
  logic _2663_;
  logic _2664_;
  logic _2665_;
  logic _2666_;
  logic _2667_;
  logic _2668_;
  logic _2669_;
  logic _2670_;
  logic _2671_;
  logic _2672_;
  logic _2673_;
  logic _2674_;
  logic _2675_;
  logic _2676_;
  logic _2677_;
  logic _2678_;
  logic _2679_;
  logic _2680_;
  logic _2681_;
  logic _2682_;
  logic _2683_;
  logic _2684_;
  logic _2685_;
  logic _2686_;
  logic _2687_;
  logic _2688_;
  logic _2689_;
  logic _2690_;
  logic _2691_;
  logic _2692_;
  logic _2693_;
  logic _2694_;
  logic _2695_;
  logic _2696_;
  logic _2697_;
  logic _2698_;
  logic _2699_;
  logic _2700_;
  logic _2701_;
  logic _2702_;
  logic _2703_;
  logic _2704_;
  logic _2705_;
  logic _2706_;
  logic _2707_;
  logic _2708_;
  logic _2709_;
  logic _2710_;
  logic _2711_;
  logic _2712_;
  logic _2713_;
  logic _2714_;
  logic _2715_;
  logic _2716_;
  logic _2717_;
  logic _2718_;
  logic _2719_;
  logic _2720_;
  logic _2721_;
  logic _2722_;
  logic _2723_;
  logic _2724_;
  logic _2725_;
  logic _2726_;
  logic _2727_;
  logic _2728_;
  logic _2729_;
  logic _2730_;
  logic _2731_;
  logic _2732_;
  logic _2733_;
  logic _2734_;
  logic _2735_;
  logic _2736_;
  logic _2737_;
  logic _2738_;
  logic _2739_;
  logic _2740_;
  logic _2741_;
  logic _2742_;
  logic _2743_;
  logic _2744_;
  logic _2745_;
  logic _2746_;
  logic _2747_;
  logic _2748_;
  logic _2749_;
  logic _2750_;
  logic _2751_;
  logic _2752_;
  logic _2753_;
  logic _2754_;
  logic _2755_;
  logic _2756_;
  logic _2757_;
  logic _2758_;
  logic _2759_;
  logic _2760_;
  logic _2761_;
  logic _2762_;
  logic _2763_;
  logic _2764_;
  logic _2765_;
  logic _2766_;
  logic _2767_;
  logic _2768_;
  logic _2769_;
  logic _2770_;
  logic _2771_;
  logic _2772_;
  logic _2773_;
  logic _2774_;
  logic _2775_;
  logic _2776_;
  logic _2777_;
  logic _2778_;
  logic _2779_;
  logic _2780_;
  logic _2781_;
  logic _2782_;
  logic _2783_;
  logic _2784_;
  logic _2785_;
  logic _2786_;
  logic _2787_;
  logic _2788_;
  logic _2789_;
  logic _2790_;
  logic _2791_;
  logic _2792_;
  logic _2793_;
  logic _2794_;
  logic _2795_;
  logic _2796_;
  logic _2797_;
  logic _2798_;
  logic _2799_;
  logic _2800_;
  logic _2801_;
  logic _2802_;
  logic _2803_;
  logic _2804_;
  logic _2805_;
  logic _2806_;
  logic _2807_;
  logic _2808_;
  logic _2809_;
  logic _2810_;
  logic _2811_;
  logic _2812_;
  logic _2813_;
  logic _2814_;
  logic _2815_;
  logic _2816_;
  logic _2817_;
  logic _2818_;
  logic _2819_;
  logic _2820_;
  logic _2821_;
  logic _2822_;
  logic _2823_;
  logic _2824_;
  logic _2825_;
  logic _2826_;
  logic _2827_;
  logic _2828_;
  logic _2829_;
  logic _2830_;
  logic _2831_;
  logic _2832_;
  logic _2833_;
  logic _2834_;
  logic _2835_;
  logic _2836_;
  logic [7:0] _2837_;
  logic [7:0] _2838_;
  logic _2839_;
  logic _2840_;
  logic _2841_;
  logic _2842_;
  logic _2843_;
  logic _2844_;
  logic _2845_;
  logic _2846_;
  logic _2847_;
  logic _2848_;
  logic _2849_;
  logic _2850_;
  logic _2851_;
  logic _2852_;
  logic _2853_;
  logic _2854_;
  logic _2855_;
  logic _2856_;
  logic _2857_;
  logic _2858_;
  logic _2859_;
  logic _2860_;
  logic _2861_;
  logic _2862_;
  logic _2863_;
  logic _2864_;
  logic _2865_;
  logic _2866_;
  logic _2867_;
  logic _2868_;
  logic _2869_;
  logic _2870_;
  logic _2871_;
  logic _2872_;
  logic _2873_;
  logic _2874_;
  logic _2875_;
  logic _2876_;
  logic _2877_;
  logic _2878_;
  logic _2879_;
  logic _2880_;
  logic _2881_;
  logic _2882_;
  logic _2883_;
  logic _2884_;
  logic _2885_;
  logic _2886_;
  logic _2887_;
  logic _2888_;
  logic _2889_;
  logic _2890_;
  logic _2891_;
  logic _2892_;
  logic _2893_;
  logic _2894_;
  logic _2895_;
  logic _2896_;
  logic _2897_;
  logic _2898_;
  logic _2899_;
  logic _2900_;
  logic _2901_;
  logic _2902_;
  logic _2903_;
  logic _2904_;
  logic _2905_;
  logic _2906_;
  logic _2907_;
  logic _2908_;
  logic _2909_;
  logic _2910_;
  logic _2911_;
  logic _2912_;
  logic _2913_;
  logic _2914_;
  logic _2915_;
  logic _2916_;
  logic _2917_;
  logic _2918_;
  logic _2919_;
  logic _2920_;
  logic _2921_;
  logic _2922_;
  logic _2923_;
  logic _2924_;
  logic _2925_;
  logic _2926_;
  logic _2927_;
  logic _2928_;
  logic _2929_;
  logic _2930_;
  logic _2931_;
  logic _2932_;
  logic _2933_;
  logic _2934_;
  logic _2935_;
  logic _2936_;
  logic _2937_;
  logic _2938_;
  logic _2939_;
  logic _2940_;
  logic _2941_;
  logic _2942_;
  logic _2943_;
  logic _2944_;
  logic _2945_;
  logic _2946_;
  logic _2947_;
  logic _2948_;
  logic _2949_;
  logic _2950_;
  logic _2951_;
  logic _2952_;
  logic _2953_;
  logic _2954_;
  logic _2955_;
  logic _2956_;
  logic _2957_;
  logic _2958_;
  logic _2959_;
  logic _2960_;
  logic _2961_;
  logic _2962_;
  logic _2963_;
  logic _2964_;
  logic _2965_;
  logic _2966_;
  logic _2967_;
  logic _2968_;
  logic _2969_;
  logic _2970_;
  logic _2971_;
  logic _2972_;
  logic _2973_;
  logic _2974_;
  logic _2975_;
  logic _2976_;
  logic _2977_;
  logic _2978_;
  logic _2979_;
  logic _2980_;
  logic _2981_;
  logic _2982_;
  logic _2983_;
  logic _2984_;
  logic _2985_;
  logic _2986_;
  logic _2987_;
  logic _2988_;
  logic _2989_;
  logic _2990_;
  logic _2991_;
  logic _2992_;
  logic _2993_;
  logic _2994_;
  logic _2995_;
  logic _2996_;
  logic _2997_;
  logic _2998_;
  logic _2999_;
  logic _3000_;
  logic _3001_;
  logic _3002_;
  logic _3003_;
  logic _3004_;
  logic _3005_;
  logic _3006_;
  logic _3007_;
  logic _3008_;
  logic _3009_;
  logic _3010_;
  logic _3011_;
  logic _3012_;
  logic _3013_;
  logic _3014_;
  logic _3015_;
  logic _3016_;
  logic _3017_;
  logic _3018_;
  logic _3019_;
  logic _3020_;
  logic _3021_;
  logic _3022_;
  logic _3023_;
  logic _3024_;
  logic _3025_;
  logic _3026_;
  logic _3027_;
  logic _3028_;
  logic _3029_;
  logic _3030_;
  logic _3031_;
  logic _3032_;
  logic _3033_;
  logic _3034_;
  logic _3035_;
  logic _3036_;
  logic _3037_;
  logic _3038_;
  logic _3039_;
  logic _3040_;
  logic _3041_;
  logic _3042_;
  logic _3043_;
  logic _3044_;
  logic _3045_;
  logic _3046_;
  logic _3047_;
  logic _3048_;
  logic _3049_;
  logic _3050_;
  logic _3051_;
  logic _3052_;
  logic _3053_;
  logic _3054_;
  logic _3055_;
  logic _3056_;
  logic _3057_;
  logic _3058_;
  logic _3059_;
  logic _3060_;
  logic _3061_;
  logic _3062_;
  logic _3063_;
  logic _3064_;
  logic _3065_;
  logic _3066_;
  logic _3067_;
  logic _3068_;
  logic _3069_;
  logic _3070_;
  logic _3071_;
  logic _3072_;
  logic _3073_;
  logic _3074_;
  logic _3075_;
  logic _3076_;
  logic _3077_;
  logic _3078_;
  logic _3079_;
  logic _3080_;
  logic _3081_;
  logic _3082_;
  logic _3083_;
  logic _3084_;
  logic _3085_;
  logic _3086_;
  logic _3087_;
  logic _3088_;
  logic _3089_;
  logic _3090_;
  logic _3091_;
  logic _3092_;
  logic _3093_;
  logic _3094_;
  logic [7:0] _3095_;
  logic [7:0] _3096_;
  logic _3097_;
  logic _3098_;
  logic _3099_;
  logic _3100_;
  logic _3101_;
  logic _3102_;
  logic _3103_;
  logic _3104_;
  logic _3105_;
  logic _3106_;
  logic _3107_;
  logic _3108_;
  logic _3109_;
  logic _3110_;
  logic _3111_;
  logic _3112_;
  logic _3113_;
  logic _3114_;
  logic _3115_;
  logic _3116_;
  logic _3117_;
  logic _3118_;
  logic _3119_;
  logic _3120_;
  logic _3121_;
  logic _3122_;
  logic _3123_;
  logic _3124_;
  logic _3125_;
  logic _3126_;
  logic _3127_;
  logic _3128_;
  logic _3129_;
  logic _3130_;
  logic _3131_;
  logic _3132_;
  logic _3133_;
  logic _3134_;
  logic _3135_;
  logic _3136_;
  logic _3137_;
  logic _3138_;
  logic _3139_;
  logic _3140_;
  logic _3141_;
  logic _3142_;
  logic _3143_;
  logic _3144_;
  logic _3145_;
  logic _3146_;
  logic _3147_;
  logic _3148_;
  logic _3149_;
  logic _3150_;
  logic _3151_;
  logic _3152_;
  logic _3153_;
  logic _3154_;
  logic _3155_;
  logic _3156_;
  logic _3157_;
  logic _3158_;
  logic _3159_;
  logic _3160_;
  logic _3161_;
  logic _3162_;
  logic _3163_;
  logic _3164_;
  logic _3165_;
  logic _3166_;
  logic _3167_;
  logic _3168_;
  logic _3169_;
  logic _3170_;
  logic _3171_;
  logic _3172_;
  logic _3173_;
  logic _3174_;
  logic _3175_;
  logic _3176_;
  logic _3177_;
  logic _3178_;
  logic _3179_;
  logic _3180_;
  logic _3181_;
  logic _3182_;
  logic _3183_;
  logic _3184_;
  logic _3185_;
  logic _3186_;
  logic _3187_;
  logic _3188_;
  logic _3189_;
  logic _3190_;
  logic _3191_;
  logic _3192_;
  logic _3193_;
  logic _3194_;
  logic _3195_;
  logic _3196_;
  logic _3197_;
  logic _3198_;
  logic _3199_;
  logic _3200_;
  logic _3201_;
  logic _3202_;
  logic _3203_;
  logic _3204_;
  logic _3205_;
  logic _3206_;
  logic _3207_;
  logic _3208_;
  logic _3209_;
  logic _3210_;
  logic _3211_;
  logic _3212_;
  logic _3213_;
  logic _3214_;
  logic _3215_;
  logic _3216_;
  logic _3217_;
  logic _3218_;
  logic _3219_;
  logic _3220_;
  logic _3221_;
  logic _3222_;
  logic _3223_;
  logic _3224_;
  logic _3225_;
  logic _3226_;
  logic _3227_;
  logic _3228_;
  logic _3229_;
  logic _3230_;
  logic _3231_;
  logic _3232_;
  logic _3233_;
  logic _3234_;
  logic _3235_;
  logic _3236_;
  logic _3237_;
  logic _3238_;
  logic _3239_;
  logic _3240_;
  logic _3241_;
  logic _3242_;
  logic _3243_;
  logic _3244_;
  logic _3245_;
  logic _3246_;
  logic _3247_;
  logic _3248_;
  logic _3249_;
  logic _3250_;
  logic _3251_;
  logic _3252_;
  logic _3253_;
  logic _3254_;
  logic _3255_;
  logic _3256_;
  logic _3257_;
  logic _3258_;
  logic _3259_;
  logic _3260_;
  logic _3261_;
  logic _3262_;
  logic _3263_;
  logic _3264_;
  logic _3265_;
  logic _3266_;
  logic _3267_;
  logic _3268_;
  logic _3269_;
  logic _3270_;
  logic _3271_;
  logic _3272_;
  logic _3273_;
  logic _3274_;
  logic _3275_;
  logic _3276_;
  logic _3277_;
  logic _3278_;
  logic _3279_;
  logic _3280_;
  logic _3281_;
  logic _3282_;
  logic _3283_;
  logic _3284_;
  logic _3285_;
  logic _3286_;
  logic _3287_;
  logic _3288_;
  logic _3289_;
  logic _3290_;
  logic _3291_;
  logic _3292_;
  logic _3293_;
  logic _3294_;
  logic _3295_;
  logic _3296_;
  logic _3297_;
  logic _3298_;
  logic _3299_;
  logic _3300_;
  logic _3301_;
  logic _3302_;
  logic _3303_;
  logic _3304_;
  logic _3305_;
  logic _3306_;
  logic _3307_;
  logic _3308_;
  logic _3309_;
  logic _3310_;
  logic _3311_;
  logic _3312_;
  logic _3313_;
  logic _3314_;
  logic _3315_;
  logic _3316_;
  logic _3317_;
  logic _3318_;
  logic _3319_;
  logic _3320_;
  logic _3321_;
  logic _3322_;
  logic _3323_;
  logic _3324_;
  logic _3325_;
  logic _3326_;
  logic _3327_;
  logic _3328_;
  logic _3329_;
  logic _3330_;
  logic _3331_;
  logic _3332_;
  logic _3333_;
  logic _3334_;
  logic _3335_;
  logic _3336_;
  logic _3337_;
  logic _3338_;
  logic _3339_;
  logic _3340_;
  logic _3341_;
  logic _3342_;
  logic _3343_;
  logic _3344_;
  logic _3345_;
  logic _3346_;
  logic _3347_;
  logic _3348_;
  logic _3349_;
  logic _3350_;
  logic _3351_;
  logic _3352_;
  logic [7:0] _3353_;
  logic [7:0] _3354_;
  logic _3355_;
  logic _3356_;
  logic _3357_;
  logic _3358_;
  logic _3359_;
  logic _3360_;
  logic _3361_;
  logic _3362_;
  logic _3363_;
  logic _3364_;
  logic _3365_;
  logic _3366_;
  logic _3367_;
  logic _3368_;
  logic _3369_;
  logic _3370_;
  logic _3371_;
  logic _3372_;
  logic _3373_;
  logic _3374_;
  logic _3375_;
  logic _3376_;
  logic _3377_;
  logic _3378_;
  logic _3379_;
  logic _3380_;
  logic _3381_;
  logic _3382_;
  logic _3383_;
  logic _3384_;
  logic _3385_;
  logic _3386_;
  logic _3387_;
  logic _3388_;
  logic _3389_;
  logic _3390_;
  logic _3391_;
  logic _3392_;
  logic _3393_;
  logic _3394_;
  logic _3395_;
  logic _3396_;
  logic _3397_;
  logic _3398_;
  logic _3399_;
  logic _3400_;
  logic _3401_;
  logic _3402_;
  logic _3403_;
  logic _3404_;
  logic _3405_;
  logic _3406_;
  logic _3407_;
  logic _3408_;
  logic _3409_;
  logic _3410_;
  logic _3411_;
  logic _3412_;
  logic _3413_;
  logic _3414_;
  logic _3415_;
  logic _3416_;
  logic _3417_;
  logic _3418_;
  logic _3419_;
  logic _3420_;
  logic _3421_;
  logic _3422_;
  logic _3423_;
  logic _3424_;
  logic _3425_;
  logic _3426_;
  logic _3427_;
  logic _3428_;
  logic _3429_;
  logic _3430_;
  logic _3431_;
  logic _3432_;
  logic _3433_;
  logic _3434_;
  logic _3435_;
  logic _3436_;
  logic _3437_;
  logic _3438_;
  logic _3439_;
  logic _3440_;
  logic _3441_;
  logic _3442_;
  logic _3443_;
  logic _3444_;
  logic _3445_;
  logic _3446_;
  logic _3447_;
  logic _3448_;
  logic _3449_;
  logic _3450_;
  logic _3451_;
  logic _3452_;
  logic _3453_;
  logic _3454_;
  logic _3455_;
  logic _3456_;
  logic _3457_;
  logic _3458_;
  logic _3459_;
  logic _3460_;
  logic _3461_;
  logic _3462_;
  logic _3463_;
  logic _3464_;
  logic _3465_;
  logic _3466_;
  logic _3467_;
  logic _3468_;
  logic _3469_;
  logic _3470_;
  logic _3471_;
  logic _3472_;
  logic _3473_;
  logic _3474_;
  logic _3475_;
  logic _3476_;
  logic _3477_;
  logic _3478_;
  logic _3479_;
  logic _3480_;
  logic _3481_;
  logic _3482_;
  logic _3483_;
  logic _3484_;
  logic _3485_;
  logic _3486_;
  logic _3487_;
  logic _3488_;
  logic _3489_;
  logic _3490_;
  logic _3491_;
  logic _3492_;
  logic _3493_;
  logic _3494_;
  logic _3495_;
  logic _3496_;
  logic _3497_;
  logic _3498_;
  logic _3499_;
  logic _3500_;
  logic _3501_;
  logic _3502_;
  logic _3503_;
  logic _3504_;
  logic _3505_;
  logic _3506_;
  logic _3507_;
  logic _3508_;
  logic _3509_;
  logic _3510_;
  logic _3511_;
  logic _3512_;
  logic _3513_;
  logic _3514_;
  logic _3515_;
  logic _3516_;
  logic _3517_;
  logic _3518_;
  logic _3519_;
  logic _3520_;
  logic _3521_;
  logic _3522_;
  logic _3523_;
  logic _3524_;
  logic _3525_;
  logic _3526_;
  logic _3527_;
  logic _3528_;
  logic _3529_;
  logic _3530_;
  logic _3531_;
  logic _3532_;
  logic _3533_;
  logic _3534_;
  logic _3535_;
  logic _3536_;
  logic _3537_;
  logic _3538_;
  logic _3539_;
  logic _3540_;
  logic _3541_;
  logic _3542_;
  logic _3543_;
  logic _3544_;
  logic _3545_;
  logic _3546_;
  logic _3547_;
  logic _3548_;
  logic _3549_;
  logic _3550_;
  logic _3551_;
  logic _3552_;
  logic _3553_;
  logic _3554_;
  logic _3555_;
  logic _3556_;
  logic _3557_;
  logic _3558_;
  logic _3559_;
  logic _3560_;
  logic _3561_;
  logic _3562_;
  logic _3563_;
  logic _3564_;
  logic _3565_;
  logic _3566_;
  logic _3567_;
  logic _3568_;
  logic _3569_;
  logic _3570_;
  logic _3571_;
  logic _3572_;
  logic _3573_;
  logic _3574_;
  logic _3575_;
  logic _3576_;
  logic _3577_;
  logic _3578_;
  logic _3579_;
  logic _3580_;
  logic _3581_;
  logic _3582_;
  logic _3583_;
  logic _3584_;
  logic _3585_;
  logic _3586_;
  logic _3587_;
  logic _3588_;
  logic _3589_;
  logic _3590_;
  logic _3591_;
  logic _3592_;
  logic _3593_;
  logic _3594_;
  logic _3595_;
  logic _3596_;
  logic _3597_;
  logic _3598_;
  logic _3599_;
  logic _3600_;
  logic _3601_;
  logic _3602_;
  logic _3603_;
  logic _3604_;
  logic _3605_;
  logic _3606_;
  logic _3607_;
  logic _3608_;
  logic _3609_;
  logic _3610_;
  logic [7:0] _3611_;
  logic [7:0] _3612_;
  logic _3613_;
  logic _3614_;
  logic _3615_;
  logic _3616_;
  logic _3617_;
  logic _3618_;
  logic _3619_;
  logic _3620_;
  logic _3621_;
  logic _3622_;
  logic _3623_;
  logic _3624_;
  logic _3625_;
  logic _3626_;
  logic _3627_;
  logic _3628_;
  logic _3629_;
  logic _3630_;
  logic _3631_;
  logic _3632_;
  logic _3633_;
  logic _3634_;
  logic _3635_;
  logic _3636_;
  logic _3637_;
  logic _3638_;
  logic _3639_;
  logic _3640_;
  logic _3641_;
  logic _3642_;
  logic _3643_;
  logic _3644_;
  logic _3645_;
  logic _3646_;
  logic _3647_;
  logic _3648_;
  logic _3649_;
  logic _3650_;
  logic _3651_;
  logic _3652_;
  logic _3653_;
  logic _3654_;
  logic _3655_;
  logic _3656_;
  logic _3657_;
  logic _3658_;
  logic _3659_;
  logic _3660_;
  logic _3661_;
  logic _3662_;
  logic _3663_;
  logic _3664_;
  logic _3665_;
  logic _3666_;
  logic _3667_;
  logic _3668_;
  logic _3669_;
  logic _3670_;
  logic _3671_;
  logic _3672_;
  logic _3673_;
  logic _3674_;
  logic _3675_;
  logic _3676_;
  logic _3677_;
  logic _3678_;
  logic _3679_;
  logic _3680_;
  logic _3681_;
  logic _3682_;
  logic _3683_;
  logic _3684_;
  logic _3685_;
  logic _3686_;
  logic _3687_;
  logic _3688_;
  logic _3689_;
  logic _3690_;
  logic _3691_;
  logic _3692_;
  logic _3693_;
  logic _3694_;
  logic _3695_;
  logic _3696_;
  logic _3697_;
  logic _3698_;
  logic _3699_;
  logic _3700_;
  logic _3701_;
  logic _3702_;
  logic _3703_;
  logic _3704_;
  logic _3705_;
  logic _3706_;
  logic _3707_;
  logic _3708_;
  logic _3709_;
  logic _3710_;
  logic _3711_;
  logic _3712_;
  logic _3713_;
  logic _3714_;
  logic _3715_;
  logic _3716_;
  logic _3717_;
  logic _3718_;
  logic _3719_;
  logic _3720_;
  logic _3721_;
  logic _3722_;
  logic _3723_;
  logic _3724_;
  logic _3725_;
  logic _3726_;
  logic _3727_;
  logic _3728_;
  logic _3729_;
  logic _3730_;
  logic _3731_;
  logic _3732_;
  logic _3733_;
  logic _3734_;
  logic _3735_;
  logic _3736_;
  logic _3737_;
  logic _3738_;
  logic _3739_;
  logic _3740_;
  logic _3741_;
  logic _3742_;
  logic _3743_;
  logic _3744_;
  logic _3745_;
  logic _3746_;
  logic _3747_;
  logic _3748_;
  logic _3749_;
  logic _3750_;
  logic _3751_;
  logic _3752_;
  logic _3753_;
  logic _3754_;
  logic _3755_;
  logic _3756_;
  logic _3757_;
  logic _3758_;
  logic _3759_;
  logic _3760_;
  logic _3761_;
  logic _3762_;
  logic _3763_;
  logic _3764_;
  logic _3765_;
  logic _3766_;
  logic _3767_;
  logic _3768_;
  logic _3769_;
  logic _3770_;
  logic _3771_;
  logic _3772_;
  logic _3773_;
  logic _3774_;
  logic _3775_;
  logic _3776_;
  logic _3777_;
  logic _3778_;
  logic _3779_;
  logic _3780_;
  logic _3781_;
  logic _3782_;
  logic _3783_;
  logic _3784_;
  logic _3785_;
  logic _3786_;
  logic _3787_;
  logic _3788_;
  logic _3789_;
  logic _3790_;
  logic _3791_;
  logic _3792_;
  logic _3793_;
  logic _3794_;
  logic _3795_;
  logic _3796_;
  logic _3797_;
  logic _3798_;
  logic _3799_;
  logic _3800_;
  logic _3801_;
  logic _3802_;
  logic _3803_;
  logic _3804_;
  logic _3805_;
  logic _3806_;
  logic _3807_;
  logic _3808_;
  logic _3809_;
  logic _3810_;
  logic _3811_;
  logic _3812_;
  logic _3813_;
  logic _3814_;
  logic _3815_;
  logic _3816_;
  logic _3817_;
  logic _3818_;
  logic _3819_;
  logic _3820_;
  logic _3821_;
  logic _3822_;
  logic _3823_;
  logic _3824_;
  logic _3825_;
  logic _3826_;
  logic _3827_;
  logic _3828_;
  logic _3829_;
  logic _3830_;
  logic _3831_;
  logic _3832_;
  logic _3833_;
  logic _3834_;
  logic _3835_;
  logic _3836_;
  logic _3837_;
  logic _3838_;
  logic _3839_;
  logic _3840_;
  logic _3841_;
  logic _3842_;
  logic _3843_;
  logic _3844_;
  logic _3845_;
  logic _3846_;
  logic _3847_;
  logic _3848_;
  logic _3849_;
  logic _3850_;
  logic _3851_;
  logic _3852_;
  logic _3853_;
  logic _3854_;
  logic _3855_;
  logic _3856_;
  logic _3857_;
  logic _3858_;
  logic _3859_;
  logic _3860_;
  logic _3861_;
  logic _3862_;
  logic _3863_;
  logic _3864_;
  logic _3865_;
  logic _3866_;
  logic _3867_;
  logic _3868_;
  logic [7:0] _3869_;
  logic [7:0] _3870_;
  logic _3871_;
  logic _3872_;
  logic _3873_;
  logic _3874_;
  logic _3875_;
  logic _3876_;
  logic _3877_;
  logic _3878_;
  logic _3879_;
  logic _3880_;
  logic _3881_;
  logic _3882_;
  logic _3883_;
  logic _3884_;
  logic _3885_;
  logic _3886_;
  logic _3887_;
  logic _3888_;
  logic _3889_;
  logic _3890_;
  logic _3891_;
  logic _3892_;
  logic _3893_;
  logic _3894_;
  logic _3895_;
  logic _3896_;
  logic _3897_;
  logic _3898_;
  logic _3899_;
  logic _3900_;
  logic _3901_;
  logic _3902_;
  logic _3903_;
  logic _3904_;
  logic _3905_;
  logic _3906_;
  logic _3907_;
  logic _3908_;
  logic _3909_;
  logic _3910_;
  logic _3911_;
  logic _3912_;
  logic _3913_;
  logic _3914_;
  logic _3915_;
  logic _3916_;
  logic _3917_;
  logic _3918_;
  logic _3919_;
  logic _3920_;
  logic _3921_;
  logic _3922_;
  logic _3923_;
  logic _3924_;
  logic _3925_;
  logic _3926_;
  logic _3927_;
  logic _3928_;
  logic _3929_;
  logic _3930_;
  logic _3931_;
  logic _3932_;
  logic _3933_;
  logic _3934_;
  logic _3935_;
  logic _3936_;
  logic _3937_;
  logic _3938_;
  logic _3939_;
  logic _3940_;
  logic _3941_;
  logic _3942_;
  logic _3943_;
  logic _3944_;
  logic _3945_;
  logic _3946_;
  logic _3947_;
  logic _3948_;
  logic _3949_;
  logic _3950_;
  logic _3951_;
  logic _3952_;
  logic _3953_;
  logic _3954_;
  logic _3955_;
  logic _3956_;
  logic _3957_;
  logic _3958_;
  logic _3959_;
  logic _3960_;
  logic _3961_;
  logic _3962_;
  logic _3963_;
  logic _3964_;
  logic _3965_;
  logic _3966_;
  logic _3967_;
  logic _3968_;
  logic _3969_;
  logic _3970_;
  logic _3971_;
  logic _3972_;
  logic _3973_;
  logic _3974_;
  logic _3975_;
  logic _3976_;
  logic _3977_;
  logic _3978_;
  logic _3979_;
  logic _3980_;
  logic _3981_;
  logic _3982_;
  logic _3983_;
  logic _3984_;
  logic _3985_;
  logic _3986_;
  logic _3987_;
  logic _3988_;
  logic _3989_;
  logic _3990_;
  logic _3991_;
  logic _3992_;
  logic _3993_;
  logic _3994_;
  logic _3995_;
  logic _3996_;
  logic _3997_;
  logic _3998_;
  logic _3999_;
  logic _4000_;
  logic _4001_;
  logic _4002_;
  logic _4003_;
  logic _4004_;
  logic _4005_;
  logic _4006_;
  logic _4007_;
  logic _4008_;
  logic _4009_;
  logic _4010_;
  logic _4011_;
  logic _4012_;
  logic _4013_;
  logic _4014_;
  logic _4015_;
  logic _4016_;
  logic _4017_;
  logic _4018_;
  logic _4019_;
  logic _4020_;
  logic _4021_;
  logic _4022_;
  logic _4023_;
  logic _4024_;
  logic _4025_;
  logic _4026_;
  logic _4027_;
  logic _4028_;
  logic _4029_;
  logic _4030_;
  logic _4031_;
  logic _4032_;
  logic _4033_;
  logic _4034_;
  logic _4035_;
  logic _4036_;
  logic _4037_;
  logic _4038_;
  logic _4039_;
  logic _4040_;
  logic _4041_;
  logic _4042_;
  logic _4043_;
  logic _4044_;
  logic _4045_;
  logic _4046_;
  logic _4047_;
  logic _4048_;
  logic _4049_;
  logic _4050_;
  logic _4051_;
  logic _4052_;
  logic _4053_;
  logic _4054_;
  logic _4055_;
  logic _4056_;
  logic _4057_;
  logic _4058_;
  logic _4059_;
  logic _4060_;
  logic _4061_;
  logic _4062_;
  logic _4063_;
  logic _4064_;
  logic _4065_;
  logic _4066_;
  logic _4067_;
  logic _4068_;
  logic _4069_;
  logic _4070_;
  logic _4071_;
  logic _4072_;
  logic _4073_;
  logic _4074_;
  logic _4075_;
  logic _4076_;
  logic _4077_;
  logic _4078_;
  logic _4079_;
  logic _4080_;
  logic _4081_;
  logic _4082_;
  logic _4083_;
  logic _4084_;
  logic _4085_;
  logic _4086_;
  logic _4087_;
  logic _4088_;
  logic _4089_;
  logic _4090_;
  logic _4091_;
  logic _4092_;
  logic _4093_;
  logic _4094_;
  logic _4095_;
  logic _4096_;
  logic _4097_;
  logic _4098_;
  logic _4099_;
  logic _4100_;
  logic _4101_;
  logic _4102_;
  logic _4103_;
  logic _4104_;
  logic _4105_;
  logic _4106_;
  logic _4107_;
  logic _4108_;
  logic _4109_;
  logic _4110_;
  logic _4111_;
  logic _4112_;
  logic _4113_;
  logic _4114_;
  logic _4115_;
  logic _4116_;
  logic _4117_;
  logic _4118_;
  logic _4119_;
  logic _4120_;
  logic _4121_;
  logic _4122_;
  logic _4123_;
  logic _4124_;
  logic _4125_;
  logic _4126_;
  logic [7:0] _4127_;
  logic [31:0] _4128_;
  logic [31:0] _4129_;
  logic [31:0] _4130_;
  logic [31:0] _4131_;
  logic [31:0] _4132_;
  logic [31:0] _4133_;
  logic [31:0] _4134_;
  logic [31:0] _4135_;
  logic [31:0] _4136_;
  logic [31:0] _4137_;
  logic [31:0] _4138_;
  logic [31:0] _4139_;
  input clk;
  logic [31:0] k0;
  logic [31:0] k1;
  logic [31:0] k2;
  logic [31:0] k3;
  input [127:0] key;
  logic [31:0] p00;
  logic [31:0] p01;
  logic [31:0] p02;
  logic [31:0] p03;
  logic [31:0] p10;
  logic [31:0] p11;
  logic [31:0] p12;
  logic [31:0] p13;
  logic [31:0] p20;
  logic [31:0] p21;
  logic [31:0] p22;
  logic [31:0] p23;
  logic [31:0] p30;
  logic [31:0] p31;
  logic [31:0] p32;
  logic [31:0] p33;
  logic [31:0] s0;
  logic [31:0] s1;
  logic [31:0] s2;
  logic [31:0] s3;
  input [127:0] state_in;
  output [127:0] state_out;
  logic [127:0] state_out;
  logic [7:0] \t0.b0 ;
  logic [7:0] \t0.b1 ;
  logic [7:0] \t0.b2 ;
  logic [7:0] \t0.b3 ;
  logic \t0.clk ;
  logic [31:0] \t0.p0 ;
  logic [31:0] \t0.p1 ;
  logic [31:0] \t0.p2 ;
  logic [31:0] \t0.p3 ;
  logic [31:0] \t0.state ;
  logic \t0.t0.clk ;
  logic [7:0] \t0.t0.in ;
  logic [31:0] \t0.t0.out ;
  logic \t0.t0.s0.clk ;
  logic [7:0] \t0.t0.s0.in ;
  logic [7:0] \t0.t0.s0.out ;
  logic \t0.t0.s4.clk ;
  logic [7:0] \t0.t0.s4.in ;
  logic [7:0] \t0.t0.s4.out ;
  logic \t0.t1.clk ;
  logic [7:0] \t0.t1.in ;
  logic [31:0] \t0.t1.out ;
  logic \t0.t1.s0.clk ;
  logic [7:0] \t0.t1.s0.in ;
  logic [7:0] \t0.t1.s0.out ;
  logic \t0.t1.s4.clk ;
  logic [7:0] \t0.t1.s4.in ;
  logic [7:0] \t0.t1.s4.out ;
  logic \t0.t2.clk ;
  logic [7:0] \t0.t2.in ;
  logic [31:0] \t0.t2.out ;
  logic \t0.t2.s0.clk ;
  logic [7:0] \t0.t2.s0.in ;
  logic [7:0] \t0.t2.s0.out ;
  logic \t0.t2.s4.clk ;
  logic [7:0] \t0.t2.s4.in ;
  logic [7:0] \t0.t2.s4.out ;
  logic \t0.t3.clk ;
  logic [7:0] \t0.t3.in ;
  logic [31:0] \t0.t3.out ;
  logic \t0.t3.s0.clk ;
  logic [7:0] \t0.t3.s0.in ;
  logic [7:0] \t0.t3.s0.out ;
  logic \t0.t3.s4.clk ;
  logic [7:0] \t0.t3.s4.in ;
  logic [7:0] \t0.t3.s4.out ;
  logic [7:0] \t1.b0 ;
  logic [7:0] \t1.b1 ;
  logic [7:0] \t1.b2 ;
  logic [7:0] \t1.b3 ;
  logic \t1.clk ;
  logic [31:0] \t1.p0 ;
  logic [31:0] \t1.p1 ;
  logic [31:0] \t1.p2 ;
  logic [31:0] \t1.p3 ;
  logic [31:0] \t1.state ;
  logic \t1.t0.clk ;
  logic [7:0] \t1.t0.in ;
  logic [31:0] \t1.t0.out ;
  logic \t1.t0.s0.clk ;
  logic [7:0] \t1.t0.s0.in ;
  logic [7:0] \t1.t0.s0.out ;
  logic \t1.t0.s4.clk ;
  logic [7:0] \t1.t0.s4.in ;
  logic [7:0] \t1.t0.s4.out ;
  logic \t1.t1.clk ;
  logic [7:0] \t1.t1.in ;
  logic [31:0] \t1.t1.out ;
  logic \t1.t1.s0.clk ;
  logic [7:0] \t1.t1.s0.in ;
  logic [7:0] \t1.t1.s0.out ;
  logic \t1.t1.s4.clk ;
  logic [7:0] \t1.t1.s4.in ;
  logic [7:0] \t1.t1.s4.out ;
  logic \t1.t2.clk ;
  logic [7:0] \t1.t2.in ;
  logic [31:0] \t1.t2.out ;
  logic \t1.t2.s0.clk ;
  logic [7:0] \t1.t2.s0.in ;
  logic [7:0] \t1.t2.s0.out ;
  logic \t1.t2.s4.clk ;
  logic [7:0] \t1.t2.s4.in ;
  logic [7:0] \t1.t2.s4.out ;
  logic \t1.t3.clk ;
  logic [7:0] \t1.t3.in ;
  logic [31:0] \t1.t3.out ;
  logic \t1.t3.s0.clk ;
  logic [7:0] \t1.t3.s0.in ;
  logic [7:0] \t1.t3.s0.out ;
  logic \t1.t3.s4.clk ;
  logic [7:0] \t1.t3.s4.in ;
  logic [7:0] \t1.t3.s4.out ;
  logic [7:0] \t2.b0 ;
  logic [7:0] \t2.b1 ;
  logic [7:0] \t2.b2 ;
  logic [7:0] \t2.b3 ;
  logic \t2.clk ;
  logic [31:0] \t2.p0 ;
  logic [31:0] \t2.p1 ;
  logic [31:0] \t2.p2 ;
  logic [31:0] \t2.p3 ;
  logic [31:0] \t2.state ;
  logic \t2.t0.clk ;
  logic [7:0] \t2.t0.in ;
  logic [31:0] \t2.t0.out ;
  logic \t2.t0.s0.clk ;
  logic [7:0] \t2.t0.s0.in ;
  logic [7:0] \t2.t0.s0.out ;
  logic \t2.t0.s4.clk ;
  logic [7:0] \t2.t0.s4.in ;
  logic [7:0] \t2.t0.s4.out ;
  logic \t2.t1.clk ;
  logic [7:0] \t2.t1.in ;
  logic [31:0] \t2.t1.out ;
  logic \t2.t1.s0.clk ;
  logic [7:0] \t2.t1.s0.in ;
  logic [7:0] \t2.t1.s0.out ;
  logic \t2.t1.s4.clk ;
  logic [7:0] \t2.t1.s4.in ;
  logic [7:0] \t2.t1.s4.out ;
  logic \t2.t2.clk ;
  logic [7:0] \t2.t2.in ;
  logic [31:0] \t2.t2.out ;
  logic \t2.t2.s0.clk ;
  logic [7:0] \t2.t2.s0.in ;
  logic [7:0] \t2.t2.s0.out ;
  logic \t2.t2.s4.clk ;
  logic [7:0] \t2.t2.s4.in ;
  logic [7:0] \t2.t2.s4.out ;
  logic \t2.t3.clk ;
  logic [7:0] \t2.t3.in ;
  logic [31:0] \t2.t3.out ;
  logic \t2.t3.s0.clk ;
  logic [7:0] \t2.t3.s0.in ;
  logic [7:0] \t2.t3.s0.out ;
  logic \t2.t3.s4.clk ;
  logic [7:0] \t2.t3.s4.in ;
  logic [7:0] \t2.t3.s4.out ;
  logic [7:0] \t3.b0 ;
  logic [7:0] \t3.b1 ;
  logic [7:0] \t3.b2 ;
  logic [7:0] \t3.b3 ;
  logic \t3.clk ;
  logic [31:0] \t3.p0 ;
  logic [31:0] \t3.p1 ;
  logic [31:0] \t3.p2 ;
  logic [31:0] \t3.p3 ;
  logic [31:0] \t3.state ;
  logic \t3.t0.clk ;
  logic [7:0] \t3.t0.in ;
  logic [31:0] \t3.t0.out ;
  logic \t3.t0.s0.clk ;
  logic [7:0] \t3.t0.s0.in ;
  logic [7:0] \t3.t0.s0.out ;
  logic \t3.t0.s4.clk ;
  logic [7:0] \t3.t0.s4.in ;
  logic [7:0] \t3.t0.s4.out ;
  logic \t3.t1.clk ;
  logic [7:0] \t3.t1.in ;
  logic [31:0] \t3.t1.out ;
  logic \t3.t1.s0.clk ;
  logic [7:0] \t3.t1.s0.in ;
  logic [7:0] \t3.t1.s0.out ;
  logic \t3.t1.s4.clk ;
  logic [7:0] \t3.t1.s4.in ;
  logic [7:0] \t3.t1.s4.out ;
  logic \t3.t2.clk ;
  logic [7:0] \t3.t2.in ;
  logic [31:0] \t3.t2.out ;
  logic \t3.t2.s0.clk ;
  logic [7:0] \t3.t2.s0.in ;
  logic [7:0] \t3.t2.s0.out ;
  logic \t3.t2.s4.clk ;
  logic [7:0] \t3.t2.s4.in ;
  logic [7:0] \t3.t2.s4.out ;
  logic \t3.t3.clk ;
  logic [7:0] \t3.t3.in ;
  logic [31:0] \t3.t3.out ;
  logic \t3.t3.s0.clk ;
  logic [7:0] \t3.t3.s0.in ;
  logic [7:0] \t3.t3.s0.out ;
  logic \t3.t3.s4.clk ;
  logic [7:0] \t3.t3.s4.in ;
  logic [7:0] \t3.t3.s4.out ;
  logic [31:0] z0;
  logic [31:0] z1;
  logic [31:0] z2;
  logic [31:0] z3;

  logic [127:0] fangyuan0;
  assign fangyuan0 = { z0, z1, z2, z3 };
  always @(posedge clk)
      state_out <= fangyuan0;
  assign p00[7:0] = \t0.t0.s0.out ^ \t0.t0.s4.out ;
  always @(posedge clk)
      \t0.t0.s0.out <= _0000_;
  logic [255:0] fangyuan1;
  assign fangyuan1 = { _0256_, _0255_, _0254_, _0253_, _0252_, _0251_, _0250_, _0249_, _0248_, _0247_, _0246_, _0245_, _0244_, _0243_, _0242_, _0241_, _0240_, _0239_, _0238_, _0237_, _0236_, _0235_, _0234_, _0233_, _0232_, _0231_, _0230_, _0229_, _0228_, _0227_, _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0220_, _0219_, _0218_, _0217_, _0216_, _0215_, _0214_, _0213_, _0212_, _0211_, _0210_, _0209_, _0208_, _0207_, _0206_, _0205_, _0204_, _0203_, _0202_, _0201_, _0200_, _0199_, _0198_, _0197_, _0196_, _0195_, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0186_, _0185_, _0184_, _0183_, _0182_, _0181_, _0180_, _0179_, _0178_, _0177_, _0176_, _0175_, _0174_, _0173_, _0172_, _0171_, _0170_, _0169_, _0168_, _0167_, _0166_, _0165_, _0164_, _0163_, _0162_, _0161_, _0160_, _0159_, _0158_, _0157_, _0156_, _0155_, _0154_, _0153_, _0152_, _0151_, _0150_, _0149_, _0148_, _0147_, _0146_, _0145_, _0144_, _0143_, _0142_, _0141_, _0140_, _0139_, _0138_, _0137_, _0136_, _0135_, _0134_, _0133_, _0132_, _0131_, _0130_, _0129_, _0128_, _0127_, _0126_, _0125_, _0124_, _0123_, _0122_, _0121_, _0120_, _0119_, _0118_, _0117_, _0116_, _0115_, _0114_, _0113_, _0112_, _0111_, _0110_, _0109_, _0108_, _0107_, _0106_, _0105_, _0104_, _0103_, _0102_, _0101_, _0100_, _0099_, _0098_, _0097_, _0096_, _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0085_, _0084_, _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0074_, _0073_, _0072_, _0071_, _0070_, _0069_, _0068_, _0067_, _0066_, _0065_, _0064_, _0063_, _0062_, _0061_, _0060_, _0059_, _0058_, _0057_, _0056_, _0055_, _0054_, _0053_, _0052_, _0051_, _0050_, _0049_, _0048_, _0047_, _0046_, _0045_, _0044_, _0043_, _0042_, _0041_, _0040_, _0039_, _0038_, _0037_, _0036_, _0035_, _0034_, _0033_, _0032_, _0031_, _0030_, _0029_, _0028_, _0027_, _0026_, _0025_, _0024_, _0023_, _0022_, _0021_, _0020_, _0019_, _0018_, _0017_, _0016_, _0015_, _0014_, _0013_, _0012_, _0011_, _0010_, _0009_, _0008_, _0007_, _0006_, _0005_, _0004_, _0003_, _0002_, _0001_ };

  always @(\t0.t0.s0.out or fangyuan1) begin
    casez (fangyuan1)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0000_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0000_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0000_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0000_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0000_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0000_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0000_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0000_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0000_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0000_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0000_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0000_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0000_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0000_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0000_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0000_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0000_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0000_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0000_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0000_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0000_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0000_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0000_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0000_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0000_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0000_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0000_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0000_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0000_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0000_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0000_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0000_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0000_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0000_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0000_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0000_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0000_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0000_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0000_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0000_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0000_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0000_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0000_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0000_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0000_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0000_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0000_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0000_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0000_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0000_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0000_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0000_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0000_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0000_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0000_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0000_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0000_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0000_ = 8'b01100011 ;
      default:
        _0000_ = \t0.t0.s0.out ;
    endcase
  end
  assign _0001_ = state_in[127:120] == 8'b11111111;
  assign _0002_ = state_in[127:120] == 8'b11111110;
  assign _0003_ = state_in[127:120] == 8'b11111101;
  assign _0004_ = state_in[127:120] == 8'b11111100;
  assign _0005_ = state_in[127:120] == 8'b11111011;
  assign _0006_ = state_in[127:120] == 8'b11111010;
  assign _0007_ = state_in[127:120] == 8'b11111001;
  assign _0008_ = state_in[127:120] == 8'b11111000;
  assign _0009_ = state_in[127:120] == 8'b11110111;
  assign _0010_ = state_in[127:120] == 8'b11110110;
  assign _0011_ = state_in[127:120] == 8'b11110101;
  assign _0012_ = state_in[127:120] == 8'b11110100;
  assign _0013_ = state_in[127:120] == 8'b11110011;
  assign _0014_ = state_in[127:120] == 8'b11110010;
  assign _0015_ = state_in[127:120] == 8'b11110001;
  assign _0016_ = state_in[127:120] == 8'b11110000;
  assign _0017_ = state_in[127:120] == 8'b11101111;
  assign _0018_ = state_in[127:120] == 8'b11101110;
  assign _0019_ = state_in[127:120] == 8'b11101101;
  assign _0020_ = state_in[127:120] == 8'b11101100;
  assign _0021_ = state_in[127:120] == 8'b11101011;
  assign _0022_ = state_in[127:120] == 8'b11101010;
  assign _0023_ = state_in[127:120] == 8'b11101001;
  assign _0024_ = state_in[127:120] == 8'b11101000;
  assign _0025_ = state_in[127:120] == 8'b11100111;
  assign _0026_ = state_in[127:120] == 8'b11100110;
  assign _0027_ = state_in[127:120] == 8'b11100101;
  assign _0028_ = state_in[127:120] == 8'b11100100;
  assign _0029_ = state_in[127:120] == 8'b11100011;
  assign _0030_ = state_in[127:120] == 8'b11100010;
  assign _0031_ = state_in[127:120] == 8'b11100001;
  assign _0032_ = state_in[127:120] == 8'b11100000;
  assign _0033_ = state_in[127:120] == 8'b11011111;
  assign _0034_ = state_in[127:120] == 8'b11011110;
  assign _0035_ = state_in[127:120] == 8'b11011101;
  assign _0036_ = state_in[127:120] == 8'b11011100;
  assign _0037_ = state_in[127:120] == 8'b11011011;
  assign _0038_ = state_in[127:120] == 8'b11011010;
  assign _0039_ = state_in[127:120] == 8'b11011001;
  assign _0040_ = state_in[127:120] == 8'b11011000;
  assign _0041_ = state_in[127:120] == 8'b11010111;
  assign _0042_ = state_in[127:120] == 8'b11010110;
  assign _0043_ = state_in[127:120] == 8'b11010101;
  assign _0044_ = state_in[127:120] == 8'b11010100;
  assign _0045_ = state_in[127:120] == 8'b11010011;
  assign _0046_ = state_in[127:120] == 8'b11010010;
  assign _0047_ = state_in[127:120] == 8'b11010001;
  assign _0048_ = state_in[127:120] == 8'b11010000;
  assign _0049_ = state_in[127:120] == 8'b11001111;
  assign _0050_ = state_in[127:120] == 8'b11001110;
  assign _0051_ = state_in[127:120] == 8'b11001101;
  assign _0052_ = state_in[127:120] == 8'b11001100;
  assign _0053_ = state_in[127:120] == 8'b11001011;
  assign _0054_ = state_in[127:120] == 8'b11001010;
  assign _0055_ = state_in[127:120] == 8'b11001001;
  assign _0056_ = state_in[127:120] == 8'b11001000;
  assign _0057_ = state_in[127:120] == 8'b11000111;
  assign _0058_ = state_in[127:120] == 8'b11000110;
  assign _0059_ = state_in[127:120] == 8'b11000101;
  assign _0060_ = state_in[127:120] == 8'b11000100;
  assign _0061_ = state_in[127:120] == 8'b11000011;
  assign _0062_ = state_in[127:120] == 8'b11000010;
  assign _0063_ = state_in[127:120] == 8'b11000001;
  assign _0064_ = state_in[127:120] == 8'b11000000;
  assign _0065_ = state_in[127:120] == 8'b10111111;
  assign _0066_ = state_in[127:120] == 8'b10111110;
  assign _0067_ = state_in[127:120] == 8'b10111101;
  assign _0068_ = state_in[127:120] == 8'b10111100;
  assign _0069_ = state_in[127:120] == 8'b10111011;
  assign _0070_ = state_in[127:120] == 8'b10111010;
  assign _0071_ = state_in[127:120] == 8'b10111001;
  assign _0072_ = state_in[127:120] == 8'b10111000;
  assign _0073_ = state_in[127:120] == 8'b10110111;
  assign _0074_ = state_in[127:120] == 8'b10110110;
  assign _0075_ = state_in[127:120] == 8'b10110101;
  assign _0076_ = state_in[127:120] == 8'b10110100;
  assign _0077_ = state_in[127:120] == 8'b10110011;
  assign _0078_ = state_in[127:120] == 8'b10110010;
  assign _0079_ = state_in[127:120] == 8'b10110001;
  assign _0080_ = state_in[127:120] == 8'b10110000;
  assign _0081_ = state_in[127:120] == 8'b10101111;
  assign _0082_ = state_in[127:120] == 8'b10101110;
  assign _0083_ = state_in[127:120] == 8'b10101101;
  assign _0084_ = state_in[127:120] == 8'b10101100;
  assign _0085_ = state_in[127:120] == 8'b10101011;
  assign _0086_ = state_in[127:120] == 8'b10101010;
  assign _0087_ = state_in[127:120] == 8'b10101001;
  assign _0088_ = state_in[127:120] == 8'b10101000;
  assign _0089_ = state_in[127:120] == 8'b10100111;
  assign _0090_ = state_in[127:120] == 8'b10100110;
  assign _0091_ = state_in[127:120] == 8'b10100101;
  assign _0092_ = state_in[127:120] == 8'b10100100;
  assign _0093_ = state_in[127:120] == 8'b10100011;
  assign _0094_ = state_in[127:120] == 8'b10100010;
  assign _0095_ = state_in[127:120] == 8'b10100001;
  assign _0096_ = state_in[127:120] == 8'b10100000;
  assign _0097_ = state_in[127:120] == 8'b10011111;
  assign _0098_ = state_in[127:120] == 8'b10011110;
  assign _0099_ = state_in[127:120] == 8'b10011101;
  assign _0100_ = state_in[127:120] == 8'b10011100;
  assign _0101_ = state_in[127:120] == 8'b10011011;
  assign _0102_ = state_in[127:120] == 8'b10011010;
  assign _0103_ = state_in[127:120] == 8'b10011001;
  assign _0104_ = state_in[127:120] == 8'b10011000;
  assign _0105_ = state_in[127:120] == 8'b10010111;
  assign _0106_ = state_in[127:120] == 8'b10010110;
  assign _0107_ = state_in[127:120] == 8'b10010101;
  assign _0108_ = state_in[127:120] == 8'b10010100;
  assign _0109_ = state_in[127:120] == 8'b10010011;
  assign _0110_ = state_in[127:120] == 8'b10010010;
  assign _0111_ = state_in[127:120] == 8'b10010001;
  assign _0112_ = state_in[127:120] == 8'b10010000;
  assign _0113_ = state_in[127:120] == 8'b10001111;
  assign _0114_ = state_in[127:120] == 8'b10001110;
  assign _0115_ = state_in[127:120] == 8'b10001101;
  assign _0116_ = state_in[127:120] == 8'b10001100;
  assign _0117_ = state_in[127:120] == 8'b10001011;
  assign _0118_ = state_in[127:120] == 8'b10001010;
  assign _0119_ = state_in[127:120] == 8'b10001001;
  assign _0120_ = state_in[127:120] == 8'b10001000;
  assign _0121_ = state_in[127:120] == 8'b10000111;
  assign _0122_ = state_in[127:120] == 8'b10000110;
  assign _0123_ = state_in[127:120] == 8'b10000101;
  assign _0124_ = state_in[127:120] == 8'b10000100;
  assign _0125_ = state_in[127:120] == 8'b10000011;
  assign _0126_ = state_in[127:120] == 8'b10000010;
  assign _0127_ = state_in[127:120] == 8'b10000001;
  assign _0128_ = state_in[127:120] == 8'b10000000;
  assign _0129_ = state_in[127:120] == 7'b1111111;
  assign _0130_ = state_in[127:120] == 7'b1111110;
  assign _0131_ = state_in[127:120] == 7'b1111101;
  assign _0132_ = state_in[127:120] == 7'b1111100;
  assign _0133_ = state_in[127:120] == 7'b1111011;
  assign _0134_ = state_in[127:120] == 7'b1111010;
  assign _0135_ = state_in[127:120] == 7'b1111001;
  assign _0136_ = state_in[127:120] == 7'b1111000;
  assign _0137_ = state_in[127:120] == 7'b1110111;
  assign _0138_ = state_in[127:120] == 7'b1110110;
  assign _0139_ = state_in[127:120] == 7'b1110101;
  assign _0140_ = state_in[127:120] == 7'b1110100;
  assign _0141_ = state_in[127:120] == 7'b1110011;
  assign _0142_ = state_in[127:120] == 7'b1110010;
  assign _0143_ = state_in[127:120] == 7'b1110001;
  assign _0144_ = state_in[127:120] == 7'b1110000;
  assign _0145_ = state_in[127:120] == 7'b1101111;
  assign _0146_ = state_in[127:120] == 7'b1101110;
  assign _0147_ = state_in[127:120] == 7'b1101101;
  assign _0148_ = state_in[127:120] == 7'b1101100;
  assign _0149_ = state_in[127:120] == 7'b1101011;
  assign _0150_ = state_in[127:120] == 7'b1101010;
  assign _0151_ = state_in[127:120] == 7'b1101001;
  assign _0152_ = state_in[127:120] == 7'b1101000;
  assign _0153_ = state_in[127:120] == 7'b1100111;
  assign _0154_ = state_in[127:120] == 7'b1100110;
  assign _0155_ = state_in[127:120] == 7'b1100101;
  assign _0156_ = state_in[127:120] == 7'b1100100;
  assign _0157_ = state_in[127:120] == 7'b1100011;
  assign _0158_ = state_in[127:120] == 7'b1100010;
  assign _0159_ = state_in[127:120] == 7'b1100001;
  assign _0160_ = state_in[127:120] == 7'b1100000;
  assign _0161_ = state_in[127:120] == 7'b1011111;
  assign _0162_ = state_in[127:120] == 7'b1011110;
  assign _0163_ = state_in[127:120] == 7'b1011101;
  assign _0164_ = state_in[127:120] == 7'b1011100;
  assign _0165_ = state_in[127:120] == 7'b1011011;
  assign _0166_ = state_in[127:120] == 7'b1011010;
  assign _0167_ = state_in[127:120] == 7'b1011001;
  assign _0168_ = state_in[127:120] == 7'b1011000;
  assign _0169_ = state_in[127:120] == 7'b1010111;
  assign _0170_ = state_in[127:120] == 7'b1010110;
  assign _0171_ = state_in[127:120] == 7'b1010101;
  assign _0172_ = state_in[127:120] == 7'b1010100;
  assign _0173_ = state_in[127:120] == 7'b1010011;
  assign _0174_ = state_in[127:120] == 7'b1010010;
  assign _0175_ = state_in[127:120] == 7'b1010001;
  assign _0176_ = state_in[127:120] == 7'b1010000;
  assign _0177_ = state_in[127:120] == 7'b1001111;
  assign _0178_ = state_in[127:120] == 7'b1001110;
  assign _0179_ = state_in[127:120] == 7'b1001101;
  assign _0180_ = state_in[127:120] == 7'b1001100;
  assign _0181_ = state_in[127:120] == 7'b1001011;
  assign _0182_ = state_in[127:120] == 7'b1001010;
  assign _0183_ = state_in[127:120] == 7'b1001001;
  assign _0184_ = state_in[127:120] == 7'b1001000;
  assign _0185_ = state_in[127:120] == 7'b1000111;
  assign _0186_ = state_in[127:120] == 7'b1000110;
  assign _0187_ = state_in[127:120] == 7'b1000101;
  assign _0188_ = state_in[127:120] == 7'b1000100;
  assign _0189_ = state_in[127:120] == 7'b1000011;
  assign _0190_ = state_in[127:120] == 7'b1000010;
  assign _0191_ = state_in[127:120] == 7'b1000001;
  assign _0192_ = state_in[127:120] == 7'b1000000;
  assign _0193_ = state_in[127:120] == 6'b111111;
  assign _0194_ = state_in[127:120] == 6'b111110;
  assign _0195_ = state_in[127:120] == 6'b111101;
  assign _0196_ = state_in[127:120] == 6'b111100;
  assign _0197_ = state_in[127:120] == 6'b111011;
  assign _0198_ = state_in[127:120] == 6'b111010;
  assign _0199_ = state_in[127:120] == 6'b111001;
  assign _0200_ = state_in[127:120] == 6'b111000;
  assign _0201_ = state_in[127:120] == 6'b110111;
  assign _0202_ = state_in[127:120] == 6'b110110;
  assign _0203_ = state_in[127:120] == 6'b110101;
  assign _0204_ = state_in[127:120] == 6'b110100;
  assign _0205_ = state_in[127:120] == 6'b110011;
  assign _0206_ = state_in[127:120] == 6'b110010;
  assign _0207_ = state_in[127:120] == 6'b110001;
  assign _0208_ = state_in[127:120] == 6'b110000;
  assign _0209_ = state_in[127:120] == 6'b101111;
  assign _0210_ = state_in[127:120] == 6'b101110;
  assign _0211_ = state_in[127:120] == 6'b101101;
  assign _0212_ = state_in[127:120] == 6'b101100;
  assign _0213_ = state_in[127:120] == 6'b101011;
  assign _0214_ = state_in[127:120] == 6'b101010;
  assign _0215_ = state_in[127:120] == 6'b101001;
  assign _0216_ = state_in[127:120] == 6'b101000;
  assign _0217_ = state_in[127:120] == 6'b100111;
  assign _0218_ = state_in[127:120] == 6'b100110;
  assign _0219_ = state_in[127:120] == 6'b100101;
  assign _0220_ = state_in[127:120] == 6'b100100;
  assign _0221_ = state_in[127:120] == 6'b100011;
  assign _0222_ = state_in[127:120] == 6'b100010;
  assign _0223_ = state_in[127:120] == 6'b100001;
  assign _0224_ = state_in[127:120] == 6'b100000;
  assign _0225_ = state_in[127:120] == 5'b11111;
  assign _0226_ = state_in[127:120] == 5'b11110;
  assign _0227_ = state_in[127:120] == 5'b11101;
  assign _0228_ = state_in[127:120] == 5'b11100;
  assign _0229_ = state_in[127:120] == 5'b11011;
  assign _0230_ = state_in[127:120] == 5'b11010;
  assign _0231_ = state_in[127:120] == 5'b11001;
  assign _0232_ = state_in[127:120] == 5'b11000;
  assign _0233_ = state_in[127:120] == 5'b10111;
  assign _0234_ = state_in[127:120] == 5'b10110;
  assign _0235_ = state_in[127:120] == 5'b10101;
  assign _0236_ = state_in[127:120] == 5'b10100;
  assign _0237_ = state_in[127:120] == 5'b10011;
  assign _0238_ = state_in[127:120] == 5'b10010;
  assign _0239_ = state_in[127:120] == 5'b10001;
  assign _0240_ = state_in[127:120] == 5'b10000;
  assign _0241_ = state_in[127:120] == 4'b1111;
  assign _0242_ = state_in[127:120] == 4'b1110;
  assign _0243_ = state_in[127:120] == 4'b1101;
  assign _0244_ = state_in[127:120] == 4'b1100;
  assign _0245_ = state_in[127:120] == 4'b1011;
  assign _0246_ = state_in[127:120] == 4'b1010;
  assign _0247_ = state_in[127:120] == 4'b1001;
  assign _0248_ = state_in[127:120] == 4'b1000;
  assign _0249_ = state_in[127:120] == 3'b111;
  assign _0250_ = state_in[127:120] == 3'b110;
  assign _0251_ = state_in[127:120] == 3'b101;
  assign _0252_ = state_in[127:120] == 3'b100;
  assign _0253_ = state_in[127:120] == 2'b11;
  assign _0254_ = state_in[127:120] == 2'b10;
  assign _0255_ = state_in[127:120] == 1'b1;
  assign _0256_ = ! state_in[127:120];
  always @(posedge clk)
      \t0.t0.s4.out <= _0257_;
  logic [255:0] fangyuan2;
  assign fangyuan2 = { _0256_, _0255_, _0254_, _0253_, _0252_, _0251_, _0250_, _0249_, _0248_, _0247_, _0246_, _0245_, _0244_, _0243_, _0242_, _0241_, _0240_, _0239_, _0238_, _0237_, _0236_, _0235_, _0234_, _0233_, _0232_, _0231_, _0230_, _0229_, _0228_, _0227_, _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0220_, _0219_, _0218_, _0217_, _0216_, _0215_, _0214_, _0213_, _0212_, _0211_, _0210_, _0209_, _0208_, _0207_, _0206_, _0205_, _0204_, _0203_, _0202_, _0201_, _0200_, _0199_, _0198_, _0197_, _0196_, _0195_, _0194_, _0193_, _0192_, _0191_, _0190_, _0189_, _0188_, _0187_, _0186_, _0185_, _0184_, _0183_, _0182_, _0181_, _0180_, _0179_, _0178_, _0177_, _0176_, _0175_, _0174_, _0173_, _0172_, _0171_, _0170_, _0169_, _0168_, _0167_, _0166_, _0165_, _0164_, _0163_, _0162_, _0161_, _0160_, _0159_, _0158_, _0157_, _0156_, _0155_, _0154_, _0153_, _0152_, _0151_, _0150_, _0149_, _0148_, _0147_, _0146_, _0145_, _0144_, _0143_, _0142_, _0141_, _0140_, _0139_, _0138_, _0137_, _0136_, _0135_, _0134_, _0133_, _0132_, _0131_, _0130_, _0129_, _0128_, _0127_, _0126_, _0125_, _0124_, _0123_, _0122_, _0121_, _0120_, _0119_, _0118_, _0117_, _0116_, _0115_, _0114_, _0113_, _0112_, _0111_, _0110_, _0109_, _0108_, _0107_, _0106_, _0105_, _0104_, _0103_, _0102_, _0101_, _0100_, _0099_, _0098_, _0097_, _0096_, _0095_, _0094_, _0093_, _0092_, _0091_, _0090_, _0089_, _0088_, _0087_, _0086_, _0085_, _0084_, _0083_, _0082_, _0081_, _0080_, _0079_, _0078_, _0077_, _0076_, _0075_, _0074_, _0073_, _0072_, _0071_, _0070_, _0069_, _0068_, _0067_, _0066_, _0065_, _0064_, _0063_, _0062_, _0061_, _0060_, _0059_, _0058_, _0057_, _0056_, _0055_, _0054_, _0053_, _0052_, _0051_, _0050_, _0049_, _0048_, _0047_, _0046_, _0045_, _0044_, _0043_, _0042_, _0041_, _0040_, _0039_, _0038_, _0037_, _0036_, _0035_, _0034_, _0033_, _0032_, _0031_, _0030_, _0029_, _0028_, _0027_, _0026_, _0025_, _0024_, _0023_, _0022_, _0021_, _0020_, _0019_, _0018_, _0017_, _0016_, _0015_, _0014_, _0013_, _0012_, _0011_, _0010_, _0009_, _0008_, _0007_, _0006_, _0005_, _0004_, _0003_, _0002_, _0001_ };

  always @(\t0.t0.s4.out or fangyuan2) begin
    casez (fangyuan2)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0257_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0257_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0257_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0257_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0257_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0257_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0257_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0257_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0257_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0257_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0257_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0257_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0257_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0257_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0257_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0257_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0257_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0257_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0257_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0257_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0257_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0257_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0257_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0257_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0257_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0257_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0257_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0257_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0257_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0257_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0257_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0257_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0257_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0257_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0257_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0257_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0257_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0257_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0257_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0257_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0257_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0257_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0257_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0257_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0257_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0257_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0257_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0257_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0257_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0257_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0257_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0257_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0257_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0257_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0257_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0257_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0257_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0257_ = 8'b11000110 ;
      default:
        _0257_ = \t0.t0.s4.out ;
    endcase
  end
  assign p01[31:24] = \t0.t1.s0.out ^ \t0.t1.s4.out ;
  always @(posedge clk)
      \t0.t1.s0.out <= _0258_;
  logic [255:0] fangyuan3;
  assign fangyuan3 = { _0514_, _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0430_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0419_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0397_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0309_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0298_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_, _0290_, _0289_, _0288_, _0287_, _0286_, _0285_, _0284_, _0283_, _0282_, _0281_, _0280_, _0279_, _0278_, _0277_, _0276_, _0275_, _0274_, _0273_, _0272_, _0271_, _0270_, _0269_, _0268_, _0267_, _0266_, _0265_, _0264_, _0263_, _0262_, _0261_, _0260_, _0259_ };

  always @(\t0.t1.s0.out or fangyuan3) begin
    casez (fangyuan3)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0258_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0258_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0258_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0258_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0258_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0258_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0258_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0258_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0258_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0258_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0258_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0258_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0258_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0258_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0258_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0258_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0258_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0258_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0258_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0258_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0258_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0258_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0258_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0258_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0258_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0258_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0258_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0258_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0258_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0258_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0258_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0258_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0258_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0258_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0258_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0258_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0258_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0258_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0258_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0258_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0258_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0258_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0258_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0258_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0258_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0258_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0258_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0258_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0258_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0258_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0258_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0258_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0258_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0258_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0258_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0258_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0258_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0258_ = 8'b01100011 ;
      default:
        _0258_ = \t0.t1.s0.out ;
    endcase
  end
  assign _0259_ = state_in[119:112] == 8'b11111111;
  assign _0260_ = state_in[119:112] == 8'b11111110;
  assign _0261_ = state_in[119:112] == 8'b11111101;
  assign _0262_ = state_in[119:112] == 8'b11111100;
  assign _0263_ = state_in[119:112] == 8'b11111011;
  assign _0264_ = state_in[119:112] == 8'b11111010;
  assign _0265_ = state_in[119:112] == 8'b11111001;
  assign _0266_ = state_in[119:112] == 8'b11111000;
  assign _0267_ = state_in[119:112] == 8'b11110111;
  assign _0268_ = state_in[119:112] == 8'b11110110;
  assign _0269_ = state_in[119:112] == 8'b11110101;
  assign _0270_ = state_in[119:112] == 8'b11110100;
  assign _0271_ = state_in[119:112] == 8'b11110011;
  assign _0272_ = state_in[119:112] == 8'b11110010;
  assign _0273_ = state_in[119:112] == 8'b11110001;
  assign _0274_ = state_in[119:112] == 8'b11110000;
  assign _0275_ = state_in[119:112] == 8'b11101111;
  assign _0276_ = state_in[119:112] == 8'b11101110;
  assign _0277_ = state_in[119:112] == 8'b11101101;
  assign _0278_ = state_in[119:112] == 8'b11101100;
  assign _0279_ = state_in[119:112] == 8'b11101011;
  assign _0280_ = state_in[119:112] == 8'b11101010;
  assign _0281_ = state_in[119:112] == 8'b11101001;
  assign _0282_ = state_in[119:112] == 8'b11101000;
  assign _0283_ = state_in[119:112] == 8'b11100111;
  assign _0284_ = state_in[119:112] == 8'b11100110;
  assign _0285_ = state_in[119:112] == 8'b11100101;
  assign _0286_ = state_in[119:112] == 8'b11100100;
  assign _0287_ = state_in[119:112] == 8'b11100011;
  assign _0288_ = state_in[119:112] == 8'b11100010;
  assign _0289_ = state_in[119:112] == 8'b11100001;
  assign _0290_ = state_in[119:112] == 8'b11100000;
  assign _0291_ = state_in[119:112] == 8'b11011111;
  assign _0292_ = state_in[119:112] == 8'b11011110;
  assign _0293_ = state_in[119:112] == 8'b11011101;
  assign _0294_ = state_in[119:112] == 8'b11011100;
  assign _0295_ = state_in[119:112] == 8'b11011011;
  assign _0296_ = state_in[119:112] == 8'b11011010;
  assign _0297_ = state_in[119:112] == 8'b11011001;
  assign _0298_ = state_in[119:112] == 8'b11011000;
  assign _0299_ = state_in[119:112] == 8'b11010111;
  assign _0300_ = state_in[119:112] == 8'b11010110;
  assign _0301_ = state_in[119:112] == 8'b11010101;
  assign _0302_ = state_in[119:112] == 8'b11010100;
  assign _0303_ = state_in[119:112] == 8'b11010011;
  assign _0304_ = state_in[119:112] == 8'b11010010;
  assign _0305_ = state_in[119:112] == 8'b11010001;
  assign _0306_ = state_in[119:112] == 8'b11010000;
  assign _0307_ = state_in[119:112] == 8'b11001111;
  assign _0308_ = state_in[119:112] == 8'b11001110;
  assign _0309_ = state_in[119:112] == 8'b11001101;
  assign _0310_ = state_in[119:112] == 8'b11001100;
  assign _0311_ = state_in[119:112] == 8'b11001011;
  assign _0312_ = state_in[119:112] == 8'b11001010;
  assign _0313_ = state_in[119:112] == 8'b11001001;
  assign _0314_ = state_in[119:112] == 8'b11001000;
  assign _0315_ = state_in[119:112] == 8'b11000111;
  assign _0316_ = state_in[119:112] == 8'b11000110;
  assign _0317_ = state_in[119:112] == 8'b11000101;
  assign _0318_ = state_in[119:112] == 8'b11000100;
  assign _0319_ = state_in[119:112] == 8'b11000011;
  assign _0320_ = state_in[119:112] == 8'b11000010;
  assign _0321_ = state_in[119:112] == 8'b11000001;
  assign _0322_ = state_in[119:112] == 8'b11000000;
  assign _0323_ = state_in[119:112] == 8'b10111111;
  assign _0324_ = state_in[119:112] == 8'b10111110;
  assign _0325_ = state_in[119:112] == 8'b10111101;
  assign _0326_ = state_in[119:112] == 8'b10111100;
  assign _0327_ = state_in[119:112] == 8'b10111011;
  assign _0328_ = state_in[119:112] == 8'b10111010;
  assign _0329_ = state_in[119:112] == 8'b10111001;
  assign _0330_ = state_in[119:112] == 8'b10111000;
  assign _0331_ = state_in[119:112] == 8'b10110111;
  assign _0332_ = state_in[119:112] == 8'b10110110;
  assign _0333_ = state_in[119:112] == 8'b10110101;
  assign _0334_ = state_in[119:112] == 8'b10110100;
  assign _0335_ = state_in[119:112] == 8'b10110011;
  assign _0336_ = state_in[119:112] == 8'b10110010;
  assign _0337_ = state_in[119:112] == 8'b10110001;
  assign _0338_ = state_in[119:112] == 8'b10110000;
  assign _0339_ = state_in[119:112] == 8'b10101111;
  assign _0340_ = state_in[119:112] == 8'b10101110;
  assign _0341_ = state_in[119:112] == 8'b10101101;
  assign _0342_ = state_in[119:112] == 8'b10101100;
  assign _0343_ = state_in[119:112] == 8'b10101011;
  assign _0344_ = state_in[119:112] == 8'b10101010;
  assign _0345_ = state_in[119:112] == 8'b10101001;
  assign _0346_ = state_in[119:112] == 8'b10101000;
  assign _0347_ = state_in[119:112] == 8'b10100111;
  assign _0348_ = state_in[119:112] == 8'b10100110;
  assign _0349_ = state_in[119:112] == 8'b10100101;
  assign _0350_ = state_in[119:112] == 8'b10100100;
  assign _0351_ = state_in[119:112] == 8'b10100011;
  assign _0352_ = state_in[119:112] == 8'b10100010;
  assign _0353_ = state_in[119:112] == 8'b10100001;
  assign _0354_ = state_in[119:112] == 8'b10100000;
  assign _0355_ = state_in[119:112] == 8'b10011111;
  assign _0356_ = state_in[119:112] == 8'b10011110;
  assign _0357_ = state_in[119:112] == 8'b10011101;
  assign _0358_ = state_in[119:112] == 8'b10011100;
  assign _0359_ = state_in[119:112] == 8'b10011011;
  assign _0360_ = state_in[119:112] == 8'b10011010;
  assign _0361_ = state_in[119:112] == 8'b10011001;
  assign _0362_ = state_in[119:112] == 8'b10011000;
  assign _0363_ = state_in[119:112] == 8'b10010111;
  assign _0364_ = state_in[119:112] == 8'b10010110;
  assign _0365_ = state_in[119:112] == 8'b10010101;
  assign _0366_ = state_in[119:112] == 8'b10010100;
  assign _0367_ = state_in[119:112] == 8'b10010011;
  assign _0368_ = state_in[119:112] == 8'b10010010;
  assign _0369_ = state_in[119:112] == 8'b10010001;
  assign _0370_ = state_in[119:112] == 8'b10010000;
  assign _0371_ = state_in[119:112] == 8'b10001111;
  assign _0372_ = state_in[119:112] == 8'b10001110;
  assign _0373_ = state_in[119:112] == 8'b10001101;
  assign _0374_ = state_in[119:112] == 8'b10001100;
  assign _0375_ = state_in[119:112] == 8'b10001011;
  assign _0376_ = state_in[119:112] == 8'b10001010;
  assign _0377_ = state_in[119:112] == 8'b10001001;
  assign _0378_ = state_in[119:112] == 8'b10001000;
  assign _0379_ = state_in[119:112] == 8'b10000111;
  assign _0380_ = state_in[119:112] == 8'b10000110;
  assign _0381_ = state_in[119:112] == 8'b10000101;
  assign _0382_ = state_in[119:112] == 8'b10000100;
  assign _0383_ = state_in[119:112] == 8'b10000011;
  assign _0384_ = state_in[119:112] == 8'b10000010;
  assign _0385_ = state_in[119:112] == 8'b10000001;
  assign _0386_ = state_in[119:112] == 8'b10000000;
  assign _0387_ = state_in[119:112] == 7'b1111111;
  assign _0388_ = state_in[119:112] == 7'b1111110;
  assign _0389_ = state_in[119:112] == 7'b1111101;
  assign _0390_ = state_in[119:112] == 7'b1111100;
  assign _0391_ = state_in[119:112] == 7'b1111011;
  assign _0392_ = state_in[119:112] == 7'b1111010;
  assign _0393_ = state_in[119:112] == 7'b1111001;
  assign _0394_ = state_in[119:112] == 7'b1111000;
  assign _0395_ = state_in[119:112] == 7'b1110111;
  assign _0396_ = state_in[119:112] == 7'b1110110;
  assign _0397_ = state_in[119:112] == 7'b1110101;
  assign _0398_ = state_in[119:112] == 7'b1110100;
  assign _0399_ = state_in[119:112] == 7'b1110011;
  assign _0400_ = state_in[119:112] == 7'b1110010;
  assign _0401_ = state_in[119:112] == 7'b1110001;
  assign _0402_ = state_in[119:112] == 7'b1110000;
  assign _0403_ = state_in[119:112] == 7'b1101111;
  assign _0404_ = state_in[119:112] == 7'b1101110;
  assign _0405_ = state_in[119:112] == 7'b1101101;
  assign _0406_ = state_in[119:112] == 7'b1101100;
  assign _0407_ = state_in[119:112] == 7'b1101011;
  assign _0408_ = state_in[119:112] == 7'b1101010;
  assign _0409_ = state_in[119:112] == 7'b1101001;
  assign _0410_ = state_in[119:112] == 7'b1101000;
  assign _0411_ = state_in[119:112] == 7'b1100111;
  assign _0412_ = state_in[119:112] == 7'b1100110;
  assign _0413_ = state_in[119:112] == 7'b1100101;
  assign _0414_ = state_in[119:112] == 7'b1100100;
  assign _0415_ = state_in[119:112] == 7'b1100011;
  assign _0416_ = state_in[119:112] == 7'b1100010;
  assign _0417_ = state_in[119:112] == 7'b1100001;
  assign _0418_ = state_in[119:112] == 7'b1100000;
  assign _0419_ = state_in[119:112] == 7'b1011111;
  assign _0420_ = state_in[119:112] == 7'b1011110;
  assign _0421_ = state_in[119:112] == 7'b1011101;
  assign _0422_ = state_in[119:112] == 7'b1011100;
  assign _0423_ = state_in[119:112] == 7'b1011011;
  assign _0424_ = state_in[119:112] == 7'b1011010;
  assign _0425_ = state_in[119:112] == 7'b1011001;
  assign _0426_ = state_in[119:112] == 7'b1011000;
  assign _0427_ = state_in[119:112] == 7'b1010111;
  assign _0428_ = state_in[119:112] == 7'b1010110;
  assign _0429_ = state_in[119:112] == 7'b1010101;
  assign _0430_ = state_in[119:112] == 7'b1010100;
  assign _0431_ = state_in[119:112] == 7'b1010011;
  assign _0432_ = state_in[119:112] == 7'b1010010;
  assign _0433_ = state_in[119:112] == 7'b1010001;
  assign _0434_ = state_in[119:112] == 7'b1010000;
  assign _0435_ = state_in[119:112] == 7'b1001111;
  assign _0436_ = state_in[119:112] == 7'b1001110;
  assign _0437_ = state_in[119:112] == 7'b1001101;
  assign _0438_ = state_in[119:112] == 7'b1001100;
  assign _0439_ = state_in[119:112] == 7'b1001011;
  assign _0440_ = state_in[119:112] == 7'b1001010;
  assign _0441_ = state_in[119:112] == 7'b1001001;
  assign _0442_ = state_in[119:112] == 7'b1001000;
  assign _0443_ = state_in[119:112] == 7'b1000111;
  assign _0444_ = state_in[119:112] == 7'b1000110;
  assign _0445_ = state_in[119:112] == 7'b1000101;
  assign _0446_ = state_in[119:112] == 7'b1000100;
  assign _0447_ = state_in[119:112] == 7'b1000011;
  assign _0448_ = state_in[119:112] == 7'b1000010;
  assign _0449_ = state_in[119:112] == 7'b1000001;
  assign _0450_ = state_in[119:112] == 7'b1000000;
  assign _0451_ = state_in[119:112] == 6'b111111;
  assign _0452_ = state_in[119:112] == 6'b111110;
  assign _0453_ = state_in[119:112] == 6'b111101;
  assign _0454_ = state_in[119:112] == 6'b111100;
  assign _0455_ = state_in[119:112] == 6'b111011;
  assign _0456_ = state_in[119:112] == 6'b111010;
  assign _0457_ = state_in[119:112] == 6'b111001;
  assign _0458_ = state_in[119:112] == 6'b111000;
  assign _0459_ = state_in[119:112] == 6'b110111;
  assign _0460_ = state_in[119:112] == 6'b110110;
  assign _0461_ = state_in[119:112] == 6'b110101;
  assign _0462_ = state_in[119:112] == 6'b110100;
  assign _0463_ = state_in[119:112] == 6'b110011;
  assign _0464_ = state_in[119:112] == 6'b110010;
  assign _0465_ = state_in[119:112] == 6'b110001;
  assign _0466_ = state_in[119:112] == 6'b110000;
  assign _0467_ = state_in[119:112] == 6'b101111;
  assign _0468_ = state_in[119:112] == 6'b101110;
  assign _0469_ = state_in[119:112] == 6'b101101;
  assign _0470_ = state_in[119:112] == 6'b101100;
  assign _0471_ = state_in[119:112] == 6'b101011;
  assign _0472_ = state_in[119:112] == 6'b101010;
  assign _0473_ = state_in[119:112] == 6'b101001;
  assign _0474_ = state_in[119:112] == 6'b101000;
  assign _0475_ = state_in[119:112] == 6'b100111;
  assign _0476_ = state_in[119:112] == 6'b100110;
  assign _0477_ = state_in[119:112] == 6'b100101;
  assign _0478_ = state_in[119:112] == 6'b100100;
  assign _0479_ = state_in[119:112] == 6'b100011;
  assign _0480_ = state_in[119:112] == 6'b100010;
  assign _0481_ = state_in[119:112] == 6'b100001;
  assign _0482_ = state_in[119:112] == 6'b100000;
  assign _0483_ = state_in[119:112] == 5'b11111;
  assign _0484_ = state_in[119:112] == 5'b11110;
  assign _0485_ = state_in[119:112] == 5'b11101;
  assign _0486_ = state_in[119:112] == 5'b11100;
  assign _0487_ = state_in[119:112] == 5'b11011;
  assign _0488_ = state_in[119:112] == 5'b11010;
  assign _0489_ = state_in[119:112] == 5'b11001;
  assign _0490_ = state_in[119:112] == 5'b11000;
  assign _0491_ = state_in[119:112] == 5'b10111;
  assign _0492_ = state_in[119:112] == 5'b10110;
  assign _0493_ = state_in[119:112] == 5'b10101;
  assign _0494_ = state_in[119:112] == 5'b10100;
  assign _0495_ = state_in[119:112] == 5'b10011;
  assign _0496_ = state_in[119:112] == 5'b10010;
  assign _0497_ = state_in[119:112] == 5'b10001;
  assign _0498_ = state_in[119:112] == 5'b10000;
  assign _0499_ = state_in[119:112] == 4'b1111;
  assign _0500_ = state_in[119:112] == 4'b1110;
  assign _0501_ = state_in[119:112] == 4'b1101;
  assign _0502_ = state_in[119:112] == 4'b1100;
  assign _0503_ = state_in[119:112] == 4'b1011;
  assign _0504_ = state_in[119:112] == 4'b1010;
  assign _0505_ = state_in[119:112] == 4'b1001;
  assign _0506_ = state_in[119:112] == 4'b1000;
  assign _0507_ = state_in[119:112] == 3'b111;
  assign _0508_ = state_in[119:112] == 3'b110;
  assign _0509_ = state_in[119:112] == 3'b101;
  assign _0510_ = state_in[119:112] == 3'b100;
  assign _0511_ = state_in[119:112] == 2'b11;
  assign _0512_ = state_in[119:112] == 2'b10;
  assign _0513_ = state_in[119:112] == 1'b1;
  assign _0514_ = ! state_in[119:112];
  always @(posedge clk)
      \t0.t1.s4.out <= _0515_;
  logic [255:0] fangyuan4;
  assign fangyuan4 = { _0514_, _0513_, _0512_, _0511_, _0510_, _0509_, _0508_, _0507_, _0506_, _0505_, _0504_, _0503_, _0502_, _0501_, _0500_, _0499_, _0498_, _0497_, _0496_, _0495_, _0494_, _0493_, _0492_, _0491_, _0490_, _0489_, _0488_, _0487_, _0486_, _0485_, _0484_, _0483_, _0482_, _0481_, _0480_, _0479_, _0478_, _0477_, _0476_, _0475_, _0474_, _0473_, _0472_, _0471_, _0470_, _0469_, _0468_, _0467_, _0466_, _0465_, _0464_, _0463_, _0462_, _0461_, _0460_, _0459_, _0458_, _0457_, _0456_, _0455_, _0454_, _0453_, _0452_, _0451_, _0450_, _0449_, _0448_, _0447_, _0446_, _0445_, _0444_, _0443_, _0442_, _0441_, _0440_, _0439_, _0438_, _0437_, _0436_, _0435_, _0434_, _0433_, _0432_, _0431_, _0430_, _0429_, _0428_, _0427_, _0426_, _0425_, _0424_, _0423_, _0422_, _0421_, _0420_, _0419_, _0418_, _0417_, _0416_, _0415_, _0414_, _0413_, _0412_, _0411_, _0410_, _0409_, _0408_, _0407_, _0406_, _0405_, _0404_, _0403_, _0402_, _0401_, _0400_, _0399_, _0398_, _0397_, _0396_, _0395_, _0394_, _0393_, _0392_, _0391_, _0390_, _0389_, _0388_, _0387_, _0386_, _0385_, _0384_, _0383_, _0382_, _0381_, _0380_, _0379_, _0378_, _0377_, _0376_, _0375_, _0374_, _0373_, _0372_, _0371_, _0370_, _0369_, _0368_, _0367_, _0366_, _0365_, _0364_, _0363_, _0362_, _0361_, _0360_, _0359_, _0358_, _0357_, _0356_, _0355_, _0354_, _0353_, _0352_, _0351_, _0350_, _0349_, _0348_, _0347_, _0346_, _0345_, _0344_, _0343_, _0342_, _0341_, _0340_, _0339_, _0338_, _0337_, _0336_, _0335_, _0334_, _0333_, _0332_, _0331_, _0330_, _0329_, _0328_, _0327_, _0326_, _0325_, _0324_, _0323_, _0322_, _0321_, _0320_, _0319_, _0318_, _0317_, _0316_, _0315_, _0314_, _0313_, _0312_, _0311_, _0310_, _0309_, _0308_, _0307_, _0306_, _0305_, _0304_, _0303_, _0302_, _0301_, _0300_, _0299_, _0298_, _0297_, _0296_, _0295_, _0294_, _0293_, _0292_, _0291_, _0290_, _0289_, _0288_, _0287_, _0286_, _0285_, _0284_, _0283_, _0282_, _0281_, _0280_, _0279_, _0278_, _0277_, _0276_, _0275_, _0274_, _0273_, _0272_, _0271_, _0270_, _0269_, _0268_, _0267_, _0266_, _0265_, _0264_, _0263_, _0262_, _0261_, _0260_, _0259_ };

  always @(\t0.t1.s4.out or fangyuan4) begin
    casez (fangyuan4)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0515_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0515_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0515_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0515_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0515_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0515_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0515_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0515_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0515_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0515_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0515_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0515_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0515_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0515_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0515_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0515_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0515_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0515_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0515_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0515_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0515_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0515_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0515_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0515_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0515_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0515_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0515_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0515_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0515_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0515_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0515_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0515_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0515_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0515_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0515_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0515_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0515_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0515_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0515_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0515_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0515_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0515_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0515_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0515_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0515_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0515_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0515_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0515_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0515_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0515_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0515_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0515_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0515_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0515_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0515_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0515_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0515_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0515_ = 8'b11000110 ;
      default:
        _0515_ = \t0.t1.s4.out ;
    endcase
  end
  assign p02[23:16] = \t0.t2.s0.out ^ \t0.t2.s4.out ;
  always @(posedge clk)
      \t0.t2.s0.out <= _0516_;
  logic [255:0] fangyuan5;
  assign fangyuan5 = { _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0676_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0665_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_, _0656_, _0655_, _0654_, _0653_, _0652_, _0651_, _0650_, _0649_, _0648_, _0647_, _0646_, _0645_, _0644_, _0643_, _0642_, _0641_, _0640_, _0639_, _0638_, _0637_, _0636_, _0635_, _0634_, _0633_, _0632_, _0631_, _0630_, _0629_, _0628_, _0627_, _0626_, _0625_, _0624_, _0623_, _0622_, _0621_, _0620_, _0619_, _0618_, _0617_, _0616_, _0615_, _0614_, _0613_, _0612_, _0611_, _0610_, _0609_, _0608_, _0607_, _0606_, _0605_, _0604_, _0603_, _0602_, _0601_, _0600_, _0599_, _0598_, _0597_, _0596_, _0595_, _0594_, _0593_, _0592_, _0591_, _0590_, _0589_, _0588_, _0587_, _0586_, _0585_, _0584_, _0583_, _0582_, _0581_, _0580_, _0579_, _0578_, _0577_, _0576_, _0575_, _0574_, _0573_, _0572_, _0571_, _0570_, _0569_, _0568_, _0567_, _0566_, _0565_, _0564_, _0563_, _0562_, _0561_, _0560_, _0559_, _0558_, _0557_, _0556_, _0555_, _0554_, _0553_, _0552_, _0551_, _0550_, _0549_, _0548_, _0547_, _0546_, _0545_, _0544_, _0543_, _0542_, _0541_, _0540_, _0539_, _0538_, _0537_, _0536_, _0535_, _0534_, _0533_, _0532_, _0531_, _0530_, _0529_, _0528_, _0527_, _0526_, _0525_, _0524_, _0523_, _0522_, _0521_, _0520_, _0519_, _0518_, _0517_ };

  always @(\t0.t2.s0.out or fangyuan5) begin
    casez (fangyuan5)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0516_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0516_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0516_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0516_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0516_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0516_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0516_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0516_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0516_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0516_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0516_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0516_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0516_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0516_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0516_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0516_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0516_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0516_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0516_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0516_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0516_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0516_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0516_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0516_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0516_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0516_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0516_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0516_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0516_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0516_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0516_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0516_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0516_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0516_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0516_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0516_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0516_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0516_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0516_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0516_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0516_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0516_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0516_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0516_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0516_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0516_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0516_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0516_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0516_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0516_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0516_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0516_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0516_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0516_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0516_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0516_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0516_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0516_ = 8'b01100011 ;
      default:
        _0516_ = \t0.t2.s0.out ;
    endcase
  end
  assign _0517_ = state_in[111:104] == 8'b11111111;
  assign _0518_ = state_in[111:104] == 8'b11111110;
  assign _0519_ = state_in[111:104] == 8'b11111101;
  assign _0520_ = state_in[111:104] == 8'b11111100;
  assign _0521_ = state_in[111:104] == 8'b11111011;
  assign _0522_ = state_in[111:104] == 8'b11111010;
  assign _0523_ = state_in[111:104] == 8'b11111001;
  assign _0524_ = state_in[111:104] == 8'b11111000;
  assign _0525_ = state_in[111:104] == 8'b11110111;
  assign _0526_ = state_in[111:104] == 8'b11110110;
  assign _0527_ = state_in[111:104] == 8'b11110101;
  assign _0528_ = state_in[111:104] == 8'b11110100;
  assign _0529_ = state_in[111:104] == 8'b11110011;
  assign _0530_ = state_in[111:104] == 8'b11110010;
  assign _0531_ = state_in[111:104] == 8'b11110001;
  assign _0532_ = state_in[111:104] == 8'b11110000;
  assign _0533_ = state_in[111:104] == 8'b11101111;
  assign _0534_ = state_in[111:104] == 8'b11101110;
  assign _0535_ = state_in[111:104] == 8'b11101101;
  assign _0536_ = state_in[111:104] == 8'b11101100;
  assign _0537_ = state_in[111:104] == 8'b11101011;
  assign _0538_ = state_in[111:104] == 8'b11101010;
  assign _0539_ = state_in[111:104] == 8'b11101001;
  assign _0540_ = state_in[111:104] == 8'b11101000;
  assign _0541_ = state_in[111:104] == 8'b11100111;
  assign _0542_ = state_in[111:104] == 8'b11100110;
  assign _0543_ = state_in[111:104] == 8'b11100101;
  assign _0544_ = state_in[111:104] == 8'b11100100;
  assign _0545_ = state_in[111:104] == 8'b11100011;
  assign _0546_ = state_in[111:104] == 8'b11100010;
  assign _0547_ = state_in[111:104] == 8'b11100001;
  assign _0548_ = state_in[111:104] == 8'b11100000;
  assign _0549_ = state_in[111:104] == 8'b11011111;
  assign _0550_ = state_in[111:104] == 8'b11011110;
  assign _0551_ = state_in[111:104] == 8'b11011101;
  assign _0552_ = state_in[111:104] == 8'b11011100;
  assign _0553_ = state_in[111:104] == 8'b11011011;
  assign _0554_ = state_in[111:104] == 8'b11011010;
  assign _0555_ = state_in[111:104] == 8'b11011001;
  assign _0556_ = state_in[111:104] == 8'b11011000;
  assign _0557_ = state_in[111:104] == 8'b11010111;
  assign _0558_ = state_in[111:104] == 8'b11010110;
  assign _0559_ = state_in[111:104] == 8'b11010101;
  assign _0560_ = state_in[111:104] == 8'b11010100;
  assign _0561_ = state_in[111:104] == 8'b11010011;
  assign _0562_ = state_in[111:104] == 8'b11010010;
  assign _0563_ = state_in[111:104] == 8'b11010001;
  assign _0564_ = state_in[111:104] == 8'b11010000;
  assign _0565_ = state_in[111:104] == 8'b11001111;
  assign _0566_ = state_in[111:104] == 8'b11001110;
  assign _0567_ = state_in[111:104] == 8'b11001101;
  assign _0568_ = state_in[111:104] == 8'b11001100;
  assign _0569_ = state_in[111:104] == 8'b11001011;
  assign _0570_ = state_in[111:104] == 8'b11001010;
  assign _0571_ = state_in[111:104] == 8'b11001001;
  assign _0572_ = state_in[111:104] == 8'b11001000;
  assign _0573_ = state_in[111:104] == 8'b11000111;
  assign _0574_ = state_in[111:104] == 8'b11000110;
  assign _0575_ = state_in[111:104] == 8'b11000101;
  assign _0576_ = state_in[111:104] == 8'b11000100;
  assign _0577_ = state_in[111:104] == 8'b11000011;
  assign _0578_ = state_in[111:104] == 8'b11000010;
  assign _0579_ = state_in[111:104] == 8'b11000001;
  assign _0580_ = state_in[111:104] == 8'b11000000;
  assign _0581_ = state_in[111:104] == 8'b10111111;
  assign _0582_ = state_in[111:104] == 8'b10111110;
  assign _0583_ = state_in[111:104] == 8'b10111101;
  assign _0584_ = state_in[111:104] == 8'b10111100;
  assign _0585_ = state_in[111:104] == 8'b10111011;
  assign _0586_ = state_in[111:104] == 8'b10111010;
  assign _0587_ = state_in[111:104] == 8'b10111001;
  assign _0588_ = state_in[111:104] == 8'b10111000;
  assign _0589_ = state_in[111:104] == 8'b10110111;
  assign _0590_ = state_in[111:104] == 8'b10110110;
  assign _0591_ = state_in[111:104] == 8'b10110101;
  assign _0592_ = state_in[111:104] == 8'b10110100;
  assign _0593_ = state_in[111:104] == 8'b10110011;
  assign _0594_ = state_in[111:104] == 8'b10110010;
  assign _0595_ = state_in[111:104] == 8'b10110001;
  assign _0596_ = state_in[111:104] == 8'b10110000;
  assign _0597_ = state_in[111:104] == 8'b10101111;
  assign _0598_ = state_in[111:104] == 8'b10101110;
  assign _0599_ = state_in[111:104] == 8'b10101101;
  assign _0600_ = state_in[111:104] == 8'b10101100;
  assign _0601_ = state_in[111:104] == 8'b10101011;
  assign _0602_ = state_in[111:104] == 8'b10101010;
  assign _0603_ = state_in[111:104] == 8'b10101001;
  assign _0604_ = state_in[111:104] == 8'b10101000;
  assign _0605_ = state_in[111:104] == 8'b10100111;
  assign _0606_ = state_in[111:104] == 8'b10100110;
  assign _0607_ = state_in[111:104] == 8'b10100101;
  assign _0608_ = state_in[111:104] == 8'b10100100;
  assign _0609_ = state_in[111:104] == 8'b10100011;
  assign _0610_ = state_in[111:104] == 8'b10100010;
  assign _0611_ = state_in[111:104] == 8'b10100001;
  assign _0612_ = state_in[111:104] == 8'b10100000;
  assign _0613_ = state_in[111:104] == 8'b10011111;
  assign _0614_ = state_in[111:104] == 8'b10011110;
  assign _0615_ = state_in[111:104] == 8'b10011101;
  assign _0616_ = state_in[111:104] == 8'b10011100;
  assign _0617_ = state_in[111:104] == 8'b10011011;
  assign _0618_ = state_in[111:104] == 8'b10011010;
  assign _0619_ = state_in[111:104] == 8'b10011001;
  assign _0620_ = state_in[111:104] == 8'b10011000;
  assign _0621_ = state_in[111:104] == 8'b10010111;
  assign _0622_ = state_in[111:104] == 8'b10010110;
  assign _0623_ = state_in[111:104] == 8'b10010101;
  assign _0624_ = state_in[111:104] == 8'b10010100;
  assign _0625_ = state_in[111:104] == 8'b10010011;
  assign _0626_ = state_in[111:104] == 8'b10010010;
  assign _0627_ = state_in[111:104] == 8'b10010001;
  assign _0628_ = state_in[111:104] == 8'b10010000;
  assign _0629_ = state_in[111:104] == 8'b10001111;
  assign _0630_ = state_in[111:104] == 8'b10001110;
  assign _0631_ = state_in[111:104] == 8'b10001101;
  assign _0632_ = state_in[111:104] == 8'b10001100;
  assign _0633_ = state_in[111:104] == 8'b10001011;
  assign _0634_ = state_in[111:104] == 8'b10001010;
  assign _0635_ = state_in[111:104] == 8'b10001001;
  assign _0636_ = state_in[111:104] == 8'b10001000;
  assign _0637_ = state_in[111:104] == 8'b10000111;
  assign _0638_ = state_in[111:104] == 8'b10000110;
  assign _0639_ = state_in[111:104] == 8'b10000101;
  assign _0640_ = state_in[111:104] == 8'b10000100;
  assign _0641_ = state_in[111:104] == 8'b10000011;
  assign _0642_ = state_in[111:104] == 8'b10000010;
  assign _0643_ = state_in[111:104] == 8'b10000001;
  assign _0644_ = state_in[111:104] == 8'b10000000;
  assign _0645_ = state_in[111:104] == 7'b1111111;
  assign _0646_ = state_in[111:104] == 7'b1111110;
  assign _0647_ = state_in[111:104] == 7'b1111101;
  assign _0648_ = state_in[111:104] == 7'b1111100;
  assign _0649_ = state_in[111:104] == 7'b1111011;
  assign _0650_ = state_in[111:104] == 7'b1111010;
  assign _0651_ = state_in[111:104] == 7'b1111001;
  assign _0652_ = state_in[111:104] == 7'b1111000;
  assign _0653_ = state_in[111:104] == 7'b1110111;
  assign _0654_ = state_in[111:104] == 7'b1110110;
  assign _0655_ = state_in[111:104] == 7'b1110101;
  assign _0656_ = state_in[111:104] == 7'b1110100;
  assign _0657_ = state_in[111:104] == 7'b1110011;
  assign _0658_ = state_in[111:104] == 7'b1110010;
  assign _0659_ = state_in[111:104] == 7'b1110001;
  assign _0660_ = state_in[111:104] == 7'b1110000;
  assign _0661_ = state_in[111:104] == 7'b1101111;
  assign _0662_ = state_in[111:104] == 7'b1101110;
  assign _0663_ = state_in[111:104] == 7'b1101101;
  assign _0664_ = state_in[111:104] == 7'b1101100;
  assign _0665_ = state_in[111:104] == 7'b1101011;
  assign _0666_ = state_in[111:104] == 7'b1101010;
  assign _0667_ = state_in[111:104] == 7'b1101001;
  assign _0668_ = state_in[111:104] == 7'b1101000;
  assign _0669_ = state_in[111:104] == 7'b1100111;
  assign _0670_ = state_in[111:104] == 7'b1100110;
  assign _0671_ = state_in[111:104] == 7'b1100101;
  assign _0672_ = state_in[111:104] == 7'b1100100;
  assign _0673_ = state_in[111:104] == 7'b1100011;
  assign _0674_ = state_in[111:104] == 7'b1100010;
  assign _0675_ = state_in[111:104] == 7'b1100001;
  assign _0676_ = state_in[111:104] == 7'b1100000;
  assign _0677_ = state_in[111:104] == 7'b1011111;
  assign _0678_ = state_in[111:104] == 7'b1011110;
  assign _0679_ = state_in[111:104] == 7'b1011101;
  assign _0680_ = state_in[111:104] == 7'b1011100;
  assign _0681_ = state_in[111:104] == 7'b1011011;
  assign _0682_ = state_in[111:104] == 7'b1011010;
  assign _0683_ = state_in[111:104] == 7'b1011001;
  assign _0684_ = state_in[111:104] == 7'b1011000;
  assign _0685_ = state_in[111:104] == 7'b1010111;
  assign _0686_ = state_in[111:104] == 7'b1010110;
  assign _0687_ = state_in[111:104] == 7'b1010101;
  assign _0688_ = state_in[111:104] == 7'b1010100;
  assign _0689_ = state_in[111:104] == 7'b1010011;
  assign _0690_ = state_in[111:104] == 7'b1010010;
  assign _0691_ = state_in[111:104] == 7'b1010001;
  assign _0692_ = state_in[111:104] == 7'b1010000;
  assign _0693_ = state_in[111:104] == 7'b1001111;
  assign _0694_ = state_in[111:104] == 7'b1001110;
  assign _0695_ = state_in[111:104] == 7'b1001101;
  assign _0696_ = state_in[111:104] == 7'b1001100;
  assign _0697_ = state_in[111:104] == 7'b1001011;
  assign _0698_ = state_in[111:104] == 7'b1001010;
  assign _0699_ = state_in[111:104] == 7'b1001001;
  assign _0700_ = state_in[111:104] == 7'b1001000;
  assign _0701_ = state_in[111:104] == 7'b1000111;
  assign _0702_ = state_in[111:104] == 7'b1000110;
  assign _0703_ = state_in[111:104] == 7'b1000101;
  assign _0704_ = state_in[111:104] == 7'b1000100;
  assign _0705_ = state_in[111:104] == 7'b1000011;
  assign _0706_ = state_in[111:104] == 7'b1000010;
  assign _0707_ = state_in[111:104] == 7'b1000001;
  assign _0708_ = state_in[111:104] == 7'b1000000;
  assign _0709_ = state_in[111:104] == 6'b111111;
  assign _0710_ = state_in[111:104] == 6'b111110;
  assign _0711_ = state_in[111:104] == 6'b111101;
  assign _0712_ = state_in[111:104] == 6'b111100;
  assign _0713_ = state_in[111:104] == 6'b111011;
  assign _0714_ = state_in[111:104] == 6'b111010;
  assign _0715_ = state_in[111:104] == 6'b111001;
  assign _0716_ = state_in[111:104] == 6'b111000;
  assign _0717_ = state_in[111:104] == 6'b110111;
  assign _0718_ = state_in[111:104] == 6'b110110;
  assign _0719_ = state_in[111:104] == 6'b110101;
  assign _0720_ = state_in[111:104] == 6'b110100;
  assign _0721_ = state_in[111:104] == 6'b110011;
  assign _0722_ = state_in[111:104] == 6'b110010;
  assign _0723_ = state_in[111:104] == 6'b110001;
  assign _0724_ = state_in[111:104] == 6'b110000;
  assign _0725_ = state_in[111:104] == 6'b101111;
  assign _0726_ = state_in[111:104] == 6'b101110;
  assign _0727_ = state_in[111:104] == 6'b101101;
  assign _0728_ = state_in[111:104] == 6'b101100;
  assign _0729_ = state_in[111:104] == 6'b101011;
  assign _0730_ = state_in[111:104] == 6'b101010;
  assign _0731_ = state_in[111:104] == 6'b101001;
  assign _0732_ = state_in[111:104] == 6'b101000;
  assign _0733_ = state_in[111:104] == 6'b100111;
  assign _0734_ = state_in[111:104] == 6'b100110;
  assign _0735_ = state_in[111:104] == 6'b100101;
  assign _0736_ = state_in[111:104] == 6'b100100;
  assign _0737_ = state_in[111:104] == 6'b100011;
  assign _0738_ = state_in[111:104] == 6'b100010;
  assign _0739_ = state_in[111:104] == 6'b100001;
  assign _0740_ = state_in[111:104] == 6'b100000;
  assign _0741_ = state_in[111:104] == 5'b11111;
  assign _0742_ = state_in[111:104] == 5'b11110;
  assign _0743_ = state_in[111:104] == 5'b11101;
  assign _0744_ = state_in[111:104] == 5'b11100;
  assign _0745_ = state_in[111:104] == 5'b11011;
  assign _0746_ = state_in[111:104] == 5'b11010;
  assign _0747_ = state_in[111:104] == 5'b11001;
  assign _0748_ = state_in[111:104] == 5'b11000;
  assign _0749_ = state_in[111:104] == 5'b10111;
  assign _0750_ = state_in[111:104] == 5'b10110;
  assign _0751_ = state_in[111:104] == 5'b10101;
  assign _0752_ = state_in[111:104] == 5'b10100;
  assign _0753_ = state_in[111:104] == 5'b10011;
  assign _0754_ = state_in[111:104] == 5'b10010;
  assign _0755_ = state_in[111:104] == 5'b10001;
  assign _0756_ = state_in[111:104] == 5'b10000;
  assign _0757_ = state_in[111:104] == 4'b1111;
  assign _0758_ = state_in[111:104] == 4'b1110;
  assign _0759_ = state_in[111:104] == 4'b1101;
  assign _0760_ = state_in[111:104] == 4'b1100;
  assign _0761_ = state_in[111:104] == 4'b1011;
  assign _0762_ = state_in[111:104] == 4'b1010;
  assign _0763_ = state_in[111:104] == 4'b1001;
  assign _0764_ = state_in[111:104] == 4'b1000;
  assign _0765_ = state_in[111:104] == 3'b111;
  assign _0766_ = state_in[111:104] == 3'b110;
  assign _0767_ = state_in[111:104] == 3'b101;
  assign _0768_ = state_in[111:104] == 3'b100;
  assign _0769_ = state_in[111:104] == 2'b11;
  assign _0770_ = state_in[111:104] == 2'b10;
  assign _0771_ = state_in[111:104] == 1'b1;
  assign _0772_ = ! state_in[111:104];
  always @(posedge clk)
      \t0.t2.s4.out <= _0773_;
  logic [255:0] fangyuan6;
  assign fangyuan6 = { _0772_, _0771_, _0770_, _0769_, _0768_, _0767_, _0766_, _0765_, _0764_, _0763_, _0762_, _0761_, _0760_, _0759_, _0758_, _0757_, _0756_, _0755_, _0754_, _0753_, _0752_, _0751_, _0750_, _0749_, _0748_, _0747_, _0746_, _0745_, _0744_, _0743_, _0742_, _0741_, _0740_, _0739_, _0738_, _0737_, _0736_, _0735_, _0734_, _0733_, _0732_, _0731_, _0730_, _0729_, _0728_, _0727_, _0726_, _0725_, _0724_, _0723_, _0722_, _0721_, _0720_, _0719_, _0718_, _0717_, _0716_, _0715_, _0714_, _0713_, _0712_, _0711_, _0710_, _0709_, _0708_, _0707_, _0706_, _0705_, _0704_, _0703_, _0702_, _0701_, _0700_, _0699_, _0698_, _0697_, _0696_, _0695_, _0694_, _0693_, _0692_, _0691_, _0690_, _0689_, _0688_, _0687_, _0686_, _0685_, _0684_, _0683_, _0682_, _0681_, _0680_, _0679_, _0678_, _0677_, _0676_, _0675_, _0674_, _0673_, _0672_, _0671_, _0670_, _0669_, _0668_, _0667_, _0666_, _0665_, _0664_, _0663_, _0662_, _0661_, _0660_, _0659_, _0658_, _0657_, _0656_, _0655_, _0654_, _0653_, _0652_, _0651_, _0650_, _0649_, _0648_, _0647_, _0646_, _0645_, _0644_, _0643_, _0642_, _0641_, _0640_, _0639_, _0638_, _0637_, _0636_, _0635_, _0634_, _0633_, _0632_, _0631_, _0630_, _0629_, _0628_, _0627_, _0626_, _0625_, _0624_, _0623_, _0622_, _0621_, _0620_, _0619_, _0618_, _0617_, _0616_, _0615_, _0614_, _0613_, _0612_, _0611_, _0610_, _0609_, _0608_, _0607_, _0606_, _0605_, _0604_, _0603_, _0602_, _0601_, _0600_, _0599_, _0598_, _0597_, _0596_, _0595_, _0594_, _0593_, _0592_, _0591_, _0590_, _0589_, _0588_, _0587_, _0586_, _0585_, _0584_, _0583_, _0582_, _0581_, _0580_, _0579_, _0578_, _0577_, _0576_, _0575_, _0574_, _0573_, _0572_, _0571_, _0570_, _0569_, _0568_, _0567_, _0566_, _0565_, _0564_, _0563_, _0562_, _0561_, _0560_, _0559_, _0558_, _0557_, _0556_, _0555_, _0554_, _0553_, _0552_, _0551_, _0550_, _0549_, _0548_, _0547_, _0546_, _0545_, _0544_, _0543_, _0542_, _0541_, _0540_, _0539_, _0538_, _0537_, _0536_, _0535_, _0534_, _0533_, _0532_, _0531_, _0530_, _0529_, _0528_, _0527_, _0526_, _0525_, _0524_, _0523_, _0522_, _0521_, _0520_, _0519_, _0518_, _0517_ };

  always @(\t0.t2.s4.out or fangyuan6) begin
    casez (fangyuan6)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0773_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0773_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0773_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0773_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0773_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0773_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0773_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0773_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0773_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0773_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0773_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0773_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0773_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0773_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0773_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0773_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0773_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0773_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0773_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0773_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0773_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0773_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0773_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0773_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0773_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0773_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0773_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0773_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0773_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0773_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0773_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0773_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0773_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0773_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0773_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0773_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0773_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0773_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0773_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0773_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0773_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0773_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0773_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0773_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0773_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0773_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0773_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0773_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0773_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0773_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0773_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0773_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0773_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0773_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0773_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0773_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0773_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0773_ = 8'b11000110 ;
      default:
        _0773_ = \t0.t2.s4.out ;
    endcase
  end
  assign p03[15:8] = \t0.t3.s0.out ^ \t0.t3.s4.out ;
  always @(posedge clk)
      \t0.t3.s0.out <= _0774_;
  logic [255:0] fangyuan7;
  assign fangyuan7 = { _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0944_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_ };

  always @(\t0.t3.s0.out or fangyuan7) begin
    casez (fangyuan7)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _0774_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _0774_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _0774_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _0774_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _0774_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _0774_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _0774_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _0774_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _0774_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _0774_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _0774_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _0774_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _0774_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _0774_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _0774_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _0774_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _0774_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _0774_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _0774_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _0774_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _0774_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _0774_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _0774_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _0774_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _0774_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _0774_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _0774_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _0774_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _0774_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _0774_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _0774_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _0774_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _0774_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _0774_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _0774_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _0774_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _0774_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _0774_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _0774_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _0774_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _0774_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _0774_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _0774_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _0774_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _0774_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _0774_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _0774_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _0774_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _0774_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _0774_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _0774_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _0774_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _0774_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _0774_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _0774_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _0774_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _0774_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _0774_ = 8'b01100011 ;
      default:
        _0774_ = \t0.t3.s0.out ;
    endcase
  end
  assign _0775_ = state_in[103:96] == 8'b11111111;
  assign _0776_ = state_in[103:96] == 8'b11111110;
  assign _0777_ = state_in[103:96] == 8'b11111101;
  assign _0778_ = state_in[103:96] == 8'b11111100;
  assign _0779_ = state_in[103:96] == 8'b11111011;
  assign _0780_ = state_in[103:96] == 8'b11111010;
  assign _0781_ = state_in[103:96] == 8'b11111001;
  assign _0782_ = state_in[103:96] == 8'b11111000;
  assign _0783_ = state_in[103:96] == 8'b11110111;
  assign _0784_ = state_in[103:96] == 8'b11110110;
  assign _0785_ = state_in[103:96] == 8'b11110101;
  assign _0786_ = state_in[103:96] == 8'b11110100;
  assign _0787_ = state_in[103:96] == 8'b11110011;
  assign _0788_ = state_in[103:96] == 8'b11110010;
  assign _0789_ = state_in[103:96] == 8'b11110001;
  assign _0790_ = state_in[103:96] == 8'b11110000;
  assign _0791_ = state_in[103:96] == 8'b11101111;
  assign _0792_ = state_in[103:96] == 8'b11101110;
  assign _0793_ = state_in[103:96] == 8'b11101101;
  assign _0794_ = state_in[103:96] == 8'b11101100;
  assign _0795_ = state_in[103:96] == 8'b11101011;
  assign _0796_ = state_in[103:96] == 8'b11101010;
  assign _0797_ = state_in[103:96] == 8'b11101001;
  assign _0798_ = state_in[103:96] == 8'b11101000;
  assign _0799_ = state_in[103:96] == 8'b11100111;
  assign _0800_ = state_in[103:96] == 8'b11100110;
  assign _0801_ = state_in[103:96] == 8'b11100101;
  assign _0802_ = state_in[103:96] == 8'b11100100;
  assign _0803_ = state_in[103:96] == 8'b11100011;
  assign _0804_ = state_in[103:96] == 8'b11100010;
  assign _0805_ = state_in[103:96] == 8'b11100001;
  assign _0806_ = state_in[103:96] == 8'b11100000;
  assign _0807_ = state_in[103:96] == 8'b11011111;
  assign _0808_ = state_in[103:96] == 8'b11011110;
  assign _0809_ = state_in[103:96] == 8'b11011101;
  assign _0810_ = state_in[103:96] == 8'b11011100;
  assign _0811_ = state_in[103:96] == 8'b11011011;
  assign _0812_ = state_in[103:96] == 8'b11011010;
  assign _0813_ = state_in[103:96] == 8'b11011001;
  assign _0814_ = state_in[103:96] == 8'b11011000;
  assign _0815_ = state_in[103:96] == 8'b11010111;
  assign _0816_ = state_in[103:96] == 8'b11010110;
  assign _0817_ = state_in[103:96] == 8'b11010101;
  assign _0818_ = state_in[103:96] == 8'b11010100;
  assign _0819_ = state_in[103:96] == 8'b11010011;
  assign _0820_ = state_in[103:96] == 8'b11010010;
  assign _0821_ = state_in[103:96] == 8'b11010001;
  assign _0822_ = state_in[103:96] == 8'b11010000;
  assign _0823_ = state_in[103:96] == 8'b11001111;
  assign _0824_ = state_in[103:96] == 8'b11001110;
  assign _0825_ = state_in[103:96] == 8'b11001101;
  assign _0826_ = state_in[103:96] == 8'b11001100;
  assign _0827_ = state_in[103:96] == 8'b11001011;
  assign _0828_ = state_in[103:96] == 8'b11001010;
  assign _0829_ = state_in[103:96] == 8'b11001001;
  assign _0830_ = state_in[103:96] == 8'b11001000;
  assign _0831_ = state_in[103:96] == 8'b11000111;
  assign _0832_ = state_in[103:96] == 8'b11000110;
  assign _0833_ = state_in[103:96] == 8'b11000101;
  assign _0834_ = state_in[103:96] == 8'b11000100;
  assign _0835_ = state_in[103:96] == 8'b11000011;
  assign _0836_ = state_in[103:96] == 8'b11000010;
  assign _0837_ = state_in[103:96] == 8'b11000001;
  assign _0838_ = state_in[103:96] == 8'b11000000;
  assign _0839_ = state_in[103:96] == 8'b10111111;
  assign _0840_ = state_in[103:96] == 8'b10111110;
  assign _0841_ = state_in[103:96] == 8'b10111101;
  assign _0842_ = state_in[103:96] == 8'b10111100;
  assign _0843_ = state_in[103:96] == 8'b10111011;
  assign _0844_ = state_in[103:96] == 8'b10111010;
  assign _0845_ = state_in[103:96] == 8'b10111001;
  assign _0846_ = state_in[103:96] == 8'b10111000;
  assign _0847_ = state_in[103:96] == 8'b10110111;
  assign _0848_ = state_in[103:96] == 8'b10110110;
  assign _0849_ = state_in[103:96] == 8'b10110101;
  assign _0850_ = state_in[103:96] == 8'b10110100;
  assign _0851_ = state_in[103:96] == 8'b10110011;
  assign _0852_ = state_in[103:96] == 8'b10110010;
  assign _0853_ = state_in[103:96] == 8'b10110001;
  assign _0854_ = state_in[103:96] == 8'b10110000;
  assign _0855_ = state_in[103:96] == 8'b10101111;
  assign _0856_ = state_in[103:96] == 8'b10101110;
  assign _0857_ = state_in[103:96] == 8'b10101101;
  assign _0858_ = state_in[103:96] == 8'b10101100;
  assign _0859_ = state_in[103:96] == 8'b10101011;
  assign _0860_ = state_in[103:96] == 8'b10101010;
  assign _0861_ = state_in[103:96] == 8'b10101001;
  assign _0862_ = state_in[103:96] == 8'b10101000;
  assign _0863_ = state_in[103:96] == 8'b10100111;
  assign _0864_ = state_in[103:96] == 8'b10100110;
  assign _0865_ = state_in[103:96] == 8'b10100101;
  assign _0866_ = state_in[103:96] == 8'b10100100;
  assign _0867_ = state_in[103:96] == 8'b10100011;
  assign _0868_ = state_in[103:96] == 8'b10100010;
  assign _0869_ = state_in[103:96] == 8'b10100001;
  assign _0870_ = state_in[103:96] == 8'b10100000;
  assign _0871_ = state_in[103:96] == 8'b10011111;
  assign _0872_ = state_in[103:96] == 8'b10011110;
  assign _0873_ = state_in[103:96] == 8'b10011101;
  assign _0874_ = state_in[103:96] == 8'b10011100;
  assign _0875_ = state_in[103:96] == 8'b10011011;
  assign _0876_ = state_in[103:96] == 8'b10011010;
  assign _0877_ = state_in[103:96] == 8'b10011001;
  assign _0878_ = state_in[103:96] == 8'b10011000;
  assign _0879_ = state_in[103:96] == 8'b10010111;
  assign _0880_ = state_in[103:96] == 8'b10010110;
  assign _0881_ = state_in[103:96] == 8'b10010101;
  assign _0882_ = state_in[103:96] == 8'b10010100;
  assign _0883_ = state_in[103:96] == 8'b10010011;
  assign _0884_ = state_in[103:96] == 8'b10010010;
  assign _0885_ = state_in[103:96] == 8'b10010001;
  assign _0886_ = state_in[103:96] == 8'b10010000;
  assign _0887_ = state_in[103:96] == 8'b10001111;
  assign _0888_ = state_in[103:96] == 8'b10001110;
  assign _0889_ = state_in[103:96] == 8'b10001101;
  assign _0890_ = state_in[103:96] == 8'b10001100;
  assign _0891_ = state_in[103:96] == 8'b10001011;
  assign _0892_ = state_in[103:96] == 8'b10001010;
  assign _0893_ = state_in[103:96] == 8'b10001001;
  assign _0894_ = state_in[103:96] == 8'b10001000;
  assign _0895_ = state_in[103:96] == 8'b10000111;
  assign _0896_ = state_in[103:96] == 8'b10000110;
  assign _0897_ = state_in[103:96] == 8'b10000101;
  assign _0898_ = state_in[103:96] == 8'b10000100;
  assign _0899_ = state_in[103:96] == 8'b10000011;
  assign _0900_ = state_in[103:96] == 8'b10000010;
  assign _0901_ = state_in[103:96] == 8'b10000001;
  assign _0902_ = state_in[103:96] == 8'b10000000;
  assign _0903_ = state_in[103:96] == 7'b1111111;
  assign _0904_ = state_in[103:96] == 7'b1111110;
  assign _0905_ = state_in[103:96] == 7'b1111101;
  assign _0906_ = state_in[103:96] == 7'b1111100;
  assign _0907_ = state_in[103:96] == 7'b1111011;
  assign _0908_ = state_in[103:96] == 7'b1111010;
  assign _0909_ = state_in[103:96] == 7'b1111001;
  assign _0910_ = state_in[103:96] == 7'b1111000;
  assign _0911_ = state_in[103:96] == 7'b1110111;
  assign _0912_ = state_in[103:96] == 7'b1110110;
  assign _0913_ = state_in[103:96] == 7'b1110101;
  assign _0914_ = state_in[103:96] == 7'b1110100;
  assign _0915_ = state_in[103:96] == 7'b1110011;
  assign _0916_ = state_in[103:96] == 7'b1110010;
  assign _0917_ = state_in[103:96] == 7'b1110001;
  assign _0918_ = state_in[103:96] == 7'b1110000;
  assign _0919_ = state_in[103:96] == 7'b1101111;
  assign _0920_ = state_in[103:96] == 7'b1101110;
  assign _0921_ = state_in[103:96] == 7'b1101101;
  assign _0922_ = state_in[103:96] == 7'b1101100;
  assign _0923_ = state_in[103:96] == 7'b1101011;
  assign _0924_ = state_in[103:96] == 7'b1101010;
  assign _0925_ = state_in[103:96] == 7'b1101001;
  assign _0926_ = state_in[103:96] == 7'b1101000;
  assign _0927_ = state_in[103:96] == 7'b1100111;
  assign _0928_ = state_in[103:96] == 7'b1100110;
  assign _0929_ = state_in[103:96] == 7'b1100101;
  assign _0930_ = state_in[103:96] == 7'b1100100;
  assign _0931_ = state_in[103:96] == 7'b1100011;
  assign _0932_ = state_in[103:96] == 7'b1100010;
  assign _0933_ = state_in[103:96] == 7'b1100001;
  assign _0934_ = state_in[103:96] == 7'b1100000;
  assign _0935_ = state_in[103:96] == 7'b1011111;
  assign _0936_ = state_in[103:96] == 7'b1011110;
  assign _0937_ = state_in[103:96] == 7'b1011101;
  assign _0938_ = state_in[103:96] == 7'b1011100;
  assign _0939_ = state_in[103:96] == 7'b1011011;
  assign _0940_ = state_in[103:96] == 7'b1011010;
  assign _0941_ = state_in[103:96] == 7'b1011001;
  assign _0942_ = state_in[103:96] == 7'b1011000;
  assign _0943_ = state_in[103:96] == 7'b1010111;
  assign _0944_ = state_in[103:96] == 7'b1010110;
  assign _0945_ = state_in[103:96] == 7'b1010101;
  assign _0946_ = state_in[103:96] == 7'b1010100;
  assign _0947_ = state_in[103:96] == 7'b1010011;
  assign _0948_ = state_in[103:96] == 7'b1010010;
  assign _0949_ = state_in[103:96] == 7'b1010001;
  assign _0950_ = state_in[103:96] == 7'b1010000;
  assign _0951_ = state_in[103:96] == 7'b1001111;
  assign _0952_ = state_in[103:96] == 7'b1001110;
  assign _0953_ = state_in[103:96] == 7'b1001101;
  assign _0954_ = state_in[103:96] == 7'b1001100;
  assign _0955_ = state_in[103:96] == 7'b1001011;
  assign _0956_ = state_in[103:96] == 7'b1001010;
  assign _0957_ = state_in[103:96] == 7'b1001001;
  assign _0958_ = state_in[103:96] == 7'b1001000;
  assign _0959_ = state_in[103:96] == 7'b1000111;
  assign _0960_ = state_in[103:96] == 7'b1000110;
  assign _0961_ = state_in[103:96] == 7'b1000101;
  assign _0962_ = state_in[103:96] == 7'b1000100;
  assign _0963_ = state_in[103:96] == 7'b1000011;
  assign _0964_ = state_in[103:96] == 7'b1000010;
  assign _0965_ = state_in[103:96] == 7'b1000001;
  assign _0966_ = state_in[103:96] == 7'b1000000;
  assign _0967_ = state_in[103:96] == 6'b111111;
  assign _0968_ = state_in[103:96] == 6'b111110;
  assign _0969_ = state_in[103:96] == 6'b111101;
  assign _0970_ = state_in[103:96] == 6'b111100;
  assign _0971_ = state_in[103:96] == 6'b111011;
  assign _0972_ = state_in[103:96] == 6'b111010;
  assign _0973_ = state_in[103:96] == 6'b111001;
  assign _0974_ = state_in[103:96] == 6'b111000;
  assign _0975_ = state_in[103:96] == 6'b110111;
  assign _0976_ = state_in[103:96] == 6'b110110;
  assign _0977_ = state_in[103:96] == 6'b110101;
  assign _0978_ = state_in[103:96] == 6'b110100;
  assign _0979_ = state_in[103:96] == 6'b110011;
  assign _0980_ = state_in[103:96] == 6'b110010;
  assign _0981_ = state_in[103:96] == 6'b110001;
  assign _0982_ = state_in[103:96] == 6'b110000;
  assign _0983_ = state_in[103:96] == 6'b101111;
  assign _0984_ = state_in[103:96] == 6'b101110;
  assign _0985_ = state_in[103:96] == 6'b101101;
  assign _0986_ = state_in[103:96] == 6'b101100;
  assign _0987_ = state_in[103:96] == 6'b101011;
  assign _0988_ = state_in[103:96] == 6'b101010;
  assign _0989_ = state_in[103:96] == 6'b101001;
  assign _0990_ = state_in[103:96] == 6'b101000;
  assign _0991_ = state_in[103:96] == 6'b100111;
  assign _0992_ = state_in[103:96] == 6'b100110;
  assign _0993_ = state_in[103:96] == 6'b100101;
  assign _0994_ = state_in[103:96] == 6'b100100;
  assign _0995_ = state_in[103:96] == 6'b100011;
  assign _0996_ = state_in[103:96] == 6'b100010;
  assign _0997_ = state_in[103:96] == 6'b100001;
  assign _0998_ = state_in[103:96] == 6'b100000;
  assign _0999_ = state_in[103:96] == 5'b11111;
  assign _1000_ = state_in[103:96] == 5'b11110;
  assign _1001_ = state_in[103:96] == 5'b11101;
  assign _1002_ = state_in[103:96] == 5'b11100;
  assign _1003_ = state_in[103:96] == 5'b11011;
  assign _1004_ = state_in[103:96] == 5'b11010;
  assign _1005_ = state_in[103:96] == 5'b11001;
  assign _1006_ = state_in[103:96] == 5'b11000;
  assign _1007_ = state_in[103:96] == 5'b10111;
  assign _1008_ = state_in[103:96] == 5'b10110;
  assign _1009_ = state_in[103:96] == 5'b10101;
  assign _1010_ = state_in[103:96] == 5'b10100;
  assign _1011_ = state_in[103:96] == 5'b10011;
  assign _1012_ = state_in[103:96] == 5'b10010;
  assign _1013_ = state_in[103:96] == 5'b10001;
  assign _1014_ = state_in[103:96] == 5'b10000;
  assign _1015_ = state_in[103:96] == 4'b1111;
  assign _1016_ = state_in[103:96] == 4'b1110;
  assign _1017_ = state_in[103:96] == 4'b1101;
  assign _1018_ = state_in[103:96] == 4'b1100;
  assign _1019_ = state_in[103:96] == 4'b1011;
  assign _1020_ = state_in[103:96] == 4'b1010;
  assign _1021_ = state_in[103:96] == 4'b1001;
  assign _1022_ = state_in[103:96] == 4'b1000;
  assign _1023_ = state_in[103:96] == 3'b111;
  assign _1024_ = state_in[103:96] == 3'b110;
  assign _1025_ = state_in[103:96] == 3'b101;
  assign _1026_ = state_in[103:96] == 3'b100;
  assign _1027_ = state_in[103:96] == 2'b11;
  assign _1028_ = state_in[103:96] == 2'b10;
  assign _1029_ = state_in[103:96] == 1'b1;
  assign _1030_ = ! state_in[103:96];
  always @(posedge clk)
      \t0.t3.s4.out <= _1031_;
  logic [255:0] fangyuan8;
  assign fangyuan8 = { _1030_, _1029_, _1028_, _1027_, _1026_, _1025_, _1024_, _1023_, _1022_, _1021_, _1020_, _1019_, _1018_, _1017_, _1016_, _1015_, _1014_, _1013_, _1012_, _1011_, _1010_, _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_, _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_, _0947_, _0946_, _0945_, _0944_, _0943_, _0942_, _0941_, _0940_, _0939_, _0938_, _0937_, _0936_, _0935_, _0934_, _0933_, _0932_, _0931_, _0930_, _0929_, _0928_, _0927_, _0926_, _0925_, _0924_, _0923_, _0922_, _0921_, _0920_, _0919_, _0918_, _0917_, _0916_, _0915_, _0914_, _0913_, _0912_, _0911_, _0910_, _0909_, _0908_, _0907_, _0906_, _0905_, _0904_, _0903_, _0902_, _0901_, _0900_, _0899_, _0898_, _0897_, _0896_, _0895_, _0894_, _0893_, _0892_, _0891_, _0890_, _0889_, _0888_, _0887_, _0886_, _0885_, _0884_, _0883_, _0882_, _0881_, _0880_, _0879_, _0878_, _0877_, _0876_, _0875_, _0874_, _0873_, _0872_, _0871_, _0870_, _0869_, _0868_, _0867_, _0866_, _0865_, _0864_, _0863_, _0862_, _0861_, _0860_, _0859_, _0858_, _0857_, _0856_, _0855_, _0854_, _0853_, _0852_, _0851_, _0850_, _0849_, _0848_, _0847_, _0846_, _0845_, _0844_, _0843_, _0842_, _0841_, _0840_, _0839_, _0838_, _0837_, _0836_, _0835_, _0834_, _0833_, _0832_, _0831_, _0830_, _0829_, _0828_, _0827_, _0826_, _0825_, _0824_, _0823_, _0822_, _0821_, _0820_, _0819_, _0818_, _0817_, _0816_, _0815_, _0814_, _0813_, _0812_, _0811_, _0810_, _0809_, _0808_, _0807_, _0806_, _0805_, _0804_, _0803_, _0802_, _0801_, _0800_, _0799_, _0798_, _0797_, _0796_, _0795_, _0794_, _0793_, _0792_, _0791_, _0790_, _0789_, _0788_, _0787_, _0786_, _0785_, _0784_, _0783_, _0782_, _0781_, _0780_, _0779_, _0778_, _0777_, _0776_, _0775_ };

  always @(\t0.t3.s4.out or fangyuan8) begin
    casez (fangyuan8)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1031_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1031_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1031_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1031_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1031_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1031_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1031_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1031_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1031_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1031_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1031_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1031_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1031_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1031_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1031_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1031_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1031_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1031_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1031_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1031_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1031_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1031_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1031_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1031_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1031_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1031_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1031_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1031_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1031_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1031_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1031_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1031_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1031_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1031_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1031_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1031_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1031_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1031_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1031_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1031_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1031_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1031_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1031_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1031_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1031_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1031_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1031_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1031_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1031_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1031_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1031_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1031_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1031_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1031_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1031_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1031_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1031_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1031_ = 8'b11000110 ;
      default:
        _1031_ = \t0.t3.s4.out ;
    endcase
  end
  assign p10[7:0] = \t1.t0.s0.out ^ \t1.t0.s4.out ;
  always @(posedge clk)
      \t1.t0.s0.out <= _1032_;
  logic [255:0] fangyuan9;
  assign fangyuan9 = { _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_, _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_ };

  always @(\t1.t0.s0.out or fangyuan9) begin
    casez (fangyuan9)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1032_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1032_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1032_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1032_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1032_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1032_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1032_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1032_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1032_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1032_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1032_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1032_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1032_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1032_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1032_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1032_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1032_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1032_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1032_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1032_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1032_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1032_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1032_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1032_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1032_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1032_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1032_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1032_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1032_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1032_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1032_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1032_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1032_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1032_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1032_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1032_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1032_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1032_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1032_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1032_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1032_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1032_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1032_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1032_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1032_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1032_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1032_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1032_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1032_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1032_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1032_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1032_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1032_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1032_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1032_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1032_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1032_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1032_ = 8'b01100011 ;
      default:
        _1032_ = \t1.t0.s0.out ;
    endcase
  end
  assign _1033_ = state_in[95:88] == 8'b11111111;
  assign _1034_ = state_in[95:88] == 8'b11111110;
  assign _1035_ = state_in[95:88] == 8'b11111101;
  assign _1036_ = state_in[95:88] == 8'b11111100;
  assign _1037_ = state_in[95:88] == 8'b11111011;
  assign _1038_ = state_in[95:88] == 8'b11111010;
  assign _1039_ = state_in[95:88] == 8'b11111001;
  assign _1040_ = state_in[95:88] == 8'b11111000;
  assign _1041_ = state_in[95:88] == 8'b11110111;
  assign _1042_ = state_in[95:88] == 8'b11110110;
  assign _1043_ = state_in[95:88] == 8'b11110101;
  assign _1044_ = state_in[95:88] == 8'b11110100;
  assign _1045_ = state_in[95:88] == 8'b11110011;
  assign _1046_ = state_in[95:88] == 8'b11110010;
  assign _1047_ = state_in[95:88] == 8'b11110001;
  assign _1048_ = state_in[95:88] == 8'b11110000;
  assign _1049_ = state_in[95:88] == 8'b11101111;
  assign _1050_ = state_in[95:88] == 8'b11101110;
  assign _1051_ = state_in[95:88] == 8'b11101101;
  assign _1052_ = state_in[95:88] == 8'b11101100;
  assign _1053_ = state_in[95:88] == 8'b11101011;
  assign _1054_ = state_in[95:88] == 8'b11101010;
  assign _1055_ = state_in[95:88] == 8'b11101001;
  assign _1056_ = state_in[95:88] == 8'b11101000;
  assign _1057_ = state_in[95:88] == 8'b11100111;
  assign _1058_ = state_in[95:88] == 8'b11100110;
  assign _1059_ = state_in[95:88] == 8'b11100101;
  assign _1060_ = state_in[95:88] == 8'b11100100;
  assign _1061_ = state_in[95:88] == 8'b11100011;
  assign _1062_ = state_in[95:88] == 8'b11100010;
  assign _1063_ = state_in[95:88] == 8'b11100001;
  assign _1064_ = state_in[95:88] == 8'b11100000;
  assign _1065_ = state_in[95:88] == 8'b11011111;
  assign _1066_ = state_in[95:88] == 8'b11011110;
  assign _1067_ = state_in[95:88] == 8'b11011101;
  assign _1068_ = state_in[95:88] == 8'b11011100;
  assign _1069_ = state_in[95:88] == 8'b11011011;
  assign _1070_ = state_in[95:88] == 8'b11011010;
  assign _1071_ = state_in[95:88] == 8'b11011001;
  assign _1072_ = state_in[95:88] == 8'b11011000;
  assign _1073_ = state_in[95:88] == 8'b11010111;
  assign _1074_ = state_in[95:88] == 8'b11010110;
  assign _1075_ = state_in[95:88] == 8'b11010101;
  assign _1076_ = state_in[95:88] == 8'b11010100;
  assign _1077_ = state_in[95:88] == 8'b11010011;
  assign _1078_ = state_in[95:88] == 8'b11010010;
  assign _1079_ = state_in[95:88] == 8'b11010001;
  assign _1080_ = state_in[95:88] == 8'b11010000;
  assign _1081_ = state_in[95:88] == 8'b11001111;
  assign _1082_ = state_in[95:88] == 8'b11001110;
  assign _1083_ = state_in[95:88] == 8'b11001101;
  assign _1084_ = state_in[95:88] == 8'b11001100;
  assign _1085_ = state_in[95:88] == 8'b11001011;
  assign _1086_ = state_in[95:88] == 8'b11001010;
  assign _1087_ = state_in[95:88] == 8'b11001001;
  assign _1088_ = state_in[95:88] == 8'b11001000;
  assign _1089_ = state_in[95:88] == 8'b11000111;
  assign _1090_ = state_in[95:88] == 8'b11000110;
  assign _1091_ = state_in[95:88] == 8'b11000101;
  assign _1092_ = state_in[95:88] == 8'b11000100;
  assign _1093_ = state_in[95:88] == 8'b11000011;
  assign _1094_ = state_in[95:88] == 8'b11000010;
  assign _1095_ = state_in[95:88] == 8'b11000001;
  assign _1096_ = state_in[95:88] == 8'b11000000;
  assign _1097_ = state_in[95:88] == 8'b10111111;
  assign _1098_ = state_in[95:88] == 8'b10111110;
  assign _1099_ = state_in[95:88] == 8'b10111101;
  assign _1100_ = state_in[95:88] == 8'b10111100;
  assign _1101_ = state_in[95:88] == 8'b10111011;
  assign _1102_ = state_in[95:88] == 8'b10111010;
  assign _1103_ = state_in[95:88] == 8'b10111001;
  assign _1104_ = state_in[95:88] == 8'b10111000;
  assign _1105_ = state_in[95:88] == 8'b10110111;
  assign _1106_ = state_in[95:88] == 8'b10110110;
  assign _1107_ = state_in[95:88] == 8'b10110101;
  assign _1108_ = state_in[95:88] == 8'b10110100;
  assign _1109_ = state_in[95:88] == 8'b10110011;
  assign _1110_ = state_in[95:88] == 8'b10110010;
  assign _1111_ = state_in[95:88] == 8'b10110001;
  assign _1112_ = state_in[95:88] == 8'b10110000;
  assign _1113_ = state_in[95:88] == 8'b10101111;
  assign _1114_ = state_in[95:88] == 8'b10101110;
  assign _1115_ = state_in[95:88] == 8'b10101101;
  assign _1116_ = state_in[95:88] == 8'b10101100;
  assign _1117_ = state_in[95:88] == 8'b10101011;
  assign _1118_ = state_in[95:88] == 8'b10101010;
  assign _1119_ = state_in[95:88] == 8'b10101001;
  assign _1120_ = state_in[95:88] == 8'b10101000;
  assign _1121_ = state_in[95:88] == 8'b10100111;
  assign _1122_ = state_in[95:88] == 8'b10100110;
  assign _1123_ = state_in[95:88] == 8'b10100101;
  assign _1124_ = state_in[95:88] == 8'b10100100;
  assign _1125_ = state_in[95:88] == 8'b10100011;
  assign _1126_ = state_in[95:88] == 8'b10100010;
  assign _1127_ = state_in[95:88] == 8'b10100001;
  assign _1128_ = state_in[95:88] == 8'b10100000;
  assign _1129_ = state_in[95:88] == 8'b10011111;
  assign _1130_ = state_in[95:88] == 8'b10011110;
  assign _1131_ = state_in[95:88] == 8'b10011101;
  assign _1132_ = state_in[95:88] == 8'b10011100;
  assign _1133_ = state_in[95:88] == 8'b10011011;
  assign _1134_ = state_in[95:88] == 8'b10011010;
  assign _1135_ = state_in[95:88] == 8'b10011001;
  assign _1136_ = state_in[95:88] == 8'b10011000;
  assign _1137_ = state_in[95:88] == 8'b10010111;
  assign _1138_ = state_in[95:88] == 8'b10010110;
  assign _1139_ = state_in[95:88] == 8'b10010101;
  assign _1140_ = state_in[95:88] == 8'b10010100;
  assign _1141_ = state_in[95:88] == 8'b10010011;
  assign _1142_ = state_in[95:88] == 8'b10010010;
  assign _1143_ = state_in[95:88] == 8'b10010001;
  assign _1144_ = state_in[95:88] == 8'b10010000;
  assign _1145_ = state_in[95:88] == 8'b10001111;
  assign _1146_ = state_in[95:88] == 8'b10001110;
  assign _1147_ = state_in[95:88] == 8'b10001101;
  assign _1148_ = state_in[95:88] == 8'b10001100;
  assign _1149_ = state_in[95:88] == 8'b10001011;
  assign _1150_ = state_in[95:88] == 8'b10001010;
  assign _1151_ = state_in[95:88] == 8'b10001001;
  assign _1152_ = state_in[95:88] == 8'b10001000;
  assign _1153_ = state_in[95:88] == 8'b10000111;
  assign _1154_ = state_in[95:88] == 8'b10000110;
  assign _1155_ = state_in[95:88] == 8'b10000101;
  assign _1156_ = state_in[95:88] == 8'b10000100;
  assign _1157_ = state_in[95:88] == 8'b10000011;
  assign _1158_ = state_in[95:88] == 8'b10000010;
  assign _1159_ = state_in[95:88] == 8'b10000001;
  assign _1160_ = state_in[95:88] == 8'b10000000;
  assign _1161_ = state_in[95:88] == 7'b1111111;
  assign _1162_ = state_in[95:88] == 7'b1111110;
  assign _1163_ = state_in[95:88] == 7'b1111101;
  assign _1164_ = state_in[95:88] == 7'b1111100;
  assign _1165_ = state_in[95:88] == 7'b1111011;
  assign _1166_ = state_in[95:88] == 7'b1111010;
  assign _1167_ = state_in[95:88] == 7'b1111001;
  assign _1168_ = state_in[95:88] == 7'b1111000;
  assign _1169_ = state_in[95:88] == 7'b1110111;
  assign _1170_ = state_in[95:88] == 7'b1110110;
  assign _1171_ = state_in[95:88] == 7'b1110101;
  assign _1172_ = state_in[95:88] == 7'b1110100;
  assign _1173_ = state_in[95:88] == 7'b1110011;
  assign _1174_ = state_in[95:88] == 7'b1110010;
  assign _1175_ = state_in[95:88] == 7'b1110001;
  assign _1176_ = state_in[95:88] == 7'b1110000;
  assign _1177_ = state_in[95:88] == 7'b1101111;
  assign _1178_ = state_in[95:88] == 7'b1101110;
  assign _1179_ = state_in[95:88] == 7'b1101101;
  assign _1180_ = state_in[95:88] == 7'b1101100;
  assign _1181_ = state_in[95:88] == 7'b1101011;
  assign _1182_ = state_in[95:88] == 7'b1101010;
  assign _1183_ = state_in[95:88] == 7'b1101001;
  assign _1184_ = state_in[95:88] == 7'b1101000;
  assign _1185_ = state_in[95:88] == 7'b1100111;
  assign _1186_ = state_in[95:88] == 7'b1100110;
  assign _1187_ = state_in[95:88] == 7'b1100101;
  assign _1188_ = state_in[95:88] == 7'b1100100;
  assign _1189_ = state_in[95:88] == 7'b1100011;
  assign _1190_ = state_in[95:88] == 7'b1100010;
  assign _1191_ = state_in[95:88] == 7'b1100001;
  assign _1192_ = state_in[95:88] == 7'b1100000;
  assign _1193_ = state_in[95:88] == 7'b1011111;
  assign _1194_ = state_in[95:88] == 7'b1011110;
  assign _1195_ = state_in[95:88] == 7'b1011101;
  assign _1196_ = state_in[95:88] == 7'b1011100;
  assign _1197_ = state_in[95:88] == 7'b1011011;
  assign _1198_ = state_in[95:88] == 7'b1011010;
  assign _1199_ = state_in[95:88] == 7'b1011001;
  assign _1200_ = state_in[95:88] == 7'b1011000;
  assign _1201_ = state_in[95:88] == 7'b1010111;
  assign _1202_ = state_in[95:88] == 7'b1010110;
  assign _1203_ = state_in[95:88] == 7'b1010101;
  assign _1204_ = state_in[95:88] == 7'b1010100;
  assign _1205_ = state_in[95:88] == 7'b1010011;
  assign _1206_ = state_in[95:88] == 7'b1010010;
  assign _1207_ = state_in[95:88] == 7'b1010001;
  assign _1208_ = state_in[95:88] == 7'b1010000;
  assign _1209_ = state_in[95:88] == 7'b1001111;
  assign _1210_ = state_in[95:88] == 7'b1001110;
  assign _1211_ = state_in[95:88] == 7'b1001101;
  assign _1212_ = state_in[95:88] == 7'b1001100;
  assign _1213_ = state_in[95:88] == 7'b1001011;
  assign _1214_ = state_in[95:88] == 7'b1001010;
  assign _1215_ = state_in[95:88] == 7'b1001001;
  assign _1216_ = state_in[95:88] == 7'b1001000;
  assign _1217_ = state_in[95:88] == 7'b1000111;
  assign _1218_ = state_in[95:88] == 7'b1000110;
  assign _1219_ = state_in[95:88] == 7'b1000101;
  assign _1220_ = state_in[95:88] == 7'b1000100;
  assign _1221_ = state_in[95:88] == 7'b1000011;
  assign _1222_ = state_in[95:88] == 7'b1000010;
  assign _1223_ = state_in[95:88] == 7'b1000001;
  assign _1224_ = state_in[95:88] == 7'b1000000;
  assign _1225_ = state_in[95:88] == 6'b111111;
  assign _1226_ = state_in[95:88] == 6'b111110;
  assign _1227_ = state_in[95:88] == 6'b111101;
  assign _1228_ = state_in[95:88] == 6'b111100;
  assign _1229_ = state_in[95:88] == 6'b111011;
  assign _1230_ = state_in[95:88] == 6'b111010;
  assign _1231_ = state_in[95:88] == 6'b111001;
  assign _1232_ = state_in[95:88] == 6'b111000;
  assign _1233_ = state_in[95:88] == 6'b110111;
  assign _1234_ = state_in[95:88] == 6'b110110;
  assign _1235_ = state_in[95:88] == 6'b110101;
  assign _1236_ = state_in[95:88] == 6'b110100;
  assign _1237_ = state_in[95:88] == 6'b110011;
  assign _1238_ = state_in[95:88] == 6'b110010;
  assign _1239_ = state_in[95:88] == 6'b110001;
  assign _1240_ = state_in[95:88] == 6'b110000;
  assign _1241_ = state_in[95:88] == 6'b101111;
  assign _1242_ = state_in[95:88] == 6'b101110;
  assign _1243_ = state_in[95:88] == 6'b101101;
  assign _1244_ = state_in[95:88] == 6'b101100;
  assign _1245_ = state_in[95:88] == 6'b101011;
  assign _1246_ = state_in[95:88] == 6'b101010;
  assign _1247_ = state_in[95:88] == 6'b101001;
  assign _1248_ = state_in[95:88] == 6'b101000;
  assign _1249_ = state_in[95:88] == 6'b100111;
  assign _1250_ = state_in[95:88] == 6'b100110;
  assign _1251_ = state_in[95:88] == 6'b100101;
  assign _1252_ = state_in[95:88] == 6'b100100;
  assign _1253_ = state_in[95:88] == 6'b100011;
  assign _1254_ = state_in[95:88] == 6'b100010;
  assign _1255_ = state_in[95:88] == 6'b100001;
  assign _1256_ = state_in[95:88] == 6'b100000;
  assign _1257_ = state_in[95:88] == 5'b11111;
  assign _1258_ = state_in[95:88] == 5'b11110;
  assign _1259_ = state_in[95:88] == 5'b11101;
  assign _1260_ = state_in[95:88] == 5'b11100;
  assign _1261_ = state_in[95:88] == 5'b11011;
  assign _1262_ = state_in[95:88] == 5'b11010;
  assign _1263_ = state_in[95:88] == 5'b11001;
  assign _1264_ = state_in[95:88] == 5'b11000;
  assign _1265_ = state_in[95:88] == 5'b10111;
  assign _1266_ = state_in[95:88] == 5'b10110;
  assign _1267_ = state_in[95:88] == 5'b10101;
  assign _1268_ = state_in[95:88] == 5'b10100;
  assign _1269_ = state_in[95:88] == 5'b10011;
  assign _1270_ = state_in[95:88] == 5'b10010;
  assign _1271_ = state_in[95:88] == 5'b10001;
  assign _1272_ = state_in[95:88] == 5'b10000;
  assign _1273_ = state_in[95:88] == 4'b1111;
  assign _1274_ = state_in[95:88] == 4'b1110;
  assign _1275_ = state_in[95:88] == 4'b1101;
  assign _1276_ = state_in[95:88] == 4'b1100;
  assign _1277_ = state_in[95:88] == 4'b1011;
  assign _1278_ = state_in[95:88] == 4'b1010;
  assign _1279_ = state_in[95:88] == 4'b1001;
  assign _1280_ = state_in[95:88] == 4'b1000;
  assign _1281_ = state_in[95:88] == 3'b111;
  assign _1282_ = state_in[95:88] == 3'b110;
  assign _1283_ = state_in[95:88] == 3'b101;
  assign _1284_ = state_in[95:88] == 3'b100;
  assign _1285_ = state_in[95:88] == 2'b11;
  assign _1286_ = state_in[95:88] == 2'b10;
  assign _1287_ = state_in[95:88] == 1'b1;
  assign _1288_ = ! state_in[95:88];
  always @(posedge clk)
      \t1.t0.s4.out <= _1289_;
  logic [255:0] fangyuan10;
  assign fangyuan10 = { _1288_, _1287_, _1286_, _1285_, _1284_, _1283_, _1282_, _1281_, _1280_, _1279_, _1278_, _1277_, _1276_, _1275_, _1274_, _1273_, _1272_, _1271_, _1270_, _1269_, _1268_, _1267_, _1266_, _1265_, _1264_, _1263_, _1262_, _1261_, _1260_, _1259_, _1258_, _1257_, _1256_, _1255_, _1254_, _1253_, _1252_, _1251_, _1250_, _1249_, _1248_, _1247_, _1246_, _1245_, _1244_, _1243_, _1242_, _1241_, _1240_, _1239_, _1238_, _1237_, _1236_, _1235_, _1234_, _1233_, _1232_, _1231_, _1230_, _1229_, _1228_, _1227_, _1226_, _1225_, _1224_, _1223_, _1222_, _1221_, _1220_, _1219_, _1218_, _1217_, _1216_, _1215_, _1214_, _1213_, _1212_, _1211_, _1210_, _1209_, _1208_, _1207_, _1206_, _1205_, _1204_, _1203_, _1202_, _1201_, _1200_, _1199_, _1198_, _1197_, _1196_, _1195_, _1194_, _1193_, _1192_, _1191_, _1190_, _1189_, _1188_, _1187_, _1186_, _1185_, _1184_, _1183_, _1182_, _1181_, _1180_, _1179_, _1178_, _1177_, _1176_, _1175_, _1174_, _1173_, _1172_, _1171_, _1170_, _1169_, _1168_, _1167_, _1166_, _1165_, _1164_, _1163_, _1162_, _1161_, _1160_, _1159_, _1158_, _1157_, _1156_, _1155_, _1154_, _1153_, _1152_, _1151_, _1150_, _1149_, _1148_, _1147_, _1146_, _1145_, _1144_, _1143_, _1142_, _1141_, _1140_, _1139_, _1138_, _1137_, _1136_, _1135_, _1134_, _1133_, _1132_, _1131_, _1130_, _1129_, _1128_, _1127_, _1126_, _1125_, _1124_, _1123_, _1122_, _1121_, _1120_, _1119_, _1118_, _1117_, _1116_, _1115_, _1114_, _1113_, _1112_, _1111_, _1110_, _1109_, _1108_, _1107_, _1106_, _1105_, _1104_, _1103_, _1102_, _1101_, _1100_, _1099_, _1098_, _1097_, _1096_, _1095_, _1094_, _1093_, _1092_, _1091_, _1090_, _1089_, _1088_, _1087_, _1086_, _1085_, _1084_, _1083_, _1082_, _1081_, _1080_, _1079_, _1078_, _1077_, _1076_, _1075_, _1074_, _1073_, _1072_, _1071_, _1070_, _1069_, _1068_, _1067_, _1066_, _1065_, _1064_, _1063_, _1062_, _1061_, _1060_, _1059_, _1058_, _1057_, _1056_, _1055_, _1054_, _1053_, _1052_, _1051_, _1050_, _1049_, _1048_, _1047_, _1046_, _1045_, _1044_, _1043_, _1042_, _1041_, _1040_, _1039_, _1038_, _1037_, _1036_, _1035_, _1034_, _1033_ };

  always @(\t1.t0.s4.out or fangyuan10) begin
    casez (fangyuan10)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1289_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1289_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1289_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1289_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1289_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1289_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1289_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1289_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1289_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1289_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1289_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1289_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1289_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1289_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1289_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1289_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1289_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1289_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1289_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1289_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1289_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1289_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1289_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1289_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1289_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1289_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1289_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1289_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1289_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1289_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1289_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1289_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1289_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1289_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1289_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1289_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1289_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1289_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1289_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1289_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1289_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1289_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1289_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1289_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1289_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1289_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1289_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1289_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1289_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1289_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1289_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1289_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1289_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1289_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1289_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1289_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1289_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1289_ = 8'b11000110 ;
      default:
        _1289_ = \t1.t0.s4.out ;
    endcase
  end
  assign p11[31:24] = \t1.t1.s0.out ^ \t1.t1.s4.out ;
  always @(posedge clk)
      \t1.t1.s0.out <= _1290_;
  logic [255:0] fangyuan11;
  assign fangyuan11 = { _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _1472_, _1471_, _1470_, _1469_, _1468_, _1467_, _1466_, _1465_, _1464_, _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_, _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_ };

  always @(\t1.t1.s0.out or fangyuan11) begin
    casez (fangyuan11)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1290_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1290_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1290_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1290_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1290_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1290_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1290_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1290_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1290_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1290_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1290_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1290_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1290_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1290_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1290_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1290_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1290_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1290_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1290_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1290_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1290_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1290_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1290_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1290_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1290_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1290_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1290_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1290_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1290_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1290_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1290_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1290_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1290_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1290_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1290_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1290_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1290_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1290_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1290_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1290_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1290_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1290_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1290_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1290_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1290_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1290_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1290_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1290_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1290_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1290_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1290_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1290_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1290_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1290_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1290_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1290_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1290_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1290_ = 8'b01100011 ;
      default:
        _1290_ = \t1.t1.s0.out ;
    endcase
  end
  assign _1291_ = state_in[87:80] == 8'b11111111;
  assign _1292_ = state_in[87:80] == 8'b11111110;
  assign _1293_ = state_in[87:80] == 8'b11111101;
  assign _1294_ = state_in[87:80] == 8'b11111100;
  assign _1295_ = state_in[87:80] == 8'b11111011;
  assign _1296_ = state_in[87:80] == 8'b11111010;
  assign _1297_ = state_in[87:80] == 8'b11111001;
  assign _1298_ = state_in[87:80] == 8'b11111000;
  assign _1299_ = state_in[87:80] == 8'b11110111;
  assign _1300_ = state_in[87:80] == 8'b11110110;
  assign _1301_ = state_in[87:80] == 8'b11110101;
  assign _1302_ = state_in[87:80] == 8'b11110100;
  assign _1303_ = state_in[87:80] == 8'b11110011;
  assign _1304_ = state_in[87:80] == 8'b11110010;
  assign _1305_ = state_in[87:80] == 8'b11110001;
  assign _1306_ = state_in[87:80] == 8'b11110000;
  assign _1307_ = state_in[87:80] == 8'b11101111;
  assign _1308_ = state_in[87:80] == 8'b11101110;
  assign _1309_ = state_in[87:80] == 8'b11101101;
  assign _1310_ = state_in[87:80] == 8'b11101100;
  assign _1311_ = state_in[87:80] == 8'b11101011;
  assign _1312_ = state_in[87:80] == 8'b11101010;
  assign _1313_ = state_in[87:80] == 8'b11101001;
  assign _1314_ = state_in[87:80] == 8'b11101000;
  assign _1315_ = state_in[87:80] == 8'b11100111;
  assign _1316_ = state_in[87:80] == 8'b11100110;
  assign _1317_ = state_in[87:80] == 8'b11100101;
  assign _1318_ = state_in[87:80] == 8'b11100100;
  assign _1319_ = state_in[87:80] == 8'b11100011;
  assign _1320_ = state_in[87:80] == 8'b11100010;
  assign _1321_ = state_in[87:80] == 8'b11100001;
  assign _1322_ = state_in[87:80] == 8'b11100000;
  assign _1323_ = state_in[87:80] == 8'b11011111;
  assign _1324_ = state_in[87:80] == 8'b11011110;
  assign _1325_ = state_in[87:80] == 8'b11011101;
  assign _1326_ = state_in[87:80] == 8'b11011100;
  assign _1327_ = state_in[87:80] == 8'b11011011;
  assign _1328_ = state_in[87:80] == 8'b11011010;
  assign _1329_ = state_in[87:80] == 8'b11011001;
  assign _1330_ = state_in[87:80] == 8'b11011000;
  assign _1331_ = state_in[87:80] == 8'b11010111;
  assign _1332_ = state_in[87:80] == 8'b11010110;
  assign _1333_ = state_in[87:80] == 8'b11010101;
  assign _1334_ = state_in[87:80] == 8'b11010100;
  assign _1335_ = state_in[87:80] == 8'b11010011;
  assign _1336_ = state_in[87:80] == 8'b11010010;
  assign _1337_ = state_in[87:80] == 8'b11010001;
  assign _1338_ = state_in[87:80] == 8'b11010000;
  assign _1339_ = state_in[87:80] == 8'b11001111;
  assign _1340_ = state_in[87:80] == 8'b11001110;
  assign _1341_ = state_in[87:80] == 8'b11001101;
  assign _1342_ = state_in[87:80] == 8'b11001100;
  assign _1343_ = state_in[87:80] == 8'b11001011;
  assign _1344_ = state_in[87:80] == 8'b11001010;
  assign _1345_ = state_in[87:80] == 8'b11001001;
  assign _1346_ = state_in[87:80] == 8'b11001000;
  assign _1347_ = state_in[87:80] == 8'b11000111;
  assign _1348_ = state_in[87:80] == 8'b11000110;
  assign _1349_ = state_in[87:80] == 8'b11000101;
  assign _1350_ = state_in[87:80] == 8'b11000100;
  assign _1351_ = state_in[87:80] == 8'b11000011;
  assign _1352_ = state_in[87:80] == 8'b11000010;
  assign _1353_ = state_in[87:80] == 8'b11000001;
  assign _1354_ = state_in[87:80] == 8'b11000000;
  assign _1355_ = state_in[87:80] == 8'b10111111;
  assign _1356_ = state_in[87:80] == 8'b10111110;
  assign _1357_ = state_in[87:80] == 8'b10111101;
  assign _1358_ = state_in[87:80] == 8'b10111100;
  assign _1359_ = state_in[87:80] == 8'b10111011;
  assign _1360_ = state_in[87:80] == 8'b10111010;
  assign _1361_ = state_in[87:80] == 8'b10111001;
  assign _1362_ = state_in[87:80] == 8'b10111000;
  assign _1363_ = state_in[87:80] == 8'b10110111;
  assign _1364_ = state_in[87:80] == 8'b10110110;
  assign _1365_ = state_in[87:80] == 8'b10110101;
  assign _1366_ = state_in[87:80] == 8'b10110100;
  assign _1367_ = state_in[87:80] == 8'b10110011;
  assign _1368_ = state_in[87:80] == 8'b10110010;
  assign _1369_ = state_in[87:80] == 8'b10110001;
  assign _1370_ = state_in[87:80] == 8'b10110000;
  assign _1371_ = state_in[87:80] == 8'b10101111;
  assign _1372_ = state_in[87:80] == 8'b10101110;
  assign _1373_ = state_in[87:80] == 8'b10101101;
  assign _1374_ = state_in[87:80] == 8'b10101100;
  assign _1375_ = state_in[87:80] == 8'b10101011;
  assign _1376_ = state_in[87:80] == 8'b10101010;
  assign _1377_ = state_in[87:80] == 8'b10101001;
  assign _1378_ = state_in[87:80] == 8'b10101000;
  assign _1379_ = state_in[87:80] == 8'b10100111;
  assign _1380_ = state_in[87:80] == 8'b10100110;
  assign _1381_ = state_in[87:80] == 8'b10100101;
  assign _1382_ = state_in[87:80] == 8'b10100100;
  assign _1383_ = state_in[87:80] == 8'b10100011;
  assign _1384_ = state_in[87:80] == 8'b10100010;
  assign _1385_ = state_in[87:80] == 8'b10100001;
  assign _1386_ = state_in[87:80] == 8'b10100000;
  assign _1387_ = state_in[87:80] == 8'b10011111;
  assign _1388_ = state_in[87:80] == 8'b10011110;
  assign _1389_ = state_in[87:80] == 8'b10011101;
  assign _1390_ = state_in[87:80] == 8'b10011100;
  assign _1391_ = state_in[87:80] == 8'b10011011;
  assign _1392_ = state_in[87:80] == 8'b10011010;
  assign _1393_ = state_in[87:80] == 8'b10011001;
  assign _1394_ = state_in[87:80] == 8'b10011000;
  assign _1395_ = state_in[87:80] == 8'b10010111;
  assign _1396_ = state_in[87:80] == 8'b10010110;
  assign _1397_ = state_in[87:80] == 8'b10010101;
  assign _1398_ = state_in[87:80] == 8'b10010100;
  assign _1399_ = state_in[87:80] == 8'b10010011;
  assign _1400_ = state_in[87:80] == 8'b10010010;
  assign _1401_ = state_in[87:80] == 8'b10010001;
  assign _1402_ = state_in[87:80] == 8'b10010000;
  assign _1403_ = state_in[87:80] == 8'b10001111;
  assign _1404_ = state_in[87:80] == 8'b10001110;
  assign _1405_ = state_in[87:80] == 8'b10001101;
  assign _1406_ = state_in[87:80] == 8'b10001100;
  assign _1407_ = state_in[87:80] == 8'b10001011;
  assign _1408_ = state_in[87:80] == 8'b10001010;
  assign _1409_ = state_in[87:80] == 8'b10001001;
  assign _1410_ = state_in[87:80] == 8'b10001000;
  assign _1411_ = state_in[87:80] == 8'b10000111;
  assign _1412_ = state_in[87:80] == 8'b10000110;
  assign _1413_ = state_in[87:80] == 8'b10000101;
  assign _1414_ = state_in[87:80] == 8'b10000100;
  assign _1415_ = state_in[87:80] == 8'b10000011;
  assign _1416_ = state_in[87:80] == 8'b10000010;
  assign _1417_ = state_in[87:80] == 8'b10000001;
  assign _1418_ = state_in[87:80] == 8'b10000000;
  assign _1419_ = state_in[87:80] == 7'b1111111;
  assign _1420_ = state_in[87:80] == 7'b1111110;
  assign _1421_ = state_in[87:80] == 7'b1111101;
  assign _1422_ = state_in[87:80] == 7'b1111100;
  assign _1423_ = state_in[87:80] == 7'b1111011;
  assign _1424_ = state_in[87:80] == 7'b1111010;
  assign _1425_ = state_in[87:80] == 7'b1111001;
  assign _1426_ = state_in[87:80] == 7'b1111000;
  assign _1427_ = state_in[87:80] == 7'b1110111;
  assign _1428_ = state_in[87:80] == 7'b1110110;
  assign _1429_ = state_in[87:80] == 7'b1110101;
  assign _1430_ = state_in[87:80] == 7'b1110100;
  assign _1431_ = state_in[87:80] == 7'b1110011;
  assign _1432_ = state_in[87:80] == 7'b1110010;
  assign _1433_ = state_in[87:80] == 7'b1110001;
  assign _1434_ = state_in[87:80] == 7'b1110000;
  assign _1435_ = state_in[87:80] == 7'b1101111;
  assign _1436_ = state_in[87:80] == 7'b1101110;
  assign _1437_ = state_in[87:80] == 7'b1101101;
  assign _1438_ = state_in[87:80] == 7'b1101100;
  assign _1439_ = state_in[87:80] == 7'b1101011;
  assign _1440_ = state_in[87:80] == 7'b1101010;
  assign _1441_ = state_in[87:80] == 7'b1101001;
  assign _1442_ = state_in[87:80] == 7'b1101000;
  assign _1443_ = state_in[87:80] == 7'b1100111;
  assign _1444_ = state_in[87:80] == 7'b1100110;
  assign _1445_ = state_in[87:80] == 7'b1100101;
  assign _1446_ = state_in[87:80] == 7'b1100100;
  assign _1447_ = state_in[87:80] == 7'b1100011;
  assign _1448_ = state_in[87:80] == 7'b1100010;
  assign _1449_ = state_in[87:80] == 7'b1100001;
  assign _1450_ = state_in[87:80] == 7'b1100000;
  assign _1451_ = state_in[87:80] == 7'b1011111;
  assign _1452_ = state_in[87:80] == 7'b1011110;
  assign _1453_ = state_in[87:80] == 7'b1011101;
  assign _1454_ = state_in[87:80] == 7'b1011100;
  assign _1455_ = state_in[87:80] == 7'b1011011;
  assign _1456_ = state_in[87:80] == 7'b1011010;
  assign _1457_ = state_in[87:80] == 7'b1011001;
  assign _1458_ = state_in[87:80] == 7'b1011000;
  assign _1459_ = state_in[87:80] == 7'b1010111;
  assign _1460_ = state_in[87:80] == 7'b1010110;
  assign _1461_ = state_in[87:80] == 7'b1010101;
  assign _1462_ = state_in[87:80] == 7'b1010100;
  assign _1463_ = state_in[87:80] == 7'b1010011;
  assign _1464_ = state_in[87:80] == 7'b1010010;
  assign _1465_ = state_in[87:80] == 7'b1010001;
  assign _1466_ = state_in[87:80] == 7'b1010000;
  assign _1467_ = state_in[87:80] == 7'b1001111;
  assign _1468_ = state_in[87:80] == 7'b1001110;
  assign _1469_ = state_in[87:80] == 7'b1001101;
  assign _1470_ = state_in[87:80] == 7'b1001100;
  assign _1471_ = state_in[87:80] == 7'b1001011;
  assign _1472_ = state_in[87:80] == 7'b1001010;
  assign _1473_ = state_in[87:80] == 7'b1001001;
  assign _1474_ = state_in[87:80] == 7'b1001000;
  assign _1475_ = state_in[87:80] == 7'b1000111;
  assign _1476_ = state_in[87:80] == 7'b1000110;
  assign _1477_ = state_in[87:80] == 7'b1000101;
  assign _1478_ = state_in[87:80] == 7'b1000100;
  assign _1479_ = state_in[87:80] == 7'b1000011;
  assign _1480_ = state_in[87:80] == 7'b1000010;
  assign _1481_ = state_in[87:80] == 7'b1000001;
  assign _1482_ = state_in[87:80] == 7'b1000000;
  assign _1483_ = state_in[87:80] == 6'b111111;
  assign _1484_ = state_in[87:80] == 6'b111110;
  assign _1485_ = state_in[87:80] == 6'b111101;
  assign _1486_ = state_in[87:80] == 6'b111100;
  assign _1487_ = state_in[87:80] == 6'b111011;
  assign _1488_ = state_in[87:80] == 6'b111010;
  assign _1489_ = state_in[87:80] == 6'b111001;
  assign _1490_ = state_in[87:80] == 6'b111000;
  assign _1491_ = state_in[87:80] == 6'b110111;
  assign _1492_ = state_in[87:80] == 6'b110110;
  assign _1493_ = state_in[87:80] == 6'b110101;
  assign _1494_ = state_in[87:80] == 6'b110100;
  assign _1495_ = state_in[87:80] == 6'b110011;
  assign _1496_ = state_in[87:80] == 6'b110010;
  assign _1497_ = state_in[87:80] == 6'b110001;
  assign _1498_ = state_in[87:80] == 6'b110000;
  assign _1499_ = state_in[87:80] == 6'b101111;
  assign _1500_ = state_in[87:80] == 6'b101110;
  assign _1501_ = state_in[87:80] == 6'b101101;
  assign _1502_ = state_in[87:80] == 6'b101100;
  assign _1503_ = state_in[87:80] == 6'b101011;
  assign _1504_ = state_in[87:80] == 6'b101010;
  assign _1505_ = state_in[87:80] == 6'b101001;
  assign _1506_ = state_in[87:80] == 6'b101000;
  assign _1507_ = state_in[87:80] == 6'b100111;
  assign _1508_ = state_in[87:80] == 6'b100110;
  assign _1509_ = state_in[87:80] == 6'b100101;
  assign _1510_ = state_in[87:80] == 6'b100100;
  assign _1511_ = state_in[87:80] == 6'b100011;
  assign _1512_ = state_in[87:80] == 6'b100010;
  assign _1513_ = state_in[87:80] == 6'b100001;
  assign _1514_ = state_in[87:80] == 6'b100000;
  assign _1515_ = state_in[87:80] == 5'b11111;
  assign _1516_ = state_in[87:80] == 5'b11110;
  assign _1517_ = state_in[87:80] == 5'b11101;
  assign _1518_ = state_in[87:80] == 5'b11100;
  assign _1519_ = state_in[87:80] == 5'b11011;
  assign _1520_ = state_in[87:80] == 5'b11010;
  assign _1521_ = state_in[87:80] == 5'b11001;
  assign _1522_ = state_in[87:80] == 5'b11000;
  assign _1523_ = state_in[87:80] == 5'b10111;
  assign _1524_ = state_in[87:80] == 5'b10110;
  assign _1525_ = state_in[87:80] == 5'b10101;
  assign _1526_ = state_in[87:80] == 5'b10100;
  assign _1527_ = state_in[87:80] == 5'b10011;
  assign _1528_ = state_in[87:80] == 5'b10010;
  assign _1529_ = state_in[87:80] == 5'b10001;
  assign _1530_ = state_in[87:80] == 5'b10000;
  assign _1531_ = state_in[87:80] == 4'b1111;
  assign _1532_ = state_in[87:80] == 4'b1110;
  assign _1533_ = state_in[87:80] == 4'b1101;
  assign _1534_ = state_in[87:80] == 4'b1100;
  assign _1535_ = state_in[87:80] == 4'b1011;
  assign _1536_ = state_in[87:80] == 4'b1010;
  assign _1537_ = state_in[87:80] == 4'b1001;
  assign _1538_ = state_in[87:80] == 4'b1000;
  assign _1539_ = state_in[87:80] == 3'b111;
  assign _1540_ = state_in[87:80] == 3'b110;
  assign _1541_ = state_in[87:80] == 3'b101;
  assign _1542_ = state_in[87:80] == 3'b100;
  assign _1543_ = state_in[87:80] == 2'b11;
  assign _1544_ = state_in[87:80] == 2'b10;
  assign _1545_ = state_in[87:80] == 1'b1;
  assign _1546_ = ! state_in[87:80];
  always @(posedge clk)
      \t1.t1.s4.out <= _1547_;
  logic [255:0] fangyuan12;
  assign fangyuan12 = { _1546_, _1545_, _1544_, _1543_, _1542_, _1541_, _1540_, _1539_, _1538_, _1537_, _1536_, _1535_, _1534_, _1533_, _1532_, _1531_, _1530_, _1529_, _1528_, _1527_, _1526_, _1525_, _1524_, _1523_, _1522_, _1521_, _1520_, _1519_, _1518_, _1517_, _1516_, _1515_, _1514_, _1513_, _1512_, _1511_, _1510_, _1509_, _1508_, _1507_, _1506_, _1505_, _1504_, _1503_, _1502_, _1501_, _1500_, _1499_, _1498_, _1497_, _1496_, _1495_, _1494_, _1493_, _1492_, _1491_, _1490_, _1489_, _1488_, _1487_, _1486_, _1485_, _1484_, _1483_, _1482_, _1481_, _1480_, _1479_, _1478_, _1477_, _1476_, _1475_, _1474_, _1473_, _1472_, _1471_, _1470_, _1469_, _1468_, _1467_, _1466_, _1465_, _1464_, _1463_, _1462_, _1461_, _1460_, _1459_, _1458_, _1457_, _1456_, _1455_, _1454_, _1453_, _1452_, _1451_, _1450_, _1449_, _1448_, _1447_, _1446_, _1445_, _1444_, _1443_, _1442_, _1441_, _1440_, _1439_, _1438_, _1437_, _1436_, _1435_, _1434_, _1433_, _1432_, _1431_, _1430_, _1429_, _1428_, _1427_, _1426_, _1425_, _1424_, _1423_, _1422_, _1421_, _1420_, _1419_, _1418_, _1417_, _1416_, _1415_, _1414_, _1413_, _1412_, _1411_, _1410_, _1409_, _1408_, _1407_, _1406_, _1405_, _1404_, _1403_, _1402_, _1401_, _1400_, _1399_, _1398_, _1397_, _1396_, _1395_, _1394_, _1393_, _1392_, _1391_, _1390_, _1389_, _1388_, _1387_, _1386_, _1385_, _1384_, _1383_, _1382_, _1381_, _1380_, _1379_, _1378_, _1377_, _1376_, _1375_, _1374_, _1373_, _1372_, _1371_, _1370_, _1369_, _1368_, _1367_, _1366_, _1365_, _1364_, _1363_, _1362_, _1361_, _1360_, _1359_, _1358_, _1357_, _1356_, _1355_, _1354_, _1353_, _1352_, _1351_, _1350_, _1349_, _1348_, _1347_, _1346_, _1345_, _1344_, _1343_, _1342_, _1341_, _1340_, _1339_, _1338_, _1337_, _1336_, _1335_, _1334_, _1333_, _1332_, _1331_, _1330_, _1329_, _1328_, _1327_, _1326_, _1325_, _1324_, _1323_, _1322_, _1321_, _1320_, _1319_, _1318_, _1317_, _1316_, _1315_, _1314_, _1313_, _1312_, _1311_, _1310_, _1309_, _1308_, _1307_, _1306_, _1305_, _1304_, _1303_, _1302_, _1301_, _1300_, _1299_, _1298_, _1297_, _1296_, _1295_, _1294_, _1293_, _1292_, _1291_ };

  always @(\t1.t1.s4.out or fangyuan12) begin
    casez (fangyuan12)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1547_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1547_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1547_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1547_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1547_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1547_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1547_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1547_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1547_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1547_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1547_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1547_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1547_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1547_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1547_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1547_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1547_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1547_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1547_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1547_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1547_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1547_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1547_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1547_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1547_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1547_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1547_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1547_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1547_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1547_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1547_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1547_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1547_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1547_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1547_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1547_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1547_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1547_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1547_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1547_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1547_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1547_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1547_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1547_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1547_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1547_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1547_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1547_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1547_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1547_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1547_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1547_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1547_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1547_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1547_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1547_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1547_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1547_ = 8'b11000110 ;
      default:
        _1547_ = \t1.t1.s4.out ;
    endcase
  end
  assign p12[23:16] = \t1.t2.s0.out ^ \t1.t2.s4.out ;
  always @(posedge clk)
      \t1.t2.s0.out <= _1548_;
  logic [255:0] fangyuan13;
  assign fangyuan13 = { _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _1735_, _1734_, _1733_, _1732_, _1731_, _1730_, _1729_, _1728_, _1727_, _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_, _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_ };

  always @(\t1.t2.s0.out or fangyuan13) begin
    casez (fangyuan13)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1548_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1548_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1548_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1548_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1548_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1548_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1548_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1548_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1548_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1548_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1548_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1548_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1548_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1548_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1548_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1548_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1548_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1548_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1548_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1548_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1548_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1548_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1548_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1548_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1548_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1548_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1548_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1548_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1548_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1548_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1548_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1548_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1548_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1548_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1548_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1548_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1548_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1548_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1548_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1548_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1548_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1548_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1548_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1548_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1548_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1548_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1548_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1548_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1548_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1548_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1548_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1548_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1548_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1548_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1548_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1548_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1548_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1548_ = 8'b01100011 ;
      default:
        _1548_ = \t1.t2.s0.out ;
    endcase
  end
  assign _1549_ = state_in[79:72] == 8'b11111111;
  assign _1550_ = state_in[79:72] == 8'b11111110;
  assign _1551_ = state_in[79:72] == 8'b11111101;
  assign _1552_ = state_in[79:72] == 8'b11111100;
  assign _1553_ = state_in[79:72] == 8'b11111011;
  assign _1554_ = state_in[79:72] == 8'b11111010;
  assign _1555_ = state_in[79:72] == 8'b11111001;
  assign _1556_ = state_in[79:72] == 8'b11111000;
  assign _1557_ = state_in[79:72] == 8'b11110111;
  assign _1558_ = state_in[79:72] == 8'b11110110;
  assign _1559_ = state_in[79:72] == 8'b11110101;
  assign _1560_ = state_in[79:72] == 8'b11110100;
  assign _1561_ = state_in[79:72] == 8'b11110011;
  assign _1562_ = state_in[79:72] == 8'b11110010;
  assign _1563_ = state_in[79:72] == 8'b11110001;
  assign _1564_ = state_in[79:72] == 8'b11110000;
  assign _1565_ = state_in[79:72] == 8'b11101111;
  assign _1566_ = state_in[79:72] == 8'b11101110;
  assign _1567_ = state_in[79:72] == 8'b11101101;
  assign _1568_ = state_in[79:72] == 8'b11101100;
  assign _1569_ = state_in[79:72] == 8'b11101011;
  assign _1570_ = state_in[79:72] == 8'b11101010;
  assign _1571_ = state_in[79:72] == 8'b11101001;
  assign _1572_ = state_in[79:72] == 8'b11101000;
  assign _1573_ = state_in[79:72] == 8'b11100111;
  assign _1574_ = state_in[79:72] == 8'b11100110;
  assign _1575_ = state_in[79:72] == 8'b11100101;
  assign _1576_ = state_in[79:72] == 8'b11100100;
  assign _1577_ = state_in[79:72] == 8'b11100011;
  assign _1578_ = state_in[79:72] == 8'b11100010;
  assign _1579_ = state_in[79:72] == 8'b11100001;
  assign _1580_ = state_in[79:72] == 8'b11100000;
  assign _1581_ = state_in[79:72] == 8'b11011111;
  assign _1582_ = state_in[79:72] == 8'b11011110;
  assign _1583_ = state_in[79:72] == 8'b11011101;
  assign _1584_ = state_in[79:72] == 8'b11011100;
  assign _1585_ = state_in[79:72] == 8'b11011011;
  assign _1586_ = state_in[79:72] == 8'b11011010;
  assign _1587_ = state_in[79:72] == 8'b11011001;
  assign _1588_ = state_in[79:72] == 8'b11011000;
  assign _1589_ = state_in[79:72] == 8'b11010111;
  assign _1590_ = state_in[79:72] == 8'b11010110;
  assign _1591_ = state_in[79:72] == 8'b11010101;
  assign _1592_ = state_in[79:72] == 8'b11010100;
  assign _1593_ = state_in[79:72] == 8'b11010011;
  assign _1594_ = state_in[79:72] == 8'b11010010;
  assign _1595_ = state_in[79:72] == 8'b11010001;
  assign _1596_ = state_in[79:72] == 8'b11010000;
  assign _1597_ = state_in[79:72] == 8'b11001111;
  assign _1598_ = state_in[79:72] == 8'b11001110;
  assign _1599_ = state_in[79:72] == 8'b11001101;
  assign _1600_ = state_in[79:72] == 8'b11001100;
  assign _1601_ = state_in[79:72] == 8'b11001011;
  assign _1602_ = state_in[79:72] == 8'b11001010;
  assign _1603_ = state_in[79:72] == 8'b11001001;
  assign _1604_ = state_in[79:72] == 8'b11001000;
  assign _1605_ = state_in[79:72] == 8'b11000111;
  assign _1606_ = state_in[79:72] == 8'b11000110;
  assign _1607_ = state_in[79:72] == 8'b11000101;
  assign _1608_ = state_in[79:72] == 8'b11000100;
  assign _1609_ = state_in[79:72] == 8'b11000011;
  assign _1610_ = state_in[79:72] == 8'b11000010;
  assign _1611_ = state_in[79:72] == 8'b11000001;
  assign _1612_ = state_in[79:72] == 8'b11000000;
  assign _1613_ = state_in[79:72] == 8'b10111111;
  assign _1614_ = state_in[79:72] == 8'b10111110;
  assign _1615_ = state_in[79:72] == 8'b10111101;
  assign _1616_ = state_in[79:72] == 8'b10111100;
  assign _1617_ = state_in[79:72] == 8'b10111011;
  assign _1618_ = state_in[79:72] == 8'b10111010;
  assign _1619_ = state_in[79:72] == 8'b10111001;
  assign _1620_ = state_in[79:72] == 8'b10111000;
  assign _1621_ = state_in[79:72] == 8'b10110111;
  assign _1622_ = state_in[79:72] == 8'b10110110;
  assign _1623_ = state_in[79:72] == 8'b10110101;
  assign _1624_ = state_in[79:72] == 8'b10110100;
  assign _1625_ = state_in[79:72] == 8'b10110011;
  assign _1626_ = state_in[79:72] == 8'b10110010;
  assign _1627_ = state_in[79:72] == 8'b10110001;
  assign _1628_ = state_in[79:72] == 8'b10110000;
  assign _1629_ = state_in[79:72] == 8'b10101111;
  assign _1630_ = state_in[79:72] == 8'b10101110;
  assign _1631_ = state_in[79:72] == 8'b10101101;
  assign _1632_ = state_in[79:72] == 8'b10101100;
  assign _1633_ = state_in[79:72] == 8'b10101011;
  assign _1634_ = state_in[79:72] == 8'b10101010;
  assign _1635_ = state_in[79:72] == 8'b10101001;
  assign _1636_ = state_in[79:72] == 8'b10101000;
  assign _1637_ = state_in[79:72] == 8'b10100111;
  assign _1638_ = state_in[79:72] == 8'b10100110;
  assign _1639_ = state_in[79:72] == 8'b10100101;
  assign _1640_ = state_in[79:72] == 8'b10100100;
  assign _1641_ = state_in[79:72] == 8'b10100011;
  assign _1642_ = state_in[79:72] == 8'b10100010;
  assign _1643_ = state_in[79:72] == 8'b10100001;
  assign _1644_ = state_in[79:72] == 8'b10100000;
  assign _1645_ = state_in[79:72] == 8'b10011111;
  assign _1646_ = state_in[79:72] == 8'b10011110;
  assign _1647_ = state_in[79:72] == 8'b10011101;
  assign _1648_ = state_in[79:72] == 8'b10011100;
  assign _1649_ = state_in[79:72] == 8'b10011011;
  assign _1650_ = state_in[79:72] == 8'b10011010;
  assign _1651_ = state_in[79:72] == 8'b10011001;
  assign _1652_ = state_in[79:72] == 8'b10011000;
  assign _1653_ = state_in[79:72] == 8'b10010111;
  assign _1654_ = state_in[79:72] == 8'b10010110;
  assign _1655_ = state_in[79:72] == 8'b10010101;
  assign _1656_ = state_in[79:72] == 8'b10010100;
  assign _1657_ = state_in[79:72] == 8'b10010011;
  assign _1658_ = state_in[79:72] == 8'b10010010;
  assign _1659_ = state_in[79:72] == 8'b10010001;
  assign _1660_ = state_in[79:72] == 8'b10010000;
  assign _1661_ = state_in[79:72] == 8'b10001111;
  assign _1662_ = state_in[79:72] == 8'b10001110;
  assign _1663_ = state_in[79:72] == 8'b10001101;
  assign _1664_ = state_in[79:72] == 8'b10001100;
  assign _1665_ = state_in[79:72] == 8'b10001011;
  assign _1666_ = state_in[79:72] == 8'b10001010;
  assign _1667_ = state_in[79:72] == 8'b10001001;
  assign _1668_ = state_in[79:72] == 8'b10001000;
  assign _1669_ = state_in[79:72] == 8'b10000111;
  assign _1670_ = state_in[79:72] == 8'b10000110;
  assign _1671_ = state_in[79:72] == 8'b10000101;
  assign _1672_ = state_in[79:72] == 8'b10000100;
  assign _1673_ = state_in[79:72] == 8'b10000011;
  assign _1674_ = state_in[79:72] == 8'b10000010;
  assign _1675_ = state_in[79:72] == 8'b10000001;
  assign _1676_ = state_in[79:72] == 8'b10000000;
  assign _1677_ = state_in[79:72] == 7'b1111111;
  assign _1678_ = state_in[79:72] == 7'b1111110;
  assign _1679_ = state_in[79:72] == 7'b1111101;
  assign _1680_ = state_in[79:72] == 7'b1111100;
  assign _1681_ = state_in[79:72] == 7'b1111011;
  assign _1682_ = state_in[79:72] == 7'b1111010;
  assign _1683_ = state_in[79:72] == 7'b1111001;
  assign _1684_ = state_in[79:72] == 7'b1111000;
  assign _1685_ = state_in[79:72] == 7'b1110111;
  assign _1686_ = state_in[79:72] == 7'b1110110;
  assign _1687_ = state_in[79:72] == 7'b1110101;
  assign _1688_ = state_in[79:72] == 7'b1110100;
  assign _1689_ = state_in[79:72] == 7'b1110011;
  assign _1690_ = state_in[79:72] == 7'b1110010;
  assign _1691_ = state_in[79:72] == 7'b1110001;
  assign _1692_ = state_in[79:72] == 7'b1110000;
  assign _1693_ = state_in[79:72] == 7'b1101111;
  assign _1694_ = state_in[79:72] == 7'b1101110;
  assign _1695_ = state_in[79:72] == 7'b1101101;
  assign _1696_ = state_in[79:72] == 7'b1101100;
  assign _1697_ = state_in[79:72] == 7'b1101011;
  assign _1698_ = state_in[79:72] == 7'b1101010;
  assign _1699_ = state_in[79:72] == 7'b1101001;
  assign _1700_ = state_in[79:72] == 7'b1101000;
  assign _1701_ = state_in[79:72] == 7'b1100111;
  assign _1702_ = state_in[79:72] == 7'b1100110;
  assign _1703_ = state_in[79:72] == 7'b1100101;
  assign _1704_ = state_in[79:72] == 7'b1100100;
  assign _1705_ = state_in[79:72] == 7'b1100011;
  assign _1706_ = state_in[79:72] == 7'b1100010;
  assign _1707_ = state_in[79:72] == 7'b1100001;
  assign _1708_ = state_in[79:72] == 7'b1100000;
  assign _1709_ = state_in[79:72] == 7'b1011111;
  assign _1710_ = state_in[79:72] == 7'b1011110;
  assign _1711_ = state_in[79:72] == 7'b1011101;
  assign _1712_ = state_in[79:72] == 7'b1011100;
  assign _1713_ = state_in[79:72] == 7'b1011011;
  assign _1714_ = state_in[79:72] == 7'b1011010;
  assign _1715_ = state_in[79:72] == 7'b1011001;
  assign _1716_ = state_in[79:72] == 7'b1011000;
  assign _1717_ = state_in[79:72] == 7'b1010111;
  assign _1718_ = state_in[79:72] == 7'b1010110;
  assign _1719_ = state_in[79:72] == 7'b1010101;
  assign _1720_ = state_in[79:72] == 7'b1010100;
  assign _1721_ = state_in[79:72] == 7'b1010011;
  assign _1722_ = state_in[79:72] == 7'b1010010;
  assign _1723_ = state_in[79:72] == 7'b1010001;
  assign _1724_ = state_in[79:72] == 7'b1010000;
  assign _1725_ = state_in[79:72] == 7'b1001111;
  assign _1726_ = state_in[79:72] == 7'b1001110;
  assign _1727_ = state_in[79:72] == 7'b1001101;
  assign _1728_ = state_in[79:72] == 7'b1001100;
  assign _1729_ = state_in[79:72] == 7'b1001011;
  assign _1730_ = state_in[79:72] == 7'b1001010;
  assign _1731_ = state_in[79:72] == 7'b1001001;
  assign _1732_ = state_in[79:72] == 7'b1001000;
  assign _1733_ = state_in[79:72] == 7'b1000111;
  assign _1734_ = state_in[79:72] == 7'b1000110;
  assign _1735_ = state_in[79:72] == 7'b1000101;
  assign _1736_ = state_in[79:72] == 7'b1000100;
  assign _1737_ = state_in[79:72] == 7'b1000011;
  assign _1738_ = state_in[79:72] == 7'b1000010;
  assign _1739_ = state_in[79:72] == 7'b1000001;
  assign _1740_ = state_in[79:72] == 7'b1000000;
  assign _1741_ = state_in[79:72] == 6'b111111;
  assign _1742_ = state_in[79:72] == 6'b111110;
  assign _1743_ = state_in[79:72] == 6'b111101;
  assign _1744_ = state_in[79:72] == 6'b111100;
  assign _1745_ = state_in[79:72] == 6'b111011;
  assign _1746_ = state_in[79:72] == 6'b111010;
  assign _1747_ = state_in[79:72] == 6'b111001;
  assign _1748_ = state_in[79:72] == 6'b111000;
  assign _1749_ = state_in[79:72] == 6'b110111;
  assign _1750_ = state_in[79:72] == 6'b110110;
  assign _1751_ = state_in[79:72] == 6'b110101;
  assign _1752_ = state_in[79:72] == 6'b110100;
  assign _1753_ = state_in[79:72] == 6'b110011;
  assign _1754_ = state_in[79:72] == 6'b110010;
  assign _1755_ = state_in[79:72] == 6'b110001;
  assign _1756_ = state_in[79:72] == 6'b110000;
  assign _1757_ = state_in[79:72] == 6'b101111;
  assign _1758_ = state_in[79:72] == 6'b101110;
  assign _1759_ = state_in[79:72] == 6'b101101;
  assign _1760_ = state_in[79:72] == 6'b101100;
  assign _1761_ = state_in[79:72] == 6'b101011;
  assign _1762_ = state_in[79:72] == 6'b101010;
  assign _1763_ = state_in[79:72] == 6'b101001;
  assign _1764_ = state_in[79:72] == 6'b101000;
  assign _1765_ = state_in[79:72] == 6'b100111;
  assign _1766_ = state_in[79:72] == 6'b100110;
  assign _1767_ = state_in[79:72] == 6'b100101;
  assign _1768_ = state_in[79:72] == 6'b100100;
  assign _1769_ = state_in[79:72] == 6'b100011;
  assign _1770_ = state_in[79:72] == 6'b100010;
  assign _1771_ = state_in[79:72] == 6'b100001;
  assign _1772_ = state_in[79:72] == 6'b100000;
  assign _1773_ = state_in[79:72] == 5'b11111;
  assign _1774_ = state_in[79:72] == 5'b11110;
  assign _1775_ = state_in[79:72] == 5'b11101;
  assign _1776_ = state_in[79:72] == 5'b11100;
  assign _1777_ = state_in[79:72] == 5'b11011;
  assign _1778_ = state_in[79:72] == 5'b11010;
  assign _1779_ = state_in[79:72] == 5'b11001;
  assign _1780_ = state_in[79:72] == 5'b11000;
  assign _1781_ = state_in[79:72] == 5'b10111;
  assign _1782_ = state_in[79:72] == 5'b10110;
  assign _1783_ = state_in[79:72] == 5'b10101;
  assign _1784_ = state_in[79:72] == 5'b10100;
  assign _1785_ = state_in[79:72] == 5'b10011;
  assign _1786_ = state_in[79:72] == 5'b10010;
  assign _1787_ = state_in[79:72] == 5'b10001;
  assign _1788_ = state_in[79:72] == 5'b10000;
  assign _1789_ = state_in[79:72] == 4'b1111;
  assign _1790_ = state_in[79:72] == 4'b1110;
  assign _1791_ = state_in[79:72] == 4'b1101;
  assign _1792_ = state_in[79:72] == 4'b1100;
  assign _1793_ = state_in[79:72] == 4'b1011;
  assign _1794_ = state_in[79:72] == 4'b1010;
  assign _1795_ = state_in[79:72] == 4'b1001;
  assign _1796_ = state_in[79:72] == 4'b1000;
  assign _1797_ = state_in[79:72] == 3'b111;
  assign _1798_ = state_in[79:72] == 3'b110;
  assign _1799_ = state_in[79:72] == 3'b101;
  assign _1800_ = state_in[79:72] == 3'b100;
  assign _1801_ = state_in[79:72] == 2'b11;
  assign _1802_ = state_in[79:72] == 2'b10;
  assign _1803_ = state_in[79:72] == 1'b1;
  assign _1804_ = ! state_in[79:72];
  always @(posedge clk)
      \t1.t2.s4.out <= _1805_;
  logic [255:0] fangyuan14;
  assign fangyuan14 = { _1804_, _1803_, _1802_, _1801_, _1800_, _1799_, _1798_, _1797_, _1796_, _1795_, _1794_, _1793_, _1792_, _1791_, _1790_, _1789_, _1788_, _1787_, _1786_, _1785_, _1784_, _1783_, _1782_, _1781_, _1780_, _1779_, _1778_, _1777_, _1776_, _1775_, _1774_, _1773_, _1772_, _1771_, _1770_, _1769_, _1768_, _1767_, _1766_, _1765_, _1764_, _1763_, _1762_, _1761_, _1760_, _1759_, _1758_, _1757_, _1756_, _1755_, _1754_, _1753_, _1752_, _1751_, _1750_, _1749_, _1748_, _1747_, _1746_, _1745_, _1744_, _1743_, _1742_, _1741_, _1740_, _1739_, _1738_, _1737_, _1736_, _1735_, _1734_, _1733_, _1732_, _1731_, _1730_, _1729_, _1728_, _1727_, _1726_, _1725_, _1724_, _1723_, _1722_, _1721_, _1720_, _1719_, _1718_, _1717_, _1716_, _1715_, _1714_, _1713_, _1712_, _1711_, _1710_, _1709_, _1708_, _1707_, _1706_, _1705_, _1704_, _1703_, _1702_, _1701_, _1700_, _1699_, _1698_, _1697_, _1696_, _1695_, _1694_, _1693_, _1692_, _1691_, _1690_, _1689_, _1688_, _1687_, _1686_, _1685_, _1684_, _1683_, _1682_, _1681_, _1680_, _1679_, _1678_, _1677_, _1676_, _1675_, _1674_, _1673_, _1672_, _1671_, _1670_, _1669_, _1668_, _1667_, _1666_, _1665_, _1664_, _1663_, _1662_, _1661_, _1660_, _1659_, _1658_, _1657_, _1656_, _1655_, _1654_, _1653_, _1652_, _1651_, _1650_, _1649_, _1648_, _1647_, _1646_, _1645_, _1644_, _1643_, _1642_, _1641_, _1640_, _1639_, _1638_, _1637_, _1636_, _1635_, _1634_, _1633_, _1632_, _1631_, _1630_, _1629_, _1628_, _1627_, _1626_, _1625_, _1624_, _1623_, _1622_, _1621_, _1620_, _1619_, _1618_, _1617_, _1616_, _1615_, _1614_, _1613_, _1612_, _1611_, _1610_, _1609_, _1608_, _1607_, _1606_, _1605_, _1604_, _1603_, _1602_, _1601_, _1600_, _1599_, _1598_, _1597_, _1596_, _1595_, _1594_, _1593_, _1592_, _1591_, _1590_, _1589_, _1588_, _1587_, _1586_, _1585_, _1584_, _1583_, _1582_, _1581_, _1580_, _1579_, _1578_, _1577_, _1576_, _1575_, _1574_, _1573_, _1572_, _1571_, _1570_, _1569_, _1568_, _1567_, _1566_, _1565_, _1564_, _1563_, _1562_, _1561_, _1560_, _1559_, _1558_, _1557_, _1556_, _1555_, _1554_, _1553_, _1552_, _1551_, _1550_, _1549_ };

  always @(\t1.t2.s4.out or fangyuan14) begin
    casez (fangyuan14)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1805_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1805_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1805_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1805_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1805_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1805_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1805_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1805_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1805_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1805_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1805_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1805_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1805_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1805_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1805_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1805_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1805_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1805_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1805_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1805_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1805_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1805_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1805_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1805_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1805_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1805_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1805_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1805_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1805_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1805_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1805_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1805_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1805_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1805_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1805_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1805_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1805_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1805_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1805_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1805_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1805_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1805_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1805_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1805_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1805_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1805_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1805_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1805_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1805_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1805_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1805_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1805_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1805_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1805_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1805_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1805_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1805_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1805_ = 8'b11000110 ;
      default:
        _1805_ = \t1.t2.s4.out ;
    endcase
  end
  assign p13[15:8] = \t1.t3.s0.out ^ \t1.t3.s4.out ;
  always @(posedge clk)
      \t1.t3.s0.out <= _1806_;
  logic [255:0] fangyuan15;
  assign fangyuan15 = { _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _1998_, _1997_, _1996_, _1995_, _1994_, _1993_, _1992_, _1991_, _1990_, _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_, _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_ };

  always @(\t1.t3.s0.out or fangyuan15) begin
    casez (fangyuan15)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _1806_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _1806_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _1806_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _1806_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _1806_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _1806_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _1806_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _1806_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _1806_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _1806_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _1806_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _1806_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _1806_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _1806_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _1806_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _1806_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _1806_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _1806_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _1806_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _1806_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _1806_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _1806_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _1806_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _1806_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _1806_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _1806_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _1806_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _1806_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _1806_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _1806_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _1806_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _1806_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _1806_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _1806_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _1806_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _1806_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _1806_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _1806_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _1806_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _1806_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _1806_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _1806_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _1806_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _1806_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _1806_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _1806_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _1806_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _1806_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _1806_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _1806_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _1806_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _1806_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _1806_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _1806_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _1806_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _1806_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _1806_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _1806_ = 8'b01100011 ;
      default:
        _1806_ = \t1.t3.s0.out ;
    endcase
  end
  assign _1807_ = state_in[71:64] == 8'b11111111;
  assign _1808_ = state_in[71:64] == 8'b11111110;
  assign _1809_ = state_in[71:64] == 8'b11111101;
  assign _1810_ = state_in[71:64] == 8'b11111100;
  assign _1811_ = state_in[71:64] == 8'b11111011;
  assign _1812_ = state_in[71:64] == 8'b11111010;
  assign _1813_ = state_in[71:64] == 8'b11111001;
  assign _1814_ = state_in[71:64] == 8'b11111000;
  assign _1815_ = state_in[71:64] == 8'b11110111;
  assign _1816_ = state_in[71:64] == 8'b11110110;
  assign _1817_ = state_in[71:64] == 8'b11110101;
  assign _1818_ = state_in[71:64] == 8'b11110100;
  assign _1819_ = state_in[71:64] == 8'b11110011;
  assign _1820_ = state_in[71:64] == 8'b11110010;
  assign _1821_ = state_in[71:64] == 8'b11110001;
  assign _1822_ = state_in[71:64] == 8'b11110000;
  assign _1823_ = state_in[71:64] == 8'b11101111;
  assign _1824_ = state_in[71:64] == 8'b11101110;
  assign _1825_ = state_in[71:64] == 8'b11101101;
  assign _1826_ = state_in[71:64] == 8'b11101100;
  assign _1827_ = state_in[71:64] == 8'b11101011;
  assign _1828_ = state_in[71:64] == 8'b11101010;
  assign _1829_ = state_in[71:64] == 8'b11101001;
  assign _1830_ = state_in[71:64] == 8'b11101000;
  assign _1831_ = state_in[71:64] == 8'b11100111;
  assign _1832_ = state_in[71:64] == 8'b11100110;
  assign _1833_ = state_in[71:64] == 8'b11100101;
  assign _1834_ = state_in[71:64] == 8'b11100100;
  assign _1835_ = state_in[71:64] == 8'b11100011;
  assign _1836_ = state_in[71:64] == 8'b11100010;
  assign _1837_ = state_in[71:64] == 8'b11100001;
  assign _1838_ = state_in[71:64] == 8'b11100000;
  assign _1839_ = state_in[71:64] == 8'b11011111;
  assign _1840_ = state_in[71:64] == 8'b11011110;
  assign _1841_ = state_in[71:64] == 8'b11011101;
  assign _1842_ = state_in[71:64] == 8'b11011100;
  assign _1843_ = state_in[71:64] == 8'b11011011;
  assign _1844_ = state_in[71:64] == 8'b11011010;
  assign _1845_ = state_in[71:64] == 8'b11011001;
  assign _1846_ = state_in[71:64] == 8'b11011000;
  assign _1847_ = state_in[71:64] == 8'b11010111;
  assign _1848_ = state_in[71:64] == 8'b11010110;
  assign _1849_ = state_in[71:64] == 8'b11010101;
  assign _1850_ = state_in[71:64] == 8'b11010100;
  assign _1851_ = state_in[71:64] == 8'b11010011;
  assign _1852_ = state_in[71:64] == 8'b11010010;
  assign _1853_ = state_in[71:64] == 8'b11010001;
  assign _1854_ = state_in[71:64] == 8'b11010000;
  assign _1855_ = state_in[71:64] == 8'b11001111;
  assign _1856_ = state_in[71:64] == 8'b11001110;
  assign _1857_ = state_in[71:64] == 8'b11001101;
  assign _1858_ = state_in[71:64] == 8'b11001100;
  assign _1859_ = state_in[71:64] == 8'b11001011;
  assign _1860_ = state_in[71:64] == 8'b11001010;
  assign _1861_ = state_in[71:64] == 8'b11001001;
  assign _1862_ = state_in[71:64] == 8'b11001000;
  assign _1863_ = state_in[71:64] == 8'b11000111;
  assign _1864_ = state_in[71:64] == 8'b11000110;
  assign _1865_ = state_in[71:64] == 8'b11000101;
  assign _1866_ = state_in[71:64] == 8'b11000100;
  assign _1867_ = state_in[71:64] == 8'b11000011;
  assign _1868_ = state_in[71:64] == 8'b11000010;
  assign _1869_ = state_in[71:64] == 8'b11000001;
  assign _1870_ = state_in[71:64] == 8'b11000000;
  assign _1871_ = state_in[71:64] == 8'b10111111;
  assign _1872_ = state_in[71:64] == 8'b10111110;
  assign _1873_ = state_in[71:64] == 8'b10111101;
  assign _1874_ = state_in[71:64] == 8'b10111100;
  assign _1875_ = state_in[71:64] == 8'b10111011;
  assign _1876_ = state_in[71:64] == 8'b10111010;
  assign _1877_ = state_in[71:64] == 8'b10111001;
  assign _1878_ = state_in[71:64] == 8'b10111000;
  assign _1879_ = state_in[71:64] == 8'b10110111;
  assign _1880_ = state_in[71:64] == 8'b10110110;
  assign _1881_ = state_in[71:64] == 8'b10110101;
  assign _1882_ = state_in[71:64] == 8'b10110100;
  assign _1883_ = state_in[71:64] == 8'b10110011;
  assign _1884_ = state_in[71:64] == 8'b10110010;
  assign _1885_ = state_in[71:64] == 8'b10110001;
  assign _1886_ = state_in[71:64] == 8'b10110000;
  assign _1887_ = state_in[71:64] == 8'b10101111;
  assign _1888_ = state_in[71:64] == 8'b10101110;
  assign _1889_ = state_in[71:64] == 8'b10101101;
  assign _1890_ = state_in[71:64] == 8'b10101100;
  assign _1891_ = state_in[71:64] == 8'b10101011;
  assign _1892_ = state_in[71:64] == 8'b10101010;
  assign _1893_ = state_in[71:64] == 8'b10101001;
  assign _1894_ = state_in[71:64] == 8'b10101000;
  assign _1895_ = state_in[71:64] == 8'b10100111;
  assign _1896_ = state_in[71:64] == 8'b10100110;
  assign _1897_ = state_in[71:64] == 8'b10100101;
  assign _1898_ = state_in[71:64] == 8'b10100100;
  assign _1899_ = state_in[71:64] == 8'b10100011;
  assign _1900_ = state_in[71:64] == 8'b10100010;
  assign _1901_ = state_in[71:64] == 8'b10100001;
  assign _1902_ = state_in[71:64] == 8'b10100000;
  assign _1903_ = state_in[71:64] == 8'b10011111;
  assign _1904_ = state_in[71:64] == 8'b10011110;
  assign _1905_ = state_in[71:64] == 8'b10011101;
  assign _1906_ = state_in[71:64] == 8'b10011100;
  assign _1907_ = state_in[71:64] == 8'b10011011;
  assign _1908_ = state_in[71:64] == 8'b10011010;
  assign _1909_ = state_in[71:64] == 8'b10011001;
  assign _1910_ = state_in[71:64] == 8'b10011000;
  assign _1911_ = state_in[71:64] == 8'b10010111;
  assign _1912_ = state_in[71:64] == 8'b10010110;
  assign _1913_ = state_in[71:64] == 8'b10010101;
  assign _1914_ = state_in[71:64] == 8'b10010100;
  assign _1915_ = state_in[71:64] == 8'b10010011;
  assign _1916_ = state_in[71:64] == 8'b10010010;
  assign _1917_ = state_in[71:64] == 8'b10010001;
  assign _1918_ = state_in[71:64] == 8'b10010000;
  assign _1919_ = state_in[71:64] == 8'b10001111;
  assign _1920_ = state_in[71:64] == 8'b10001110;
  assign _1921_ = state_in[71:64] == 8'b10001101;
  assign _1922_ = state_in[71:64] == 8'b10001100;
  assign _1923_ = state_in[71:64] == 8'b10001011;
  assign _1924_ = state_in[71:64] == 8'b10001010;
  assign _1925_ = state_in[71:64] == 8'b10001001;
  assign _1926_ = state_in[71:64] == 8'b10001000;
  assign _1927_ = state_in[71:64] == 8'b10000111;
  assign _1928_ = state_in[71:64] == 8'b10000110;
  assign _1929_ = state_in[71:64] == 8'b10000101;
  assign _1930_ = state_in[71:64] == 8'b10000100;
  assign _1931_ = state_in[71:64] == 8'b10000011;
  assign _1932_ = state_in[71:64] == 8'b10000010;
  assign _1933_ = state_in[71:64] == 8'b10000001;
  assign _1934_ = state_in[71:64] == 8'b10000000;
  assign _1935_ = state_in[71:64] == 7'b1111111;
  assign _1936_ = state_in[71:64] == 7'b1111110;
  assign _1937_ = state_in[71:64] == 7'b1111101;
  assign _1938_ = state_in[71:64] == 7'b1111100;
  assign _1939_ = state_in[71:64] == 7'b1111011;
  assign _1940_ = state_in[71:64] == 7'b1111010;
  assign _1941_ = state_in[71:64] == 7'b1111001;
  assign _1942_ = state_in[71:64] == 7'b1111000;
  assign _1943_ = state_in[71:64] == 7'b1110111;
  assign _1944_ = state_in[71:64] == 7'b1110110;
  assign _1945_ = state_in[71:64] == 7'b1110101;
  assign _1946_ = state_in[71:64] == 7'b1110100;
  assign _1947_ = state_in[71:64] == 7'b1110011;
  assign _1948_ = state_in[71:64] == 7'b1110010;
  assign _1949_ = state_in[71:64] == 7'b1110001;
  assign _1950_ = state_in[71:64] == 7'b1110000;
  assign _1951_ = state_in[71:64] == 7'b1101111;
  assign _1952_ = state_in[71:64] == 7'b1101110;
  assign _1953_ = state_in[71:64] == 7'b1101101;
  assign _1954_ = state_in[71:64] == 7'b1101100;
  assign _1955_ = state_in[71:64] == 7'b1101011;
  assign _1956_ = state_in[71:64] == 7'b1101010;
  assign _1957_ = state_in[71:64] == 7'b1101001;
  assign _1958_ = state_in[71:64] == 7'b1101000;
  assign _1959_ = state_in[71:64] == 7'b1100111;
  assign _1960_ = state_in[71:64] == 7'b1100110;
  assign _1961_ = state_in[71:64] == 7'b1100101;
  assign _1962_ = state_in[71:64] == 7'b1100100;
  assign _1963_ = state_in[71:64] == 7'b1100011;
  assign _1964_ = state_in[71:64] == 7'b1100010;
  assign _1965_ = state_in[71:64] == 7'b1100001;
  assign _1966_ = state_in[71:64] == 7'b1100000;
  assign _1967_ = state_in[71:64] == 7'b1011111;
  assign _1968_ = state_in[71:64] == 7'b1011110;
  assign _1969_ = state_in[71:64] == 7'b1011101;
  assign _1970_ = state_in[71:64] == 7'b1011100;
  assign _1971_ = state_in[71:64] == 7'b1011011;
  assign _1972_ = state_in[71:64] == 7'b1011010;
  assign _1973_ = state_in[71:64] == 7'b1011001;
  assign _1974_ = state_in[71:64] == 7'b1011000;
  assign _1975_ = state_in[71:64] == 7'b1010111;
  assign _1976_ = state_in[71:64] == 7'b1010110;
  assign _1977_ = state_in[71:64] == 7'b1010101;
  assign _1978_ = state_in[71:64] == 7'b1010100;
  assign _1979_ = state_in[71:64] == 7'b1010011;
  assign _1980_ = state_in[71:64] == 7'b1010010;
  assign _1981_ = state_in[71:64] == 7'b1010001;
  assign _1982_ = state_in[71:64] == 7'b1010000;
  assign _1983_ = state_in[71:64] == 7'b1001111;
  assign _1984_ = state_in[71:64] == 7'b1001110;
  assign _1985_ = state_in[71:64] == 7'b1001101;
  assign _1986_ = state_in[71:64] == 7'b1001100;
  assign _1987_ = state_in[71:64] == 7'b1001011;
  assign _1988_ = state_in[71:64] == 7'b1001010;
  assign _1989_ = state_in[71:64] == 7'b1001001;
  assign _1990_ = state_in[71:64] == 7'b1001000;
  assign _1991_ = state_in[71:64] == 7'b1000111;
  assign _1992_ = state_in[71:64] == 7'b1000110;
  assign _1993_ = state_in[71:64] == 7'b1000101;
  assign _1994_ = state_in[71:64] == 7'b1000100;
  assign _1995_ = state_in[71:64] == 7'b1000011;
  assign _1996_ = state_in[71:64] == 7'b1000010;
  assign _1997_ = state_in[71:64] == 7'b1000001;
  assign _1998_ = state_in[71:64] == 7'b1000000;
  assign _1999_ = state_in[71:64] == 6'b111111;
  assign _2000_ = state_in[71:64] == 6'b111110;
  assign _2001_ = state_in[71:64] == 6'b111101;
  assign _2002_ = state_in[71:64] == 6'b111100;
  assign _2003_ = state_in[71:64] == 6'b111011;
  assign _2004_ = state_in[71:64] == 6'b111010;
  assign _2005_ = state_in[71:64] == 6'b111001;
  assign _2006_ = state_in[71:64] == 6'b111000;
  assign _2007_ = state_in[71:64] == 6'b110111;
  assign _2008_ = state_in[71:64] == 6'b110110;
  assign _2009_ = state_in[71:64] == 6'b110101;
  assign _2010_ = state_in[71:64] == 6'b110100;
  assign _2011_ = state_in[71:64] == 6'b110011;
  assign _2012_ = state_in[71:64] == 6'b110010;
  assign _2013_ = state_in[71:64] == 6'b110001;
  assign _2014_ = state_in[71:64] == 6'b110000;
  assign _2015_ = state_in[71:64] == 6'b101111;
  assign _2016_ = state_in[71:64] == 6'b101110;
  assign _2017_ = state_in[71:64] == 6'b101101;
  assign _2018_ = state_in[71:64] == 6'b101100;
  assign _2019_ = state_in[71:64] == 6'b101011;
  assign _2020_ = state_in[71:64] == 6'b101010;
  assign _2021_ = state_in[71:64] == 6'b101001;
  assign _2022_ = state_in[71:64] == 6'b101000;
  assign _2023_ = state_in[71:64] == 6'b100111;
  assign _2024_ = state_in[71:64] == 6'b100110;
  assign _2025_ = state_in[71:64] == 6'b100101;
  assign _2026_ = state_in[71:64] == 6'b100100;
  assign _2027_ = state_in[71:64] == 6'b100011;
  assign _2028_ = state_in[71:64] == 6'b100010;
  assign _2029_ = state_in[71:64] == 6'b100001;
  assign _2030_ = state_in[71:64] == 6'b100000;
  assign _2031_ = state_in[71:64] == 5'b11111;
  assign _2032_ = state_in[71:64] == 5'b11110;
  assign _2033_ = state_in[71:64] == 5'b11101;
  assign _2034_ = state_in[71:64] == 5'b11100;
  assign _2035_ = state_in[71:64] == 5'b11011;
  assign _2036_ = state_in[71:64] == 5'b11010;
  assign _2037_ = state_in[71:64] == 5'b11001;
  assign _2038_ = state_in[71:64] == 5'b11000;
  assign _2039_ = state_in[71:64] == 5'b10111;
  assign _2040_ = state_in[71:64] == 5'b10110;
  assign _2041_ = state_in[71:64] == 5'b10101;
  assign _2042_ = state_in[71:64] == 5'b10100;
  assign _2043_ = state_in[71:64] == 5'b10011;
  assign _2044_ = state_in[71:64] == 5'b10010;
  assign _2045_ = state_in[71:64] == 5'b10001;
  assign _2046_ = state_in[71:64] == 5'b10000;
  assign _2047_ = state_in[71:64] == 4'b1111;
  assign _2048_ = state_in[71:64] == 4'b1110;
  assign _2049_ = state_in[71:64] == 4'b1101;
  assign _2050_ = state_in[71:64] == 4'b1100;
  assign _2051_ = state_in[71:64] == 4'b1011;
  assign _2052_ = state_in[71:64] == 4'b1010;
  assign _2053_ = state_in[71:64] == 4'b1001;
  assign _2054_ = state_in[71:64] == 4'b1000;
  assign _2055_ = state_in[71:64] == 3'b111;
  assign _2056_ = state_in[71:64] == 3'b110;
  assign _2057_ = state_in[71:64] == 3'b101;
  assign _2058_ = state_in[71:64] == 3'b100;
  assign _2059_ = state_in[71:64] == 2'b11;
  assign _2060_ = state_in[71:64] == 2'b10;
  assign _2061_ = state_in[71:64] == 1'b1;
  assign _2062_ = ! state_in[71:64];
  always @(posedge clk)
      \t1.t3.s4.out <= _2063_;
  logic [255:0] fangyuan16;
  assign fangyuan16 = { _2062_, _2061_, _2060_, _2059_, _2058_, _2057_, _2056_, _2055_, _2054_, _2053_, _2052_, _2051_, _2050_, _2049_, _2048_, _2047_, _2046_, _2045_, _2044_, _2043_, _2042_, _2041_, _2040_, _2039_, _2038_, _2037_, _2036_, _2035_, _2034_, _2033_, _2032_, _2031_, _2030_, _2029_, _2028_, _2027_, _2026_, _2025_, _2024_, _2023_, _2022_, _2021_, _2020_, _2019_, _2018_, _2017_, _2016_, _2015_, _2014_, _2013_, _2012_, _2011_, _2010_, _2009_, _2008_, _2007_, _2006_, _2005_, _2004_, _2003_, _2002_, _2001_, _2000_, _1999_, _1998_, _1997_, _1996_, _1995_, _1994_, _1993_, _1992_, _1991_, _1990_, _1989_, _1988_, _1987_, _1986_, _1985_, _1984_, _1983_, _1982_, _1981_, _1980_, _1979_, _1978_, _1977_, _1976_, _1975_, _1974_, _1973_, _1972_, _1971_, _1970_, _1969_, _1968_, _1967_, _1966_, _1965_, _1964_, _1963_, _1962_, _1961_, _1960_, _1959_, _1958_, _1957_, _1956_, _1955_, _1954_, _1953_, _1952_, _1951_, _1950_, _1949_, _1948_, _1947_, _1946_, _1945_, _1944_, _1943_, _1942_, _1941_, _1940_, _1939_, _1938_, _1937_, _1936_, _1935_, _1934_, _1933_, _1932_, _1931_, _1930_, _1929_, _1928_, _1927_, _1926_, _1925_, _1924_, _1923_, _1922_, _1921_, _1920_, _1919_, _1918_, _1917_, _1916_, _1915_, _1914_, _1913_, _1912_, _1911_, _1910_, _1909_, _1908_, _1907_, _1906_, _1905_, _1904_, _1903_, _1902_, _1901_, _1900_, _1899_, _1898_, _1897_, _1896_, _1895_, _1894_, _1893_, _1892_, _1891_, _1890_, _1889_, _1888_, _1887_, _1886_, _1885_, _1884_, _1883_, _1882_, _1881_, _1880_, _1879_, _1878_, _1877_, _1876_, _1875_, _1874_, _1873_, _1872_, _1871_, _1870_, _1869_, _1868_, _1867_, _1866_, _1865_, _1864_, _1863_, _1862_, _1861_, _1860_, _1859_, _1858_, _1857_, _1856_, _1855_, _1854_, _1853_, _1852_, _1851_, _1850_, _1849_, _1848_, _1847_, _1846_, _1845_, _1844_, _1843_, _1842_, _1841_, _1840_, _1839_, _1838_, _1837_, _1836_, _1835_, _1834_, _1833_, _1832_, _1831_, _1830_, _1829_, _1828_, _1827_, _1826_, _1825_, _1824_, _1823_, _1822_, _1821_, _1820_, _1819_, _1818_, _1817_, _1816_, _1815_, _1814_, _1813_, _1812_, _1811_, _1810_, _1809_, _1808_, _1807_ };

  always @(\t1.t3.s4.out or fangyuan16) begin
    casez (fangyuan16)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2063_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2063_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2063_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2063_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2063_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2063_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2063_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2063_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2063_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2063_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2063_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2063_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2063_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2063_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2063_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2063_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2063_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2063_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2063_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2063_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2063_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2063_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2063_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2063_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2063_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2063_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2063_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2063_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2063_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2063_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2063_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2063_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2063_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2063_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2063_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2063_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2063_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2063_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2063_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2063_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2063_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2063_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2063_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2063_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2063_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2063_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2063_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2063_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2063_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2063_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2063_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2063_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2063_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2063_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2063_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2063_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2063_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2063_ = 8'b11000110 ;
      default:
        _2063_ = \t1.t3.s4.out ;
    endcase
  end
  assign p20[7:0] = \t2.t0.s0.out ^ \t2.t0.s4.out ;
  always @(posedge clk)
      \t2.t0.s0.out <= _2064_;
  logic [255:0] fangyuan17;
  assign fangyuan17 = { _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _2261_, _2260_, _2259_, _2258_, _2257_, _2256_, _2255_, _2254_, _2253_, _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_, _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_ };

  always @(\t2.t0.s0.out or fangyuan17) begin
    casez (fangyuan17)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2064_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2064_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2064_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2064_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2064_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2064_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2064_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2064_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2064_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2064_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2064_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2064_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2064_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2064_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2064_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2064_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2064_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2064_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2064_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2064_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2064_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2064_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2064_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2064_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2064_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2064_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2064_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2064_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2064_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2064_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2064_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2064_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2064_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2064_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2064_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2064_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2064_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2064_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2064_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2064_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2064_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2064_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2064_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2064_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2064_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2064_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2064_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2064_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2064_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2064_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2064_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2064_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2064_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2064_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2064_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2064_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2064_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2064_ = 8'b01100011 ;
      default:
        _2064_ = \t2.t0.s0.out ;
    endcase
  end
  assign _2065_ = state_in[63:56] == 8'b11111111;
  assign _2066_ = state_in[63:56] == 8'b11111110;
  assign _2067_ = state_in[63:56] == 8'b11111101;
  assign _2068_ = state_in[63:56] == 8'b11111100;
  assign _2069_ = state_in[63:56] == 8'b11111011;
  assign _2070_ = state_in[63:56] == 8'b11111010;
  assign _2071_ = state_in[63:56] == 8'b11111001;
  assign _2072_ = state_in[63:56] == 8'b11111000;
  assign _2073_ = state_in[63:56] == 8'b11110111;
  assign _2074_ = state_in[63:56] == 8'b11110110;
  assign _2075_ = state_in[63:56] == 8'b11110101;
  assign _2076_ = state_in[63:56] == 8'b11110100;
  assign _2077_ = state_in[63:56] == 8'b11110011;
  assign _2078_ = state_in[63:56] == 8'b11110010;
  assign _2079_ = state_in[63:56] == 8'b11110001;
  assign _2080_ = state_in[63:56] == 8'b11110000;
  assign _2081_ = state_in[63:56] == 8'b11101111;
  assign _2082_ = state_in[63:56] == 8'b11101110;
  assign _2083_ = state_in[63:56] == 8'b11101101;
  assign _2084_ = state_in[63:56] == 8'b11101100;
  assign _2085_ = state_in[63:56] == 8'b11101011;
  assign _2086_ = state_in[63:56] == 8'b11101010;
  assign _2087_ = state_in[63:56] == 8'b11101001;
  assign _2088_ = state_in[63:56] == 8'b11101000;
  assign _2089_ = state_in[63:56] == 8'b11100111;
  assign _2090_ = state_in[63:56] == 8'b11100110;
  assign _2091_ = state_in[63:56] == 8'b11100101;
  assign _2092_ = state_in[63:56] == 8'b11100100;
  assign _2093_ = state_in[63:56] == 8'b11100011;
  assign _2094_ = state_in[63:56] == 8'b11100010;
  assign _2095_ = state_in[63:56] == 8'b11100001;
  assign _2096_ = state_in[63:56] == 8'b11100000;
  assign _2097_ = state_in[63:56] == 8'b11011111;
  assign _2098_ = state_in[63:56] == 8'b11011110;
  assign _2099_ = state_in[63:56] == 8'b11011101;
  assign _2100_ = state_in[63:56] == 8'b11011100;
  assign _2101_ = state_in[63:56] == 8'b11011011;
  assign _2102_ = state_in[63:56] == 8'b11011010;
  assign _2103_ = state_in[63:56] == 8'b11011001;
  assign _2104_ = state_in[63:56] == 8'b11011000;
  assign _2105_ = state_in[63:56] == 8'b11010111;
  assign _2106_ = state_in[63:56] == 8'b11010110;
  assign _2107_ = state_in[63:56] == 8'b11010101;
  assign _2108_ = state_in[63:56] == 8'b11010100;
  assign _2109_ = state_in[63:56] == 8'b11010011;
  assign _2110_ = state_in[63:56] == 8'b11010010;
  assign _2111_ = state_in[63:56] == 8'b11010001;
  assign _2112_ = state_in[63:56] == 8'b11010000;
  assign _2113_ = state_in[63:56] == 8'b11001111;
  assign _2114_ = state_in[63:56] == 8'b11001110;
  assign _2115_ = state_in[63:56] == 8'b11001101;
  assign _2116_ = state_in[63:56] == 8'b11001100;
  assign _2117_ = state_in[63:56] == 8'b11001011;
  assign _2118_ = state_in[63:56] == 8'b11001010;
  assign _2119_ = state_in[63:56] == 8'b11001001;
  assign _2120_ = state_in[63:56] == 8'b11001000;
  assign _2121_ = state_in[63:56] == 8'b11000111;
  assign _2122_ = state_in[63:56] == 8'b11000110;
  assign _2123_ = state_in[63:56] == 8'b11000101;
  assign _2124_ = state_in[63:56] == 8'b11000100;
  assign _2125_ = state_in[63:56] == 8'b11000011;
  assign _2126_ = state_in[63:56] == 8'b11000010;
  assign _2127_ = state_in[63:56] == 8'b11000001;
  assign _2128_ = state_in[63:56] == 8'b11000000;
  assign _2129_ = state_in[63:56] == 8'b10111111;
  assign _2130_ = state_in[63:56] == 8'b10111110;
  assign _2131_ = state_in[63:56] == 8'b10111101;
  assign _2132_ = state_in[63:56] == 8'b10111100;
  assign _2133_ = state_in[63:56] == 8'b10111011;
  assign _2134_ = state_in[63:56] == 8'b10111010;
  assign _2135_ = state_in[63:56] == 8'b10111001;
  assign _2136_ = state_in[63:56] == 8'b10111000;
  assign _2137_ = state_in[63:56] == 8'b10110111;
  assign _2138_ = state_in[63:56] == 8'b10110110;
  assign _2139_ = state_in[63:56] == 8'b10110101;
  assign _2140_ = state_in[63:56] == 8'b10110100;
  assign _2141_ = state_in[63:56] == 8'b10110011;
  assign _2142_ = state_in[63:56] == 8'b10110010;
  assign _2143_ = state_in[63:56] == 8'b10110001;
  assign _2144_ = state_in[63:56] == 8'b10110000;
  assign _2145_ = state_in[63:56] == 8'b10101111;
  assign _2146_ = state_in[63:56] == 8'b10101110;
  assign _2147_ = state_in[63:56] == 8'b10101101;
  assign _2148_ = state_in[63:56] == 8'b10101100;
  assign _2149_ = state_in[63:56] == 8'b10101011;
  assign _2150_ = state_in[63:56] == 8'b10101010;
  assign _2151_ = state_in[63:56] == 8'b10101001;
  assign _2152_ = state_in[63:56] == 8'b10101000;
  assign _2153_ = state_in[63:56] == 8'b10100111;
  assign _2154_ = state_in[63:56] == 8'b10100110;
  assign _2155_ = state_in[63:56] == 8'b10100101;
  assign _2156_ = state_in[63:56] == 8'b10100100;
  assign _2157_ = state_in[63:56] == 8'b10100011;
  assign _2158_ = state_in[63:56] == 8'b10100010;
  assign _2159_ = state_in[63:56] == 8'b10100001;
  assign _2160_ = state_in[63:56] == 8'b10100000;
  assign _2161_ = state_in[63:56] == 8'b10011111;
  assign _2162_ = state_in[63:56] == 8'b10011110;
  assign _2163_ = state_in[63:56] == 8'b10011101;
  assign _2164_ = state_in[63:56] == 8'b10011100;
  assign _2165_ = state_in[63:56] == 8'b10011011;
  assign _2166_ = state_in[63:56] == 8'b10011010;
  assign _2167_ = state_in[63:56] == 8'b10011001;
  assign _2168_ = state_in[63:56] == 8'b10011000;
  assign _2169_ = state_in[63:56] == 8'b10010111;
  assign _2170_ = state_in[63:56] == 8'b10010110;
  assign _2171_ = state_in[63:56] == 8'b10010101;
  assign _2172_ = state_in[63:56] == 8'b10010100;
  assign _2173_ = state_in[63:56] == 8'b10010011;
  assign _2174_ = state_in[63:56] == 8'b10010010;
  assign _2175_ = state_in[63:56] == 8'b10010001;
  assign _2176_ = state_in[63:56] == 8'b10010000;
  assign _2177_ = state_in[63:56] == 8'b10001111;
  assign _2178_ = state_in[63:56] == 8'b10001110;
  assign _2179_ = state_in[63:56] == 8'b10001101;
  assign _2180_ = state_in[63:56] == 8'b10001100;
  assign _2181_ = state_in[63:56] == 8'b10001011;
  assign _2182_ = state_in[63:56] == 8'b10001010;
  assign _2183_ = state_in[63:56] == 8'b10001001;
  assign _2184_ = state_in[63:56] == 8'b10001000;
  assign _2185_ = state_in[63:56] == 8'b10000111;
  assign _2186_ = state_in[63:56] == 8'b10000110;
  assign _2187_ = state_in[63:56] == 8'b10000101;
  assign _2188_ = state_in[63:56] == 8'b10000100;
  assign _2189_ = state_in[63:56] == 8'b10000011;
  assign _2190_ = state_in[63:56] == 8'b10000010;
  assign _2191_ = state_in[63:56] == 8'b10000001;
  assign _2192_ = state_in[63:56] == 8'b10000000;
  assign _2193_ = state_in[63:56] == 7'b1111111;
  assign _2194_ = state_in[63:56] == 7'b1111110;
  assign _2195_ = state_in[63:56] == 7'b1111101;
  assign _2196_ = state_in[63:56] == 7'b1111100;
  assign _2197_ = state_in[63:56] == 7'b1111011;
  assign _2198_ = state_in[63:56] == 7'b1111010;
  assign _2199_ = state_in[63:56] == 7'b1111001;
  assign _2200_ = state_in[63:56] == 7'b1111000;
  assign _2201_ = state_in[63:56] == 7'b1110111;
  assign _2202_ = state_in[63:56] == 7'b1110110;
  assign _2203_ = state_in[63:56] == 7'b1110101;
  assign _2204_ = state_in[63:56] == 7'b1110100;
  assign _2205_ = state_in[63:56] == 7'b1110011;
  assign _2206_ = state_in[63:56] == 7'b1110010;
  assign _2207_ = state_in[63:56] == 7'b1110001;
  assign _2208_ = state_in[63:56] == 7'b1110000;
  assign _2209_ = state_in[63:56] == 7'b1101111;
  assign _2210_ = state_in[63:56] == 7'b1101110;
  assign _2211_ = state_in[63:56] == 7'b1101101;
  assign _2212_ = state_in[63:56] == 7'b1101100;
  assign _2213_ = state_in[63:56] == 7'b1101011;
  assign _2214_ = state_in[63:56] == 7'b1101010;
  assign _2215_ = state_in[63:56] == 7'b1101001;
  assign _2216_ = state_in[63:56] == 7'b1101000;
  assign _2217_ = state_in[63:56] == 7'b1100111;
  assign _2218_ = state_in[63:56] == 7'b1100110;
  assign _2219_ = state_in[63:56] == 7'b1100101;
  assign _2220_ = state_in[63:56] == 7'b1100100;
  assign _2221_ = state_in[63:56] == 7'b1100011;
  assign _2222_ = state_in[63:56] == 7'b1100010;
  assign _2223_ = state_in[63:56] == 7'b1100001;
  assign _2224_ = state_in[63:56] == 7'b1100000;
  assign _2225_ = state_in[63:56] == 7'b1011111;
  assign _2226_ = state_in[63:56] == 7'b1011110;
  assign _2227_ = state_in[63:56] == 7'b1011101;
  assign _2228_ = state_in[63:56] == 7'b1011100;
  assign _2229_ = state_in[63:56] == 7'b1011011;
  assign _2230_ = state_in[63:56] == 7'b1011010;
  assign _2231_ = state_in[63:56] == 7'b1011001;
  assign _2232_ = state_in[63:56] == 7'b1011000;
  assign _2233_ = state_in[63:56] == 7'b1010111;
  assign _2234_ = state_in[63:56] == 7'b1010110;
  assign _2235_ = state_in[63:56] == 7'b1010101;
  assign _2236_ = state_in[63:56] == 7'b1010100;
  assign _2237_ = state_in[63:56] == 7'b1010011;
  assign _2238_ = state_in[63:56] == 7'b1010010;
  assign _2239_ = state_in[63:56] == 7'b1010001;
  assign _2240_ = state_in[63:56] == 7'b1010000;
  assign _2241_ = state_in[63:56] == 7'b1001111;
  assign _2242_ = state_in[63:56] == 7'b1001110;
  assign _2243_ = state_in[63:56] == 7'b1001101;
  assign _2244_ = state_in[63:56] == 7'b1001100;
  assign _2245_ = state_in[63:56] == 7'b1001011;
  assign _2246_ = state_in[63:56] == 7'b1001010;
  assign _2247_ = state_in[63:56] == 7'b1001001;
  assign _2248_ = state_in[63:56] == 7'b1001000;
  assign _2249_ = state_in[63:56] == 7'b1000111;
  assign _2250_ = state_in[63:56] == 7'b1000110;
  assign _2251_ = state_in[63:56] == 7'b1000101;
  assign _2252_ = state_in[63:56] == 7'b1000100;
  assign _2253_ = state_in[63:56] == 7'b1000011;
  assign _2254_ = state_in[63:56] == 7'b1000010;
  assign _2255_ = state_in[63:56] == 7'b1000001;
  assign _2256_ = state_in[63:56] == 7'b1000000;
  assign _2257_ = state_in[63:56] == 6'b111111;
  assign _2258_ = state_in[63:56] == 6'b111110;
  assign _2259_ = state_in[63:56] == 6'b111101;
  assign _2260_ = state_in[63:56] == 6'b111100;
  assign _2261_ = state_in[63:56] == 6'b111011;
  assign _2262_ = state_in[63:56] == 6'b111010;
  assign _2263_ = state_in[63:56] == 6'b111001;
  assign _2264_ = state_in[63:56] == 6'b111000;
  assign _2265_ = state_in[63:56] == 6'b110111;
  assign _2266_ = state_in[63:56] == 6'b110110;
  assign _2267_ = state_in[63:56] == 6'b110101;
  assign _2268_ = state_in[63:56] == 6'b110100;
  assign _2269_ = state_in[63:56] == 6'b110011;
  assign _2270_ = state_in[63:56] == 6'b110010;
  assign _2271_ = state_in[63:56] == 6'b110001;
  assign _2272_ = state_in[63:56] == 6'b110000;
  assign _2273_ = state_in[63:56] == 6'b101111;
  assign _2274_ = state_in[63:56] == 6'b101110;
  assign _2275_ = state_in[63:56] == 6'b101101;
  assign _2276_ = state_in[63:56] == 6'b101100;
  assign _2277_ = state_in[63:56] == 6'b101011;
  assign _2278_ = state_in[63:56] == 6'b101010;
  assign _2279_ = state_in[63:56] == 6'b101001;
  assign _2280_ = state_in[63:56] == 6'b101000;
  assign _2281_ = state_in[63:56] == 6'b100111;
  assign _2282_ = state_in[63:56] == 6'b100110;
  assign _2283_ = state_in[63:56] == 6'b100101;
  assign _2284_ = state_in[63:56] == 6'b100100;
  assign _2285_ = state_in[63:56] == 6'b100011;
  assign _2286_ = state_in[63:56] == 6'b100010;
  assign _2287_ = state_in[63:56] == 6'b100001;
  assign _2288_ = state_in[63:56] == 6'b100000;
  assign _2289_ = state_in[63:56] == 5'b11111;
  assign _2290_ = state_in[63:56] == 5'b11110;
  assign _2291_ = state_in[63:56] == 5'b11101;
  assign _2292_ = state_in[63:56] == 5'b11100;
  assign _2293_ = state_in[63:56] == 5'b11011;
  assign _2294_ = state_in[63:56] == 5'b11010;
  assign _2295_ = state_in[63:56] == 5'b11001;
  assign _2296_ = state_in[63:56] == 5'b11000;
  assign _2297_ = state_in[63:56] == 5'b10111;
  assign _2298_ = state_in[63:56] == 5'b10110;
  assign _2299_ = state_in[63:56] == 5'b10101;
  assign _2300_ = state_in[63:56] == 5'b10100;
  assign _2301_ = state_in[63:56] == 5'b10011;
  assign _2302_ = state_in[63:56] == 5'b10010;
  assign _2303_ = state_in[63:56] == 5'b10001;
  assign _2304_ = state_in[63:56] == 5'b10000;
  assign _2305_ = state_in[63:56] == 4'b1111;
  assign _2306_ = state_in[63:56] == 4'b1110;
  assign _2307_ = state_in[63:56] == 4'b1101;
  assign _2308_ = state_in[63:56] == 4'b1100;
  assign _2309_ = state_in[63:56] == 4'b1011;
  assign _2310_ = state_in[63:56] == 4'b1010;
  assign _2311_ = state_in[63:56] == 4'b1001;
  assign _2312_ = state_in[63:56] == 4'b1000;
  assign _2313_ = state_in[63:56] == 3'b111;
  assign _2314_ = state_in[63:56] == 3'b110;
  assign _2315_ = state_in[63:56] == 3'b101;
  assign _2316_ = state_in[63:56] == 3'b100;
  assign _2317_ = state_in[63:56] == 2'b11;
  assign _2318_ = state_in[63:56] == 2'b10;
  assign _2319_ = state_in[63:56] == 1'b1;
  assign _2320_ = ! state_in[63:56];
  always @(posedge clk)
      \t2.t0.s4.out <= _2321_;
  logic [255:0] fangyuan18;
  assign fangyuan18 = { _2320_, _2319_, _2318_, _2317_, _2316_, _2315_, _2314_, _2313_, _2312_, _2311_, _2310_, _2309_, _2308_, _2307_, _2306_, _2305_, _2304_, _2303_, _2302_, _2301_, _2300_, _2299_, _2298_, _2297_, _2296_, _2295_, _2294_, _2293_, _2292_, _2291_, _2290_, _2289_, _2288_, _2287_, _2286_, _2285_, _2284_, _2283_, _2282_, _2281_, _2280_, _2279_, _2278_, _2277_, _2276_, _2275_, _2274_, _2273_, _2272_, _2271_, _2270_, _2269_, _2268_, _2267_, _2266_, _2265_, _2264_, _2263_, _2262_, _2261_, _2260_, _2259_, _2258_, _2257_, _2256_, _2255_, _2254_, _2253_, _2252_, _2251_, _2250_, _2249_, _2248_, _2247_, _2246_, _2245_, _2244_, _2243_, _2242_, _2241_, _2240_, _2239_, _2238_, _2237_, _2236_, _2235_, _2234_, _2233_, _2232_, _2231_, _2230_, _2229_, _2228_, _2227_, _2226_, _2225_, _2224_, _2223_, _2222_, _2221_, _2220_, _2219_, _2218_, _2217_, _2216_, _2215_, _2214_, _2213_, _2212_, _2211_, _2210_, _2209_, _2208_, _2207_, _2206_, _2205_, _2204_, _2203_, _2202_, _2201_, _2200_, _2199_, _2198_, _2197_, _2196_, _2195_, _2194_, _2193_, _2192_, _2191_, _2190_, _2189_, _2188_, _2187_, _2186_, _2185_, _2184_, _2183_, _2182_, _2181_, _2180_, _2179_, _2178_, _2177_, _2176_, _2175_, _2174_, _2173_, _2172_, _2171_, _2170_, _2169_, _2168_, _2167_, _2166_, _2165_, _2164_, _2163_, _2162_, _2161_, _2160_, _2159_, _2158_, _2157_, _2156_, _2155_, _2154_, _2153_, _2152_, _2151_, _2150_, _2149_, _2148_, _2147_, _2146_, _2145_, _2144_, _2143_, _2142_, _2141_, _2140_, _2139_, _2138_, _2137_, _2136_, _2135_, _2134_, _2133_, _2132_, _2131_, _2130_, _2129_, _2128_, _2127_, _2126_, _2125_, _2124_, _2123_, _2122_, _2121_, _2120_, _2119_, _2118_, _2117_, _2116_, _2115_, _2114_, _2113_, _2112_, _2111_, _2110_, _2109_, _2108_, _2107_, _2106_, _2105_, _2104_, _2103_, _2102_, _2101_, _2100_, _2099_, _2098_, _2097_, _2096_, _2095_, _2094_, _2093_, _2092_, _2091_, _2090_, _2089_, _2088_, _2087_, _2086_, _2085_, _2084_, _2083_, _2082_, _2081_, _2080_, _2079_, _2078_, _2077_, _2076_, _2075_, _2074_, _2073_, _2072_, _2071_, _2070_, _2069_, _2068_, _2067_, _2066_, _2065_ };

  always @(\t2.t0.s4.out or fangyuan18) begin
    casez (fangyuan18)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2321_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2321_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2321_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2321_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2321_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2321_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2321_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2321_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2321_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2321_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2321_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2321_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2321_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2321_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2321_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2321_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2321_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2321_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2321_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2321_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2321_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2321_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2321_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2321_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2321_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2321_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2321_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2321_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2321_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2321_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2321_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2321_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2321_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2321_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2321_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2321_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2321_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2321_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2321_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2321_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2321_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2321_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2321_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2321_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2321_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2321_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2321_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2321_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2321_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2321_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2321_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2321_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2321_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2321_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2321_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2321_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2321_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2321_ = 8'b11000110 ;
      default:
        _2321_ = \t2.t0.s4.out ;
    endcase
  end
  assign p21[31:24] = \t2.t1.s0.out ^ \t2.t1.s4.out ;
  always @(posedge clk)
      \t2.t1.s0.out <= _2322_;
  logic [255:0] fangyuan19;
  assign fangyuan19 = { _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _2524_, _2523_, _2522_, _2521_, _2520_, _2519_, _2518_, _2517_, _2516_, _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_, _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_ };

  always @(\t2.t1.s0.out or fangyuan19) begin
    casez (fangyuan19)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2322_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2322_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2322_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2322_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2322_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2322_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2322_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2322_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2322_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2322_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2322_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2322_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2322_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2322_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2322_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2322_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2322_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2322_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2322_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2322_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2322_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2322_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2322_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2322_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2322_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2322_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2322_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2322_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2322_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2322_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2322_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2322_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2322_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2322_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2322_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2322_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2322_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2322_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2322_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2322_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2322_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2322_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2322_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2322_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2322_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2322_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2322_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2322_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2322_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2322_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2322_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2322_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2322_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2322_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2322_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2322_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2322_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2322_ = 8'b01100011 ;
      default:
        _2322_ = \t2.t1.s0.out ;
    endcase
  end
  assign _2323_ = state_in[55:48] == 8'b11111111;
  assign _2324_ = state_in[55:48] == 8'b11111110;
  assign _2325_ = state_in[55:48] == 8'b11111101;
  assign _2326_ = state_in[55:48] == 8'b11111100;
  assign _2327_ = state_in[55:48] == 8'b11111011;
  assign _2328_ = state_in[55:48] == 8'b11111010;
  assign _2329_ = state_in[55:48] == 8'b11111001;
  assign _2330_ = state_in[55:48] == 8'b11111000;
  assign _2331_ = state_in[55:48] == 8'b11110111;
  assign _2332_ = state_in[55:48] == 8'b11110110;
  assign _2333_ = state_in[55:48] == 8'b11110101;
  assign _2334_ = state_in[55:48] == 8'b11110100;
  assign _2335_ = state_in[55:48] == 8'b11110011;
  assign _2336_ = state_in[55:48] == 8'b11110010;
  assign _2337_ = state_in[55:48] == 8'b11110001;
  assign _2338_ = state_in[55:48] == 8'b11110000;
  assign _2339_ = state_in[55:48] == 8'b11101111;
  assign _2340_ = state_in[55:48] == 8'b11101110;
  assign _2341_ = state_in[55:48] == 8'b11101101;
  assign _2342_ = state_in[55:48] == 8'b11101100;
  assign _2343_ = state_in[55:48] == 8'b11101011;
  assign _2344_ = state_in[55:48] == 8'b11101010;
  assign _2345_ = state_in[55:48] == 8'b11101001;
  assign _2346_ = state_in[55:48] == 8'b11101000;
  assign _2347_ = state_in[55:48] == 8'b11100111;
  assign _2348_ = state_in[55:48] == 8'b11100110;
  assign _2349_ = state_in[55:48] == 8'b11100101;
  assign _2350_ = state_in[55:48] == 8'b11100100;
  assign _2351_ = state_in[55:48] == 8'b11100011;
  assign _2352_ = state_in[55:48] == 8'b11100010;
  assign _2353_ = state_in[55:48] == 8'b11100001;
  assign _2354_ = state_in[55:48] == 8'b11100000;
  assign _2355_ = state_in[55:48] == 8'b11011111;
  assign _2356_ = state_in[55:48] == 8'b11011110;
  assign _2357_ = state_in[55:48] == 8'b11011101;
  assign _2358_ = state_in[55:48] == 8'b11011100;
  assign _2359_ = state_in[55:48] == 8'b11011011;
  assign _2360_ = state_in[55:48] == 8'b11011010;
  assign _2361_ = state_in[55:48] == 8'b11011001;
  assign _2362_ = state_in[55:48] == 8'b11011000;
  assign _2363_ = state_in[55:48] == 8'b11010111;
  assign _2364_ = state_in[55:48] == 8'b11010110;
  assign _2365_ = state_in[55:48] == 8'b11010101;
  assign _2366_ = state_in[55:48] == 8'b11010100;
  assign _2367_ = state_in[55:48] == 8'b11010011;
  assign _2368_ = state_in[55:48] == 8'b11010010;
  assign _2369_ = state_in[55:48] == 8'b11010001;
  assign _2370_ = state_in[55:48] == 8'b11010000;
  assign _2371_ = state_in[55:48] == 8'b11001111;
  assign _2372_ = state_in[55:48] == 8'b11001110;
  assign _2373_ = state_in[55:48] == 8'b11001101;
  assign _2374_ = state_in[55:48] == 8'b11001100;
  assign _2375_ = state_in[55:48] == 8'b11001011;
  assign _2376_ = state_in[55:48] == 8'b11001010;
  assign _2377_ = state_in[55:48] == 8'b11001001;
  assign _2378_ = state_in[55:48] == 8'b11001000;
  assign _2379_ = state_in[55:48] == 8'b11000111;
  assign _2380_ = state_in[55:48] == 8'b11000110;
  assign _2381_ = state_in[55:48] == 8'b11000101;
  assign _2382_ = state_in[55:48] == 8'b11000100;
  assign _2383_ = state_in[55:48] == 8'b11000011;
  assign _2384_ = state_in[55:48] == 8'b11000010;
  assign _2385_ = state_in[55:48] == 8'b11000001;
  assign _2386_ = state_in[55:48] == 8'b11000000;
  assign _2387_ = state_in[55:48] == 8'b10111111;
  assign _2388_ = state_in[55:48] == 8'b10111110;
  assign _2389_ = state_in[55:48] == 8'b10111101;
  assign _2390_ = state_in[55:48] == 8'b10111100;
  assign _2391_ = state_in[55:48] == 8'b10111011;
  assign _2392_ = state_in[55:48] == 8'b10111010;
  assign _2393_ = state_in[55:48] == 8'b10111001;
  assign _2394_ = state_in[55:48] == 8'b10111000;
  assign _2395_ = state_in[55:48] == 8'b10110111;
  assign _2396_ = state_in[55:48] == 8'b10110110;
  assign _2397_ = state_in[55:48] == 8'b10110101;
  assign _2398_ = state_in[55:48] == 8'b10110100;
  assign _2399_ = state_in[55:48] == 8'b10110011;
  assign _2400_ = state_in[55:48] == 8'b10110010;
  assign _2401_ = state_in[55:48] == 8'b10110001;
  assign _2402_ = state_in[55:48] == 8'b10110000;
  assign _2403_ = state_in[55:48] == 8'b10101111;
  assign _2404_ = state_in[55:48] == 8'b10101110;
  assign _2405_ = state_in[55:48] == 8'b10101101;
  assign _2406_ = state_in[55:48] == 8'b10101100;
  assign _2407_ = state_in[55:48] == 8'b10101011;
  assign _2408_ = state_in[55:48] == 8'b10101010;
  assign _2409_ = state_in[55:48] == 8'b10101001;
  assign _2410_ = state_in[55:48] == 8'b10101000;
  assign _2411_ = state_in[55:48] == 8'b10100111;
  assign _2412_ = state_in[55:48] == 8'b10100110;
  assign _2413_ = state_in[55:48] == 8'b10100101;
  assign _2414_ = state_in[55:48] == 8'b10100100;
  assign _2415_ = state_in[55:48] == 8'b10100011;
  assign _2416_ = state_in[55:48] == 8'b10100010;
  assign _2417_ = state_in[55:48] == 8'b10100001;
  assign _2418_ = state_in[55:48] == 8'b10100000;
  assign _2419_ = state_in[55:48] == 8'b10011111;
  assign _2420_ = state_in[55:48] == 8'b10011110;
  assign _2421_ = state_in[55:48] == 8'b10011101;
  assign _2422_ = state_in[55:48] == 8'b10011100;
  assign _2423_ = state_in[55:48] == 8'b10011011;
  assign _2424_ = state_in[55:48] == 8'b10011010;
  assign _2425_ = state_in[55:48] == 8'b10011001;
  assign _2426_ = state_in[55:48] == 8'b10011000;
  assign _2427_ = state_in[55:48] == 8'b10010111;
  assign _2428_ = state_in[55:48] == 8'b10010110;
  assign _2429_ = state_in[55:48] == 8'b10010101;
  assign _2430_ = state_in[55:48] == 8'b10010100;
  assign _2431_ = state_in[55:48] == 8'b10010011;
  assign _2432_ = state_in[55:48] == 8'b10010010;
  assign _2433_ = state_in[55:48] == 8'b10010001;
  assign _2434_ = state_in[55:48] == 8'b10010000;
  assign _2435_ = state_in[55:48] == 8'b10001111;
  assign _2436_ = state_in[55:48] == 8'b10001110;
  assign _2437_ = state_in[55:48] == 8'b10001101;
  assign _2438_ = state_in[55:48] == 8'b10001100;
  assign _2439_ = state_in[55:48] == 8'b10001011;
  assign _2440_ = state_in[55:48] == 8'b10001010;
  assign _2441_ = state_in[55:48] == 8'b10001001;
  assign _2442_ = state_in[55:48] == 8'b10001000;
  assign _2443_ = state_in[55:48] == 8'b10000111;
  assign _2444_ = state_in[55:48] == 8'b10000110;
  assign _2445_ = state_in[55:48] == 8'b10000101;
  assign _2446_ = state_in[55:48] == 8'b10000100;
  assign _2447_ = state_in[55:48] == 8'b10000011;
  assign _2448_ = state_in[55:48] == 8'b10000010;
  assign _2449_ = state_in[55:48] == 8'b10000001;
  assign _2450_ = state_in[55:48] == 8'b10000000;
  assign _2451_ = state_in[55:48] == 7'b1111111;
  assign _2452_ = state_in[55:48] == 7'b1111110;
  assign _2453_ = state_in[55:48] == 7'b1111101;
  assign _2454_ = state_in[55:48] == 7'b1111100;
  assign _2455_ = state_in[55:48] == 7'b1111011;
  assign _2456_ = state_in[55:48] == 7'b1111010;
  assign _2457_ = state_in[55:48] == 7'b1111001;
  assign _2458_ = state_in[55:48] == 7'b1111000;
  assign _2459_ = state_in[55:48] == 7'b1110111;
  assign _2460_ = state_in[55:48] == 7'b1110110;
  assign _2461_ = state_in[55:48] == 7'b1110101;
  assign _2462_ = state_in[55:48] == 7'b1110100;
  assign _2463_ = state_in[55:48] == 7'b1110011;
  assign _2464_ = state_in[55:48] == 7'b1110010;
  assign _2465_ = state_in[55:48] == 7'b1110001;
  assign _2466_ = state_in[55:48] == 7'b1110000;
  assign _2467_ = state_in[55:48] == 7'b1101111;
  assign _2468_ = state_in[55:48] == 7'b1101110;
  assign _2469_ = state_in[55:48] == 7'b1101101;
  assign _2470_ = state_in[55:48] == 7'b1101100;
  assign _2471_ = state_in[55:48] == 7'b1101011;
  assign _2472_ = state_in[55:48] == 7'b1101010;
  assign _2473_ = state_in[55:48] == 7'b1101001;
  assign _2474_ = state_in[55:48] == 7'b1101000;
  assign _2475_ = state_in[55:48] == 7'b1100111;
  assign _2476_ = state_in[55:48] == 7'b1100110;
  assign _2477_ = state_in[55:48] == 7'b1100101;
  assign _2478_ = state_in[55:48] == 7'b1100100;
  assign _2479_ = state_in[55:48] == 7'b1100011;
  assign _2480_ = state_in[55:48] == 7'b1100010;
  assign _2481_ = state_in[55:48] == 7'b1100001;
  assign _2482_ = state_in[55:48] == 7'b1100000;
  assign _2483_ = state_in[55:48] == 7'b1011111;
  assign _2484_ = state_in[55:48] == 7'b1011110;
  assign _2485_ = state_in[55:48] == 7'b1011101;
  assign _2486_ = state_in[55:48] == 7'b1011100;
  assign _2487_ = state_in[55:48] == 7'b1011011;
  assign _2488_ = state_in[55:48] == 7'b1011010;
  assign _2489_ = state_in[55:48] == 7'b1011001;
  assign _2490_ = state_in[55:48] == 7'b1011000;
  assign _2491_ = state_in[55:48] == 7'b1010111;
  assign _2492_ = state_in[55:48] == 7'b1010110;
  assign _2493_ = state_in[55:48] == 7'b1010101;
  assign _2494_ = state_in[55:48] == 7'b1010100;
  assign _2495_ = state_in[55:48] == 7'b1010011;
  assign _2496_ = state_in[55:48] == 7'b1010010;
  assign _2497_ = state_in[55:48] == 7'b1010001;
  assign _2498_ = state_in[55:48] == 7'b1010000;
  assign _2499_ = state_in[55:48] == 7'b1001111;
  assign _2500_ = state_in[55:48] == 7'b1001110;
  assign _2501_ = state_in[55:48] == 7'b1001101;
  assign _2502_ = state_in[55:48] == 7'b1001100;
  assign _2503_ = state_in[55:48] == 7'b1001011;
  assign _2504_ = state_in[55:48] == 7'b1001010;
  assign _2505_ = state_in[55:48] == 7'b1001001;
  assign _2506_ = state_in[55:48] == 7'b1001000;
  assign _2507_ = state_in[55:48] == 7'b1000111;
  assign _2508_ = state_in[55:48] == 7'b1000110;
  assign _2509_ = state_in[55:48] == 7'b1000101;
  assign _2510_ = state_in[55:48] == 7'b1000100;
  assign _2511_ = state_in[55:48] == 7'b1000011;
  assign _2512_ = state_in[55:48] == 7'b1000010;
  assign _2513_ = state_in[55:48] == 7'b1000001;
  assign _2514_ = state_in[55:48] == 7'b1000000;
  assign _2515_ = state_in[55:48] == 6'b111111;
  assign _2516_ = state_in[55:48] == 6'b111110;
  assign _2517_ = state_in[55:48] == 6'b111101;
  assign _2518_ = state_in[55:48] == 6'b111100;
  assign _2519_ = state_in[55:48] == 6'b111011;
  assign _2520_ = state_in[55:48] == 6'b111010;
  assign _2521_ = state_in[55:48] == 6'b111001;
  assign _2522_ = state_in[55:48] == 6'b111000;
  assign _2523_ = state_in[55:48] == 6'b110111;
  assign _2524_ = state_in[55:48] == 6'b110110;
  assign _2525_ = state_in[55:48] == 6'b110101;
  assign _2526_ = state_in[55:48] == 6'b110100;
  assign _2527_ = state_in[55:48] == 6'b110011;
  assign _2528_ = state_in[55:48] == 6'b110010;
  assign _2529_ = state_in[55:48] == 6'b110001;
  assign _2530_ = state_in[55:48] == 6'b110000;
  assign _2531_ = state_in[55:48] == 6'b101111;
  assign _2532_ = state_in[55:48] == 6'b101110;
  assign _2533_ = state_in[55:48] == 6'b101101;
  assign _2534_ = state_in[55:48] == 6'b101100;
  assign _2535_ = state_in[55:48] == 6'b101011;
  assign _2536_ = state_in[55:48] == 6'b101010;
  assign _2537_ = state_in[55:48] == 6'b101001;
  assign _2538_ = state_in[55:48] == 6'b101000;
  assign _2539_ = state_in[55:48] == 6'b100111;
  assign _2540_ = state_in[55:48] == 6'b100110;
  assign _2541_ = state_in[55:48] == 6'b100101;
  assign _2542_ = state_in[55:48] == 6'b100100;
  assign _2543_ = state_in[55:48] == 6'b100011;
  assign _2544_ = state_in[55:48] == 6'b100010;
  assign _2545_ = state_in[55:48] == 6'b100001;
  assign _2546_ = state_in[55:48] == 6'b100000;
  assign _2547_ = state_in[55:48] == 5'b11111;
  assign _2548_ = state_in[55:48] == 5'b11110;
  assign _2549_ = state_in[55:48] == 5'b11101;
  assign _2550_ = state_in[55:48] == 5'b11100;
  assign _2551_ = state_in[55:48] == 5'b11011;
  assign _2552_ = state_in[55:48] == 5'b11010;
  assign _2553_ = state_in[55:48] == 5'b11001;
  assign _2554_ = state_in[55:48] == 5'b11000;
  assign _2555_ = state_in[55:48] == 5'b10111;
  assign _2556_ = state_in[55:48] == 5'b10110;
  assign _2557_ = state_in[55:48] == 5'b10101;
  assign _2558_ = state_in[55:48] == 5'b10100;
  assign _2559_ = state_in[55:48] == 5'b10011;
  assign _2560_ = state_in[55:48] == 5'b10010;
  assign _2561_ = state_in[55:48] == 5'b10001;
  assign _2562_ = state_in[55:48] == 5'b10000;
  assign _2563_ = state_in[55:48] == 4'b1111;
  assign _2564_ = state_in[55:48] == 4'b1110;
  assign _2565_ = state_in[55:48] == 4'b1101;
  assign _2566_ = state_in[55:48] == 4'b1100;
  assign _2567_ = state_in[55:48] == 4'b1011;
  assign _2568_ = state_in[55:48] == 4'b1010;
  assign _2569_ = state_in[55:48] == 4'b1001;
  assign _2570_ = state_in[55:48] == 4'b1000;
  assign _2571_ = state_in[55:48] == 3'b111;
  assign _2572_ = state_in[55:48] == 3'b110;
  assign _2573_ = state_in[55:48] == 3'b101;
  assign _2574_ = state_in[55:48] == 3'b100;
  assign _2575_ = state_in[55:48] == 2'b11;
  assign _2576_ = state_in[55:48] == 2'b10;
  assign _2577_ = state_in[55:48] == 1'b1;
  assign _2578_ = ! state_in[55:48];
  always @(posedge clk)
      \t2.t1.s4.out <= _2579_;
  logic [255:0] fangyuan20;
  assign fangyuan20 = { _2578_, _2577_, _2576_, _2575_, _2574_, _2573_, _2572_, _2571_, _2570_, _2569_, _2568_, _2567_, _2566_, _2565_, _2564_, _2563_, _2562_, _2561_, _2560_, _2559_, _2558_, _2557_, _2556_, _2555_, _2554_, _2553_, _2552_, _2551_, _2550_, _2549_, _2548_, _2547_, _2546_, _2545_, _2544_, _2543_, _2542_, _2541_, _2540_, _2539_, _2538_, _2537_, _2536_, _2535_, _2534_, _2533_, _2532_, _2531_, _2530_, _2529_, _2528_, _2527_, _2526_, _2525_, _2524_, _2523_, _2522_, _2521_, _2520_, _2519_, _2518_, _2517_, _2516_, _2515_, _2514_, _2513_, _2512_, _2511_, _2510_, _2509_, _2508_, _2507_, _2506_, _2505_, _2504_, _2503_, _2502_, _2501_, _2500_, _2499_, _2498_, _2497_, _2496_, _2495_, _2494_, _2493_, _2492_, _2491_, _2490_, _2489_, _2488_, _2487_, _2486_, _2485_, _2484_, _2483_, _2482_, _2481_, _2480_, _2479_, _2478_, _2477_, _2476_, _2475_, _2474_, _2473_, _2472_, _2471_, _2470_, _2469_, _2468_, _2467_, _2466_, _2465_, _2464_, _2463_, _2462_, _2461_, _2460_, _2459_, _2458_, _2457_, _2456_, _2455_, _2454_, _2453_, _2452_, _2451_, _2450_, _2449_, _2448_, _2447_, _2446_, _2445_, _2444_, _2443_, _2442_, _2441_, _2440_, _2439_, _2438_, _2437_, _2436_, _2435_, _2434_, _2433_, _2432_, _2431_, _2430_, _2429_, _2428_, _2427_, _2426_, _2425_, _2424_, _2423_, _2422_, _2421_, _2420_, _2419_, _2418_, _2417_, _2416_, _2415_, _2414_, _2413_, _2412_, _2411_, _2410_, _2409_, _2408_, _2407_, _2406_, _2405_, _2404_, _2403_, _2402_, _2401_, _2400_, _2399_, _2398_, _2397_, _2396_, _2395_, _2394_, _2393_, _2392_, _2391_, _2390_, _2389_, _2388_, _2387_, _2386_, _2385_, _2384_, _2383_, _2382_, _2381_, _2380_, _2379_, _2378_, _2377_, _2376_, _2375_, _2374_, _2373_, _2372_, _2371_, _2370_, _2369_, _2368_, _2367_, _2366_, _2365_, _2364_, _2363_, _2362_, _2361_, _2360_, _2359_, _2358_, _2357_, _2356_, _2355_, _2354_, _2353_, _2352_, _2351_, _2350_, _2349_, _2348_, _2347_, _2346_, _2345_, _2344_, _2343_, _2342_, _2341_, _2340_, _2339_, _2338_, _2337_, _2336_, _2335_, _2334_, _2333_, _2332_, _2331_, _2330_, _2329_, _2328_, _2327_, _2326_, _2325_, _2324_, _2323_ };

  always @(\t2.t1.s4.out or fangyuan20) begin
    casez (fangyuan20)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2579_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2579_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2579_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2579_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2579_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2579_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2579_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2579_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2579_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2579_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2579_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2579_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2579_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2579_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2579_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2579_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2579_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2579_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2579_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2579_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2579_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2579_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2579_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2579_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2579_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2579_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2579_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2579_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2579_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2579_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2579_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2579_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2579_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2579_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2579_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2579_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2579_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2579_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2579_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2579_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2579_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2579_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2579_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2579_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2579_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2579_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2579_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2579_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2579_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2579_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2579_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2579_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2579_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2579_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2579_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2579_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2579_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2579_ = 8'b11000110 ;
      default:
        _2579_ = \t2.t1.s4.out ;
    endcase
  end
  assign p22[23:16] = \t2.t2.s0.out ^ \t2.t2.s4.out ;
  always @(posedge clk)
      \t2.t2.s0.out <= _2580_;
  logic [255:0] fangyuan21;
  assign fangyuan21 = { _2836_, _2835_, _2834_, _2833_, _2832_, _2831_, _2830_, _2829_, _2828_, _2827_, _2826_, _2825_, _2824_, _2823_, _2822_, _2821_, _2820_, _2819_, _2818_, _2817_, _2816_, _2815_, _2814_, _2813_, _2812_, _2811_, _2810_, _2809_, _2808_, _2807_, _2806_, _2805_, _2804_, _2803_, _2802_, _2801_, _2800_, _2799_, _2798_, _2797_, _2796_, _2795_, _2794_, _2793_, _2792_, _2791_, _2790_, _2789_, _2788_, _2787_, _2786_, _2785_, _2784_, _2783_, _2782_, _2781_, _2780_, _2779_, _2778_, _2777_, _2776_, _2775_, _2774_, _2773_, _2772_, _2771_, _2770_, _2769_, _2768_, _2767_, _2766_, _2765_, _2764_, _2763_, _2762_, _2761_, _2760_, _2759_, _2758_, _2757_, _2756_, _2755_, _2754_, _2753_, _2752_, _2751_, _2750_, _2749_, _2748_, _2747_, _2746_, _2745_, _2744_, _2743_, _2742_, _2741_, _2740_, _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_, _2732_, _2731_, _2730_, _2729_, _2728_, _2727_, _2726_, _2725_, _2724_, _2723_, _2722_, _2721_, _2720_, _2719_, _2718_, _2717_, _2716_, _2715_, _2714_, _2713_, _2712_, _2711_, _2710_, _2709_, _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_ };

  always @(\t2.t2.s0.out or fangyuan21) begin
    casez (fangyuan21)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2580_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2580_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2580_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2580_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2580_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2580_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2580_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2580_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2580_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2580_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2580_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2580_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2580_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2580_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2580_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2580_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2580_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2580_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2580_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2580_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2580_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2580_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2580_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2580_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2580_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2580_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2580_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2580_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2580_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2580_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2580_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2580_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2580_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2580_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2580_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2580_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2580_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2580_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2580_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2580_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2580_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2580_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2580_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2580_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2580_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2580_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2580_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2580_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2580_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2580_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2580_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2580_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2580_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2580_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2580_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2580_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2580_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2580_ = 8'b01100011 ;
      default:
        _2580_ = \t2.t2.s0.out ;
    endcase
  end
  assign _2581_ = state_in[47:40] == 8'b11111111;
  assign _2582_ = state_in[47:40] == 8'b11111110;
  assign _2583_ = state_in[47:40] == 8'b11111101;
  assign _2584_ = state_in[47:40] == 8'b11111100;
  assign _2585_ = state_in[47:40] == 8'b11111011;
  assign _2586_ = state_in[47:40] == 8'b11111010;
  assign _2587_ = state_in[47:40] == 8'b11111001;
  assign _2588_ = state_in[47:40] == 8'b11111000;
  assign _2589_ = state_in[47:40] == 8'b11110111;
  assign _2590_ = state_in[47:40] == 8'b11110110;
  assign _2591_ = state_in[47:40] == 8'b11110101;
  assign _2592_ = state_in[47:40] == 8'b11110100;
  assign _2593_ = state_in[47:40] == 8'b11110011;
  assign _2594_ = state_in[47:40] == 8'b11110010;
  assign _2595_ = state_in[47:40] == 8'b11110001;
  assign _2596_ = state_in[47:40] == 8'b11110000;
  assign _2597_ = state_in[47:40] == 8'b11101111;
  assign _2598_ = state_in[47:40] == 8'b11101110;
  assign _2599_ = state_in[47:40] == 8'b11101101;
  assign _2600_ = state_in[47:40] == 8'b11101100;
  assign _2601_ = state_in[47:40] == 8'b11101011;
  assign _2602_ = state_in[47:40] == 8'b11101010;
  assign _2603_ = state_in[47:40] == 8'b11101001;
  assign _2604_ = state_in[47:40] == 8'b11101000;
  assign _2605_ = state_in[47:40] == 8'b11100111;
  assign _2606_ = state_in[47:40] == 8'b11100110;
  assign _2607_ = state_in[47:40] == 8'b11100101;
  assign _2608_ = state_in[47:40] == 8'b11100100;
  assign _2609_ = state_in[47:40] == 8'b11100011;
  assign _2610_ = state_in[47:40] == 8'b11100010;
  assign _2611_ = state_in[47:40] == 8'b11100001;
  assign _2612_ = state_in[47:40] == 8'b11100000;
  assign _2613_ = state_in[47:40] == 8'b11011111;
  assign _2614_ = state_in[47:40] == 8'b11011110;
  assign _2615_ = state_in[47:40] == 8'b11011101;
  assign _2616_ = state_in[47:40] == 8'b11011100;
  assign _2617_ = state_in[47:40] == 8'b11011011;
  assign _2618_ = state_in[47:40] == 8'b11011010;
  assign _2619_ = state_in[47:40] == 8'b11011001;
  assign _2620_ = state_in[47:40] == 8'b11011000;
  assign _2621_ = state_in[47:40] == 8'b11010111;
  assign _2622_ = state_in[47:40] == 8'b11010110;
  assign _2623_ = state_in[47:40] == 8'b11010101;
  assign _2624_ = state_in[47:40] == 8'b11010100;
  assign _2625_ = state_in[47:40] == 8'b11010011;
  assign _2626_ = state_in[47:40] == 8'b11010010;
  assign _2627_ = state_in[47:40] == 8'b11010001;
  assign _2628_ = state_in[47:40] == 8'b11010000;
  assign _2629_ = state_in[47:40] == 8'b11001111;
  assign _2630_ = state_in[47:40] == 8'b11001110;
  assign _2631_ = state_in[47:40] == 8'b11001101;
  assign _2632_ = state_in[47:40] == 8'b11001100;
  assign _2633_ = state_in[47:40] == 8'b11001011;
  assign _2634_ = state_in[47:40] == 8'b11001010;
  assign _2635_ = state_in[47:40] == 8'b11001001;
  assign _2636_ = state_in[47:40] == 8'b11001000;
  assign _2637_ = state_in[47:40] == 8'b11000111;
  assign _2638_ = state_in[47:40] == 8'b11000110;
  assign _2639_ = state_in[47:40] == 8'b11000101;
  assign _2640_ = state_in[47:40] == 8'b11000100;
  assign _2641_ = state_in[47:40] == 8'b11000011;
  assign _2642_ = state_in[47:40] == 8'b11000010;
  assign _2643_ = state_in[47:40] == 8'b11000001;
  assign _2644_ = state_in[47:40] == 8'b11000000;
  assign _2645_ = state_in[47:40] == 8'b10111111;
  assign _2646_ = state_in[47:40] == 8'b10111110;
  assign _2647_ = state_in[47:40] == 8'b10111101;
  assign _2648_ = state_in[47:40] == 8'b10111100;
  assign _2649_ = state_in[47:40] == 8'b10111011;
  assign _2650_ = state_in[47:40] == 8'b10111010;
  assign _2651_ = state_in[47:40] == 8'b10111001;
  assign _2652_ = state_in[47:40] == 8'b10111000;
  assign _2653_ = state_in[47:40] == 8'b10110111;
  assign _2654_ = state_in[47:40] == 8'b10110110;
  assign _2655_ = state_in[47:40] == 8'b10110101;
  assign _2656_ = state_in[47:40] == 8'b10110100;
  assign _2657_ = state_in[47:40] == 8'b10110011;
  assign _2658_ = state_in[47:40] == 8'b10110010;
  assign _2659_ = state_in[47:40] == 8'b10110001;
  assign _2660_ = state_in[47:40] == 8'b10110000;
  assign _2661_ = state_in[47:40] == 8'b10101111;
  assign _2662_ = state_in[47:40] == 8'b10101110;
  assign _2663_ = state_in[47:40] == 8'b10101101;
  assign _2664_ = state_in[47:40] == 8'b10101100;
  assign _2665_ = state_in[47:40] == 8'b10101011;
  assign _2666_ = state_in[47:40] == 8'b10101010;
  assign _2667_ = state_in[47:40] == 8'b10101001;
  assign _2668_ = state_in[47:40] == 8'b10101000;
  assign _2669_ = state_in[47:40] == 8'b10100111;
  assign _2670_ = state_in[47:40] == 8'b10100110;
  assign _2671_ = state_in[47:40] == 8'b10100101;
  assign _2672_ = state_in[47:40] == 8'b10100100;
  assign _2673_ = state_in[47:40] == 8'b10100011;
  assign _2674_ = state_in[47:40] == 8'b10100010;
  assign _2675_ = state_in[47:40] == 8'b10100001;
  assign _2676_ = state_in[47:40] == 8'b10100000;
  assign _2677_ = state_in[47:40] == 8'b10011111;
  assign _2678_ = state_in[47:40] == 8'b10011110;
  assign _2679_ = state_in[47:40] == 8'b10011101;
  assign _2680_ = state_in[47:40] == 8'b10011100;
  assign _2681_ = state_in[47:40] == 8'b10011011;
  assign _2682_ = state_in[47:40] == 8'b10011010;
  assign _2683_ = state_in[47:40] == 8'b10011001;
  assign _2684_ = state_in[47:40] == 8'b10011000;
  assign _2685_ = state_in[47:40] == 8'b10010111;
  assign _2686_ = state_in[47:40] == 8'b10010110;
  assign _2687_ = state_in[47:40] == 8'b10010101;
  assign _2688_ = state_in[47:40] == 8'b10010100;
  assign _2689_ = state_in[47:40] == 8'b10010011;
  assign _2690_ = state_in[47:40] == 8'b10010010;
  assign _2691_ = state_in[47:40] == 8'b10010001;
  assign _2692_ = state_in[47:40] == 8'b10010000;
  assign _2693_ = state_in[47:40] == 8'b10001111;
  assign _2694_ = state_in[47:40] == 8'b10001110;
  assign _2695_ = state_in[47:40] == 8'b10001101;
  assign _2696_ = state_in[47:40] == 8'b10001100;
  assign _2697_ = state_in[47:40] == 8'b10001011;
  assign _2698_ = state_in[47:40] == 8'b10001010;
  assign _2699_ = state_in[47:40] == 8'b10001001;
  assign _2700_ = state_in[47:40] == 8'b10001000;
  assign _2701_ = state_in[47:40] == 8'b10000111;
  assign _2702_ = state_in[47:40] == 8'b10000110;
  assign _2703_ = state_in[47:40] == 8'b10000101;
  assign _2704_ = state_in[47:40] == 8'b10000100;
  assign _2705_ = state_in[47:40] == 8'b10000011;
  assign _2706_ = state_in[47:40] == 8'b10000010;
  assign _2707_ = state_in[47:40] == 8'b10000001;
  assign _2708_ = state_in[47:40] == 8'b10000000;
  assign _2709_ = state_in[47:40] == 7'b1111111;
  assign _2710_ = state_in[47:40] == 7'b1111110;
  assign _2711_ = state_in[47:40] == 7'b1111101;
  assign _2712_ = state_in[47:40] == 7'b1111100;
  assign _2713_ = state_in[47:40] == 7'b1111011;
  assign _2714_ = state_in[47:40] == 7'b1111010;
  assign _2715_ = state_in[47:40] == 7'b1111001;
  assign _2716_ = state_in[47:40] == 7'b1111000;
  assign _2717_ = state_in[47:40] == 7'b1110111;
  assign _2718_ = state_in[47:40] == 7'b1110110;
  assign _2719_ = state_in[47:40] == 7'b1110101;
  assign _2720_ = state_in[47:40] == 7'b1110100;
  assign _2721_ = state_in[47:40] == 7'b1110011;
  assign _2722_ = state_in[47:40] == 7'b1110010;
  assign _2723_ = state_in[47:40] == 7'b1110001;
  assign _2724_ = state_in[47:40] == 7'b1110000;
  assign _2725_ = state_in[47:40] == 7'b1101111;
  assign _2726_ = state_in[47:40] == 7'b1101110;
  assign _2727_ = state_in[47:40] == 7'b1101101;
  assign _2728_ = state_in[47:40] == 7'b1101100;
  assign _2729_ = state_in[47:40] == 7'b1101011;
  assign _2730_ = state_in[47:40] == 7'b1101010;
  assign _2731_ = state_in[47:40] == 7'b1101001;
  assign _2732_ = state_in[47:40] == 7'b1101000;
  assign _2733_ = state_in[47:40] == 7'b1100111;
  assign _2734_ = state_in[47:40] == 7'b1100110;
  assign _2735_ = state_in[47:40] == 7'b1100101;
  assign _2736_ = state_in[47:40] == 7'b1100100;
  assign _2737_ = state_in[47:40] == 7'b1100011;
  assign _2738_ = state_in[47:40] == 7'b1100010;
  assign _2739_ = state_in[47:40] == 7'b1100001;
  assign _2740_ = state_in[47:40] == 7'b1100000;
  assign _2741_ = state_in[47:40] == 7'b1011111;
  assign _2742_ = state_in[47:40] == 7'b1011110;
  assign _2743_ = state_in[47:40] == 7'b1011101;
  assign _2744_ = state_in[47:40] == 7'b1011100;
  assign _2745_ = state_in[47:40] == 7'b1011011;
  assign _2746_ = state_in[47:40] == 7'b1011010;
  assign _2747_ = state_in[47:40] == 7'b1011001;
  assign _2748_ = state_in[47:40] == 7'b1011000;
  assign _2749_ = state_in[47:40] == 7'b1010111;
  assign _2750_ = state_in[47:40] == 7'b1010110;
  assign _2751_ = state_in[47:40] == 7'b1010101;
  assign _2752_ = state_in[47:40] == 7'b1010100;
  assign _2753_ = state_in[47:40] == 7'b1010011;
  assign _2754_ = state_in[47:40] == 7'b1010010;
  assign _2755_ = state_in[47:40] == 7'b1010001;
  assign _2756_ = state_in[47:40] == 7'b1010000;
  assign _2757_ = state_in[47:40] == 7'b1001111;
  assign _2758_ = state_in[47:40] == 7'b1001110;
  assign _2759_ = state_in[47:40] == 7'b1001101;
  assign _2760_ = state_in[47:40] == 7'b1001100;
  assign _2761_ = state_in[47:40] == 7'b1001011;
  assign _2762_ = state_in[47:40] == 7'b1001010;
  assign _2763_ = state_in[47:40] == 7'b1001001;
  assign _2764_ = state_in[47:40] == 7'b1001000;
  assign _2765_ = state_in[47:40] == 7'b1000111;
  assign _2766_ = state_in[47:40] == 7'b1000110;
  assign _2767_ = state_in[47:40] == 7'b1000101;
  assign _2768_ = state_in[47:40] == 7'b1000100;
  assign _2769_ = state_in[47:40] == 7'b1000011;
  assign _2770_ = state_in[47:40] == 7'b1000010;
  assign _2771_ = state_in[47:40] == 7'b1000001;
  assign _2772_ = state_in[47:40] == 7'b1000000;
  assign _2773_ = state_in[47:40] == 6'b111111;
  assign _2774_ = state_in[47:40] == 6'b111110;
  assign _2775_ = state_in[47:40] == 6'b111101;
  assign _2776_ = state_in[47:40] == 6'b111100;
  assign _2777_ = state_in[47:40] == 6'b111011;
  assign _2778_ = state_in[47:40] == 6'b111010;
  assign _2779_ = state_in[47:40] == 6'b111001;
  assign _2780_ = state_in[47:40] == 6'b111000;
  assign _2781_ = state_in[47:40] == 6'b110111;
  assign _2782_ = state_in[47:40] == 6'b110110;
  assign _2783_ = state_in[47:40] == 6'b110101;
  assign _2784_ = state_in[47:40] == 6'b110100;
  assign _2785_ = state_in[47:40] == 6'b110011;
  assign _2786_ = state_in[47:40] == 6'b110010;
  assign _2787_ = state_in[47:40] == 6'b110001;
  assign _2788_ = state_in[47:40] == 6'b110000;
  assign _2789_ = state_in[47:40] == 6'b101111;
  assign _2790_ = state_in[47:40] == 6'b101110;
  assign _2791_ = state_in[47:40] == 6'b101101;
  assign _2792_ = state_in[47:40] == 6'b101100;
  assign _2793_ = state_in[47:40] == 6'b101011;
  assign _2794_ = state_in[47:40] == 6'b101010;
  assign _2795_ = state_in[47:40] == 6'b101001;
  assign _2796_ = state_in[47:40] == 6'b101000;
  assign _2797_ = state_in[47:40] == 6'b100111;
  assign _2798_ = state_in[47:40] == 6'b100110;
  assign _2799_ = state_in[47:40] == 6'b100101;
  assign _2800_ = state_in[47:40] == 6'b100100;
  assign _2801_ = state_in[47:40] == 6'b100011;
  assign _2802_ = state_in[47:40] == 6'b100010;
  assign _2803_ = state_in[47:40] == 6'b100001;
  assign _2804_ = state_in[47:40] == 6'b100000;
  assign _2805_ = state_in[47:40] == 5'b11111;
  assign _2806_ = state_in[47:40] == 5'b11110;
  assign _2807_ = state_in[47:40] == 5'b11101;
  assign _2808_ = state_in[47:40] == 5'b11100;
  assign _2809_ = state_in[47:40] == 5'b11011;
  assign _2810_ = state_in[47:40] == 5'b11010;
  assign _2811_ = state_in[47:40] == 5'b11001;
  assign _2812_ = state_in[47:40] == 5'b11000;
  assign _2813_ = state_in[47:40] == 5'b10111;
  assign _2814_ = state_in[47:40] == 5'b10110;
  assign _2815_ = state_in[47:40] == 5'b10101;
  assign _2816_ = state_in[47:40] == 5'b10100;
  assign _2817_ = state_in[47:40] == 5'b10011;
  assign _2818_ = state_in[47:40] == 5'b10010;
  assign _2819_ = state_in[47:40] == 5'b10001;
  assign _2820_ = state_in[47:40] == 5'b10000;
  assign _2821_ = state_in[47:40] == 4'b1111;
  assign _2822_ = state_in[47:40] == 4'b1110;
  assign _2823_ = state_in[47:40] == 4'b1101;
  assign _2824_ = state_in[47:40] == 4'b1100;
  assign _2825_ = state_in[47:40] == 4'b1011;
  assign _2826_ = state_in[47:40] == 4'b1010;
  assign _2827_ = state_in[47:40] == 4'b1001;
  assign _2828_ = state_in[47:40] == 4'b1000;
  assign _2829_ = state_in[47:40] == 3'b111;
  assign _2830_ = state_in[47:40] == 3'b110;
  assign _2831_ = state_in[47:40] == 3'b101;
  assign _2832_ = state_in[47:40] == 3'b100;
  assign _2833_ = state_in[47:40] == 2'b11;
  assign _2834_ = state_in[47:40] == 2'b10;
  assign _2835_ = state_in[47:40] == 1'b1;
  assign _2836_ = ! state_in[47:40];
  always @(posedge clk)
      \t2.t2.s4.out <= _2837_;
  logic [255:0] fangyuan22;
  assign fangyuan22 = { _2836_, _2835_, _2834_, _2833_, _2832_, _2831_, _2830_, _2829_, _2828_, _2827_, _2826_, _2825_, _2824_, _2823_, _2822_, _2821_, _2820_, _2819_, _2818_, _2817_, _2816_, _2815_, _2814_, _2813_, _2812_, _2811_, _2810_, _2809_, _2808_, _2807_, _2806_, _2805_, _2804_, _2803_, _2802_, _2801_, _2800_, _2799_, _2798_, _2797_, _2796_, _2795_, _2794_, _2793_, _2792_, _2791_, _2790_, _2789_, _2788_, _2787_, _2786_, _2785_, _2784_, _2783_, _2782_, _2781_, _2780_, _2779_, _2778_, _2777_, _2776_, _2775_, _2774_, _2773_, _2772_, _2771_, _2770_, _2769_, _2768_, _2767_, _2766_, _2765_, _2764_, _2763_, _2762_, _2761_, _2760_, _2759_, _2758_, _2757_, _2756_, _2755_, _2754_, _2753_, _2752_, _2751_, _2750_, _2749_, _2748_, _2747_, _2746_, _2745_, _2744_, _2743_, _2742_, _2741_, _2740_, _2739_, _2738_, _2737_, _2736_, _2735_, _2734_, _2733_, _2732_, _2731_, _2730_, _2729_, _2728_, _2727_, _2726_, _2725_, _2724_, _2723_, _2722_, _2721_, _2720_, _2719_, _2718_, _2717_, _2716_, _2715_, _2714_, _2713_, _2712_, _2711_, _2710_, _2709_, _2708_, _2707_, _2706_, _2705_, _2704_, _2703_, _2702_, _2701_, _2700_, _2699_, _2698_, _2697_, _2696_, _2695_, _2694_, _2693_, _2692_, _2691_, _2690_, _2689_, _2688_, _2687_, _2686_, _2685_, _2684_, _2683_, _2682_, _2681_, _2680_, _2679_, _2678_, _2677_, _2676_, _2675_, _2674_, _2673_, _2672_, _2671_, _2670_, _2669_, _2668_, _2667_, _2666_, _2665_, _2664_, _2663_, _2662_, _2661_, _2660_, _2659_, _2658_, _2657_, _2656_, _2655_, _2654_, _2653_, _2652_, _2651_, _2650_, _2649_, _2648_, _2647_, _2646_, _2645_, _2644_, _2643_, _2642_, _2641_, _2640_, _2639_, _2638_, _2637_, _2636_, _2635_, _2634_, _2633_, _2632_, _2631_, _2630_, _2629_, _2628_, _2627_, _2626_, _2625_, _2624_, _2623_, _2622_, _2621_, _2620_, _2619_, _2618_, _2617_, _2616_, _2615_, _2614_, _2613_, _2612_, _2611_, _2610_, _2609_, _2608_, _2607_, _2606_, _2605_, _2604_, _2603_, _2602_, _2601_, _2600_, _2599_, _2598_, _2597_, _2596_, _2595_, _2594_, _2593_, _2592_, _2591_, _2590_, _2589_, _2588_, _2587_, _2586_, _2585_, _2584_, _2583_, _2582_, _2581_ };

  always @(\t2.t2.s4.out or fangyuan22) begin
    casez (fangyuan22)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2837_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2837_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2837_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2837_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2837_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2837_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2837_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2837_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2837_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2837_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2837_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2837_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2837_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2837_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2837_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2837_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2837_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2837_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2837_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2837_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2837_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2837_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2837_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2837_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2837_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2837_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2837_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2837_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2837_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2837_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2837_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2837_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2837_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2837_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2837_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2837_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2837_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2837_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2837_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2837_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2837_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2837_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2837_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2837_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2837_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2837_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2837_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2837_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2837_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2837_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2837_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2837_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2837_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2837_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2837_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2837_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2837_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2837_ = 8'b11000110 ;
      default:
        _2837_ = \t2.t2.s4.out ;
    endcase
  end
  assign p23[15:8] = \t2.t3.s0.out ^ \t2.t3.s4.out ;
  always @(posedge clk)
      \t2.t3.s0.out <= _2838_;
  logic [255:0] fangyuan23;
  assign fangyuan23 = { _3094_, _3093_, _3092_, _3091_, _3090_, _3089_, _3088_, _3087_, _3086_, _3085_, _3084_, _3083_, _3082_, _3081_, _3080_, _3079_, _3078_, _3077_, _3076_, _3075_, _3074_, _3073_, _3072_, _3071_, _3070_, _3069_, _3068_, _3067_, _3066_, _3065_, _3064_, _3063_, _3062_, _3061_, _3060_, _3059_, _3058_, _3057_, _3056_, _3055_, _3054_, _3053_, _3052_, _3051_, _3050_, _3049_, _3048_, _3047_, _3046_, _3045_, _3044_, _3043_, _3042_, _3041_, _3040_, _3039_, _3038_, _3037_, _3036_, _3035_, _3034_, _3033_, _3032_, _3031_, _3030_, _3029_, _3028_, _3027_, _3026_, _3025_, _3024_, _3023_, _3022_, _3021_, _3020_, _3019_, _3018_, _3017_, _3016_, _3015_, _3014_, _3013_, _3012_, _3011_, _3010_, _3009_, _3008_, _3007_, _3006_, _3005_, _3004_, _3003_, _3002_, _3001_, _3000_, _2999_, _2998_, _2997_, _2996_, _2995_, _2994_, _2993_, _2992_, _2991_, _2990_, _2989_, _2988_, _2987_, _2986_, _2985_, _2984_, _2983_, _2982_, _2981_, _2980_, _2979_, _2978_, _2977_, _2976_, _2975_, _2974_, _2973_, _2972_, _2971_, _2970_, _2969_, _2968_, _2967_, _2966_, _2965_, _2964_, _2963_, _2962_, _2961_, _2960_, _2959_, _2958_, _2957_, _2956_, _2955_, _2954_, _2953_, _2952_, _2951_, _2950_, _2949_, _2948_, _2947_, _2946_, _2945_, _2944_, _2943_, _2942_, _2941_, _2940_, _2939_, _2938_, _2937_, _2936_, _2935_, _2934_, _2933_, _2932_, _2931_, _2930_, _2929_, _2928_, _2927_, _2926_, _2925_, _2924_, _2923_, _2922_, _2921_, _2920_, _2919_, _2918_, _2917_, _2916_, _2915_, _2914_, _2913_, _2912_, _2911_, _2910_, _2909_, _2908_, _2907_, _2906_, _2905_, _2904_, _2903_, _2902_, _2901_, _2900_, _2899_, _2898_, _2897_, _2896_, _2895_, _2894_, _2893_, _2892_, _2891_, _2890_, _2889_, _2888_, _2887_, _2886_, _2885_, _2884_, _2883_, _2882_, _2881_, _2880_, _2879_, _2878_, _2877_, _2876_, _2875_, _2874_, _2873_, _2872_, _2871_, _2870_, _2869_, _2868_, _2867_, _2866_, _2865_, _2864_, _2863_, _2862_, _2861_, _2860_, _2859_, _2858_, _2857_, _2856_, _2855_, _2854_, _2853_, _2852_, _2851_, _2850_, _2849_, _2848_, _2847_, _2846_, _2845_, _2844_, _2843_, _2842_, _2841_, _2840_, _2839_ };

  always @(\t2.t3.s0.out or fangyuan23) begin
    casez (fangyuan23)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _2838_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _2838_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _2838_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _2838_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _2838_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _2838_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _2838_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _2838_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _2838_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _2838_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _2838_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _2838_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _2838_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _2838_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _2838_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _2838_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _2838_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _2838_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _2838_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _2838_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _2838_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _2838_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _2838_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _2838_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _2838_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _2838_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _2838_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _2838_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _2838_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _2838_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _2838_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _2838_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _2838_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _2838_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _2838_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _2838_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _2838_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _2838_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _2838_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _2838_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _2838_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _2838_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _2838_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _2838_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _2838_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _2838_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _2838_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _2838_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _2838_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _2838_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _2838_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _2838_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _2838_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _2838_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _2838_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _2838_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _2838_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _2838_ = 8'b01100011 ;
      default:
        _2838_ = \t2.t3.s0.out ;
    endcase
  end
  assign _2839_ = state_in[39:32] == 8'b11111111;
  assign _2840_ = state_in[39:32] == 8'b11111110;
  assign _2841_ = state_in[39:32] == 8'b11111101;
  assign _2842_ = state_in[39:32] == 8'b11111100;
  assign _2843_ = state_in[39:32] == 8'b11111011;
  assign _2844_ = state_in[39:32] == 8'b11111010;
  assign _2845_ = state_in[39:32] == 8'b11111001;
  assign _2846_ = state_in[39:32] == 8'b11111000;
  assign _2847_ = state_in[39:32] == 8'b11110111;
  assign _2848_ = state_in[39:32] == 8'b11110110;
  assign _2849_ = state_in[39:32] == 8'b11110101;
  assign _2850_ = state_in[39:32] == 8'b11110100;
  assign _2851_ = state_in[39:32] == 8'b11110011;
  assign _2852_ = state_in[39:32] == 8'b11110010;
  assign _2853_ = state_in[39:32] == 8'b11110001;
  assign _2854_ = state_in[39:32] == 8'b11110000;
  assign _2855_ = state_in[39:32] == 8'b11101111;
  assign _2856_ = state_in[39:32] == 8'b11101110;
  assign _2857_ = state_in[39:32] == 8'b11101101;
  assign _2858_ = state_in[39:32] == 8'b11101100;
  assign _2859_ = state_in[39:32] == 8'b11101011;
  assign _2860_ = state_in[39:32] == 8'b11101010;
  assign _2861_ = state_in[39:32] == 8'b11101001;
  assign _2862_ = state_in[39:32] == 8'b11101000;
  assign _2863_ = state_in[39:32] == 8'b11100111;
  assign _2864_ = state_in[39:32] == 8'b11100110;
  assign _2865_ = state_in[39:32] == 8'b11100101;
  assign _2866_ = state_in[39:32] == 8'b11100100;
  assign _2867_ = state_in[39:32] == 8'b11100011;
  assign _2868_ = state_in[39:32] == 8'b11100010;
  assign _2869_ = state_in[39:32] == 8'b11100001;
  assign _2870_ = state_in[39:32] == 8'b11100000;
  assign _2871_ = state_in[39:32] == 8'b11011111;
  assign _2872_ = state_in[39:32] == 8'b11011110;
  assign _2873_ = state_in[39:32] == 8'b11011101;
  assign _2874_ = state_in[39:32] == 8'b11011100;
  assign _2875_ = state_in[39:32] == 8'b11011011;
  assign _2876_ = state_in[39:32] == 8'b11011010;
  assign _2877_ = state_in[39:32] == 8'b11011001;
  assign _2878_ = state_in[39:32] == 8'b11011000;
  assign _2879_ = state_in[39:32] == 8'b11010111;
  assign _2880_ = state_in[39:32] == 8'b11010110;
  assign _2881_ = state_in[39:32] == 8'b11010101;
  assign _2882_ = state_in[39:32] == 8'b11010100;
  assign _2883_ = state_in[39:32] == 8'b11010011;
  assign _2884_ = state_in[39:32] == 8'b11010010;
  assign _2885_ = state_in[39:32] == 8'b11010001;
  assign _2886_ = state_in[39:32] == 8'b11010000;
  assign _2887_ = state_in[39:32] == 8'b11001111;
  assign _2888_ = state_in[39:32] == 8'b11001110;
  assign _2889_ = state_in[39:32] == 8'b11001101;
  assign _2890_ = state_in[39:32] == 8'b11001100;
  assign _2891_ = state_in[39:32] == 8'b11001011;
  assign _2892_ = state_in[39:32] == 8'b11001010;
  assign _2893_ = state_in[39:32] == 8'b11001001;
  assign _2894_ = state_in[39:32] == 8'b11001000;
  assign _2895_ = state_in[39:32] == 8'b11000111;
  assign _2896_ = state_in[39:32] == 8'b11000110;
  assign _2897_ = state_in[39:32] == 8'b11000101;
  assign _2898_ = state_in[39:32] == 8'b11000100;
  assign _2899_ = state_in[39:32] == 8'b11000011;
  assign _2900_ = state_in[39:32] == 8'b11000010;
  assign _2901_ = state_in[39:32] == 8'b11000001;
  assign _2902_ = state_in[39:32] == 8'b11000000;
  assign _2903_ = state_in[39:32] == 8'b10111111;
  assign _2904_ = state_in[39:32] == 8'b10111110;
  assign _2905_ = state_in[39:32] == 8'b10111101;
  assign _2906_ = state_in[39:32] == 8'b10111100;
  assign _2907_ = state_in[39:32] == 8'b10111011;
  assign _2908_ = state_in[39:32] == 8'b10111010;
  assign _2909_ = state_in[39:32] == 8'b10111001;
  assign _2910_ = state_in[39:32] == 8'b10111000;
  assign _2911_ = state_in[39:32] == 8'b10110111;
  assign _2912_ = state_in[39:32] == 8'b10110110;
  assign _2913_ = state_in[39:32] == 8'b10110101;
  assign _2914_ = state_in[39:32] == 8'b10110100;
  assign _2915_ = state_in[39:32] == 8'b10110011;
  assign _2916_ = state_in[39:32] == 8'b10110010;
  assign _2917_ = state_in[39:32] == 8'b10110001;
  assign _2918_ = state_in[39:32] == 8'b10110000;
  assign _2919_ = state_in[39:32] == 8'b10101111;
  assign _2920_ = state_in[39:32] == 8'b10101110;
  assign _2921_ = state_in[39:32] == 8'b10101101;
  assign _2922_ = state_in[39:32] == 8'b10101100;
  assign _2923_ = state_in[39:32] == 8'b10101011;
  assign _2924_ = state_in[39:32] == 8'b10101010;
  assign _2925_ = state_in[39:32] == 8'b10101001;
  assign _2926_ = state_in[39:32] == 8'b10101000;
  assign _2927_ = state_in[39:32] == 8'b10100111;
  assign _2928_ = state_in[39:32] == 8'b10100110;
  assign _2929_ = state_in[39:32] == 8'b10100101;
  assign _2930_ = state_in[39:32] == 8'b10100100;
  assign _2931_ = state_in[39:32] == 8'b10100011;
  assign _2932_ = state_in[39:32] == 8'b10100010;
  assign _2933_ = state_in[39:32] == 8'b10100001;
  assign _2934_ = state_in[39:32] == 8'b10100000;
  assign _2935_ = state_in[39:32] == 8'b10011111;
  assign _2936_ = state_in[39:32] == 8'b10011110;
  assign _2937_ = state_in[39:32] == 8'b10011101;
  assign _2938_ = state_in[39:32] == 8'b10011100;
  assign _2939_ = state_in[39:32] == 8'b10011011;
  assign _2940_ = state_in[39:32] == 8'b10011010;
  assign _2941_ = state_in[39:32] == 8'b10011001;
  assign _2942_ = state_in[39:32] == 8'b10011000;
  assign _2943_ = state_in[39:32] == 8'b10010111;
  assign _2944_ = state_in[39:32] == 8'b10010110;
  assign _2945_ = state_in[39:32] == 8'b10010101;
  assign _2946_ = state_in[39:32] == 8'b10010100;
  assign _2947_ = state_in[39:32] == 8'b10010011;
  assign _2948_ = state_in[39:32] == 8'b10010010;
  assign _2949_ = state_in[39:32] == 8'b10010001;
  assign _2950_ = state_in[39:32] == 8'b10010000;
  assign _2951_ = state_in[39:32] == 8'b10001111;
  assign _2952_ = state_in[39:32] == 8'b10001110;
  assign _2953_ = state_in[39:32] == 8'b10001101;
  assign _2954_ = state_in[39:32] == 8'b10001100;
  assign _2955_ = state_in[39:32] == 8'b10001011;
  assign _2956_ = state_in[39:32] == 8'b10001010;
  assign _2957_ = state_in[39:32] == 8'b10001001;
  assign _2958_ = state_in[39:32] == 8'b10001000;
  assign _2959_ = state_in[39:32] == 8'b10000111;
  assign _2960_ = state_in[39:32] == 8'b10000110;
  assign _2961_ = state_in[39:32] == 8'b10000101;
  assign _2962_ = state_in[39:32] == 8'b10000100;
  assign _2963_ = state_in[39:32] == 8'b10000011;
  assign _2964_ = state_in[39:32] == 8'b10000010;
  assign _2965_ = state_in[39:32] == 8'b10000001;
  assign _2966_ = state_in[39:32] == 8'b10000000;
  assign _2967_ = state_in[39:32] == 7'b1111111;
  assign _2968_ = state_in[39:32] == 7'b1111110;
  assign _2969_ = state_in[39:32] == 7'b1111101;
  assign _2970_ = state_in[39:32] == 7'b1111100;
  assign _2971_ = state_in[39:32] == 7'b1111011;
  assign _2972_ = state_in[39:32] == 7'b1111010;
  assign _2973_ = state_in[39:32] == 7'b1111001;
  assign _2974_ = state_in[39:32] == 7'b1111000;
  assign _2975_ = state_in[39:32] == 7'b1110111;
  assign _2976_ = state_in[39:32] == 7'b1110110;
  assign _2977_ = state_in[39:32] == 7'b1110101;
  assign _2978_ = state_in[39:32] == 7'b1110100;
  assign _2979_ = state_in[39:32] == 7'b1110011;
  assign _2980_ = state_in[39:32] == 7'b1110010;
  assign _2981_ = state_in[39:32] == 7'b1110001;
  assign _2982_ = state_in[39:32] == 7'b1110000;
  assign _2983_ = state_in[39:32] == 7'b1101111;
  assign _2984_ = state_in[39:32] == 7'b1101110;
  assign _2985_ = state_in[39:32] == 7'b1101101;
  assign _2986_ = state_in[39:32] == 7'b1101100;
  assign _2987_ = state_in[39:32] == 7'b1101011;
  assign _2988_ = state_in[39:32] == 7'b1101010;
  assign _2989_ = state_in[39:32] == 7'b1101001;
  assign _2990_ = state_in[39:32] == 7'b1101000;
  assign _2991_ = state_in[39:32] == 7'b1100111;
  assign _2992_ = state_in[39:32] == 7'b1100110;
  assign _2993_ = state_in[39:32] == 7'b1100101;
  assign _2994_ = state_in[39:32] == 7'b1100100;
  assign _2995_ = state_in[39:32] == 7'b1100011;
  assign _2996_ = state_in[39:32] == 7'b1100010;
  assign _2997_ = state_in[39:32] == 7'b1100001;
  assign _2998_ = state_in[39:32] == 7'b1100000;
  assign _2999_ = state_in[39:32] == 7'b1011111;
  assign _3000_ = state_in[39:32] == 7'b1011110;
  assign _3001_ = state_in[39:32] == 7'b1011101;
  assign _3002_ = state_in[39:32] == 7'b1011100;
  assign _3003_ = state_in[39:32] == 7'b1011011;
  assign _3004_ = state_in[39:32] == 7'b1011010;
  assign _3005_ = state_in[39:32] == 7'b1011001;
  assign _3006_ = state_in[39:32] == 7'b1011000;
  assign _3007_ = state_in[39:32] == 7'b1010111;
  assign _3008_ = state_in[39:32] == 7'b1010110;
  assign _3009_ = state_in[39:32] == 7'b1010101;
  assign _3010_ = state_in[39:32] == 7'b1010100;
  assign _3011_ = state_in[39:32] == 7'b1010011;
  assign _3012_ = state_in[39:32] == 7'b1010010;
  assign _3013_ = state_in[39:32] == 7'b1010001;
  assign _3014_ = state_in[39:32] == 7'b1010000;
  assign _3015_ = state_in[39:32] == 7'b1001111;
  assign _3016_ = state_in[39:32] == 7'b1001110;
  assign _3017_ = state_in[39:32] == 7'b1001101;
  assign _3018_ = state_in[39:32] == 7'b1001100;
  assign _3019_ = state_in[39:32] == 7'b1001011;
  assign _3020_ = state_in[39:32] == 7'b1001010;
  assign _3021_ = state_in[39:32] == 7'b1001001;
  assign _3022_ = state_in[39:32] == 7'b1001000;
  assign _3023_ = state_in[39:32] == 7'b1000111;
  assign _3024_ = state_in[39:32] == 7'b1000110;
  assign _3025_ = state_in[39:32] == 7'b1000101;
  assign _3026_ = state_in[39:32] == 7'b1000100;
  assign _3027_ = state_in[39:32] == 7'b1000011;
  assign _3028_ = state_in[39:32] == 7'b1000010;
  assign _3029_ = state_in[39:32] == 7'b1000001;
  assign _3030_ = state_in[39:32] == 7'b1000000;
  assign _3031_ = state_in[39:32] == 6'b111111;
  assign _3032_ = state_in[39:32] == 6'b111110;
  assign _3033_ = state_in[39:32] == 6'b111101;
  assign _3034_ = state_in[39:32] == 6'b111100;
  assign _3035_ = state_in[39:32] == 6'b111011;
  assign _3036_ = state_in[39:32] == 6'b111010;
  assign _3037_ = state_in[39:32] == 6'b111001;
  assign _3038_ = state_in[39:32] == 6'b111000;
  assign _3039_ = state_in[39:32] == 6'b110111;
  assign _3040_ = state_in[39:32] == 6'b110110;
  assign _3041_ = state_in[39:32] == 6'b110101;
  assign _3042_ = state_in[39:32] == 6'b110100;
  assign _3043_ = state_in[39:32] == 6'b110011;
  assign _3044_ = state_in[39:32] == 6'b110010;
  assign _3045_ = state_in[39:32] == 6'b110001;
  assign _3046_ = state_in[39:32] == 6'b110000;
  assign _3047_ = state_in[39:32] == 6'b101111;
  assign _3048_ = state_in[39:32] == 6'b101110;
  assign _3049_ = state_in[39:32] == 6'b101101;
  assign _3050_ = state_in[39:32] == 6'b101100;
  assign _3051_ = state_in[39:32] == 6'b101011;
  assign _3052_ = state_in[39:32] == 6'b101010;
  assign _3053_ = state_in[39:32] == 6'b101001;
  assign _3054_ = state_in[39:32] == 6'b101000;
  assign _3055_ = state_in[39:32] == 6'b100111;
  assign _3056_ = state_in[39:32] == 6'b100110;
  assign _3057_ = state_in[39:32] == 6'b100101;
  assign _3058_ = state_in[39:32] == 6'b100100;
  assign _3059_ = state_in[39:32] == 6'b100011;
  assign _3060_ = state_in[39:32] == 6'b100010;
  assign _3061_ = state_in[39:32] == 6'b100001;
  assign _3062_ = state_in[39:32] == 6'b100000;
  assign _3063_ = state_in[39:32] == 5'b11111;
  assign _3064_ = state_in[39:32] == 5'b11110;
  assign _3065_ = state_in[39:32] == 5'b11101;
  assign _3066_ = state_in[39:32] == 5'b11100;
  assign _3067_ = state_in[39:32] == 5'b11011;
  assign _3068_ = state_in[39:32] == 5'b11010;
  assign _3069_ = state_in[39:32] == 5'b11001;
  assign _3070_ = state_in[39:32] == 5'b11000;
  assign _3071_ = state_in[39:32] == 5'b10111;
  assign _3072_ = state_in[39:32] == 5'b10110;
  assign _3073_ = state_in[39:32] == 5'b10101;
  assign _3074_ = state_in[39:32] == 5'b10100;
  assign _3075_ = state_in[39:32] == 5'b10011;
  assign _3076_ = state_in[39:32] == 5'b10010;
  assign _3077_ = state_in[39:32] == 5'b10001;
  assign _3078_ = state_in[39:32] == 5'b10000;
  assign _3079_ = state_in[39:32] == 4'b1111;
  assign _3080_ = state_in[39:32] == 4'b1110;
  assign _3081_ = state_in[39:32] == 4'b1101;
  assign _3082_ = state_in[39:32] == 4'b1100;
  assign _3083_ = state_in[39:32] == 4'b1011;
  assign _3084_ = state_in[39:32] == 4'b1010;
  assign _3085_ = state_in[39:32] == 4'b1001;
  assign _3086_ = state_in[39:32] == 4'b1000;
  assign _3087_ = state_in[39:32] == 3'b111;
  assign _3088_ = state_in[39:32] == 3'b110;
  assign _3089_ = state_in[39:32] == 3'b101;
  assign _3090_ = state_in[39:32] == 3'b100;
  assign _3091_ = state_in[39:32] == 2'b11;
  assign _3092_ = state_in[39:32] == 2'b10;
  assign _3093_ = state_in[39:32] == 1'b1;
  assign _3094_ = ! state_in[39:32];
  always @(posedge clk)
      \t2.t3.s4.out <= _3095_;
  logic [255:0] fangyuan24;
  assign fangyuan24 = { _3094_, _3093_, _3092_, _3091_, _3090_, _3089_, _3088_, _3087_, _3086_, _3085_, _3084_, _3083_, _3082_, _3081_, _3080_, _3079_, _3078_, _3077_, _3076_, _3075_, _3074_, _3073_, _3072_, _3071_, _3070_, _3069_, _3068_, _3067_, _3066_, _3065_, _3064_, _3063_, _3062_, _3061_, _3060_, _3059_, _3058_, _3057_, _3056_, _3055_, _3054_, _3053_, _3052_, _3051_, _3050_, _3049_, _3048_, _3047_, _3046_, _3045_, _3044_, _3043_, _3042_, _3041_, _3040_, _3039_, _3038_, _3037_, _3036_, _3035_, _3034_, _3033_, _3032_, _3031_, _3030_, _3029_, _3028_, _3027_, _3026_, _3025_, _3024_, _3023_, _3022_, _3021_, _3020_, _3019_, _3018_, _3017_, _3016_, _3015_, _3014_, _3013_, _3012_, _3011_, _3010_, _3009_, _3008_, _3007_, _3006_, _3005_, _3004_, _3003_, _3002_, _3001_, _3000_, _2999_, _2998_, _2997_, _2996_, _2995_, _2994_, _2993_, _2992_, _2991_, _2990_, _2989_, _2988_, _2987_, _2986_, _2985_, _2984_, _2983_, _2982_, _2981_, _2980_, _2979_, _2978_, _2977_, _2976_, _2975_, _2974_, _2973_, _2972_, _2971_, _2970_, _2969_, _2968_, _2967_, _2966_, _2965_, _2964_, _2963_, _2962_, _2961_, _2960_, _2959_, _2958_, _2957_, _2956_, _2955_, _2954_, _2953_, _2952_, _2951_, _2950_, _2949_, _2948_, _2947_, _2946_, _2945_, _2944_, _2943_, _2942_, _2941_, _2940_, _2939_, _2938_, _2937_, _2936_, _2935_, _2934_, _2933_, _2932_, _2931_, _2930_, _2929_, _2928_, _2927_, _2926_, _2925_, _2924_, _2923_, _2922_, _2921_, _2920_, _2919_, _2918_, _2917_, _2916_, _2915_, _2914_, _2913_, _2912_, _2911_, _2910_, _2909_, _2908_, _2907_, _2906_, _2905_, _2904_, _2903_, _2902_, _2901_, _2900_, _2899_, _2898_, _2897_, _2896_, _2895_, _2894_, _2893_, _2892_, _2891_, _2890_, _2889_, _2888_, _2887_, _2886_, _2885_, _2884_, _2883_, _2882_, _2881_, _2880_, _2879_, _2878_, _2877_, _2876_, _2875_, _2874_, _2873_, _2872_, _2871_, _2870_, _2869_, _2868_, _2867_, _2866_, _2865_, _2864_, _2863_, _2862_, _2861_, _2860_, _2859_, _2858_, _2857_, _2856_, _2855_, _2854_, _2853_, _2852_, _2851_, _2850_, _2849_, _2848_, _2847_, _2846_, _2845_, _2844_, _2843_, _2842_, _2841_, _2840_, _2839_ };

  always @(\t2.t3.s4.out or fangyuan24) begin
    casez (fangyuan24)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3095_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3095_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3095_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3095_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3095_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3095_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3095_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3095_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3095_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3095_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3095_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3095_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3095_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3095_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3095_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3095_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3095_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3095_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3095_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3095_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3095_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3095_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3095_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3095_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3095_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3095_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3095_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3095_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3095_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3095_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3095_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3095_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3095_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3095_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3095_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3095_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3095_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3095_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3095_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3095_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3095_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3095_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3095_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3095_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3095_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3095_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3095_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3095_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3095_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3095_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3095_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3095_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3095_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3095_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3095_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3095_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3095_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3095_ = 8'b11000110 ;
      default:
        _3095_ = \t2.t3.s4.out ;
    endcase
  end
  assign p30[7:0] = \t3.t0.s0.out ^ \t3.t0.s4.out ;
  always @(posedge clk)
      \t3.t0.s0.out <= _3096_;
  logic [255:0] fangyuan25;
  assign fangyuan25 = { _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_, _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_, _3309_, _3308_, _3307_, _3306_, _3305_, _3304_, _3303_, _3302_, _3301_, _3300_, _3299_, _3298_, _3297_, _3296_, _3295_, _3294_, _3293_, _3292_, _3291_, _3290_, _3289_, _3288_, _3287_, _3286_, _3285_, _3284_, _3283_, _3282_, _3281_, _3280_, _3279_, _3278_, _3277_, _3276_, _3275_, _3274_, _3273_, _3272_, _3271_, _3270_, _3269_, _3268_, _3267_, _3266_, _3265_, _3264_, _3263_, _3262_, _3261_, _3260_, _3259_, _3258_, _3257_, _3256_, _3255_, _3254_, _3253_, _3252_, _3251_, _3250_, _3249_, _3248_, _3247_, _3246_, _3245_, _3244_, _3243_, _3242_, _3241_, _3240_, _3239_, _3238_, _3237_, _3236_, _3235_, _3234_, _3233_, _3232_, _3231_, _3230_, _3229_, _3228_, _3227_, _3226_, _3225_, _3224_, _3223_, _3222_, _3221_, _3220_, _3219_, _3218_, _3217_, _3216_, _3215_, _3214_, _3213_, _3212_, _3211_, _3210_, _3209_, _3208_, _3207_, _3206_, _3205_, _3204_, _3203_, _3202_, _3201_, _3200_, _3199_, _3198_, _3197_, _3196_, _3195_, _3194_, _3193_, _3192_, _3191_, _3190_, _3189_, _3188_, _3187_, _3186_, _3185_, _3184_, _3183_, _3182_, _3181_, _3180_, _3179_, _3178_, _3177_, _3176_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3169_, _3168_, _3167_, _3166_, _3165_, _3164_, _3163_, _3162_, _3161_, _3160_, _3159_, _3158_, _3157_, _3156_, _3155_, _3154_, _3153_, _3152_, _3151_, _3150_, _3149_, _3148_, _3147_, _3146_, _3145_, _3144_, _3143_, _3142_, _3141_, _3140_, _3139_, _3138_, _3137_, _3136_, _3135_, _3134_, _3133_, _3132_, _3131_, _3130_, _3129_, _3128_, _3127_, _3126_, _3125_, _3124_, _3123_, _3122_, _3121_, _3120_, _3119_, _3118_, _3117_, _3116_, _3115_, _3114_, _3113_, _3112_, _3111_, _3110_, _3109_, _3108_, _3107_, _3106_, _3105_, _3104_, _3103_, _3102_, _3101_, _3100_, _3099_, _3098_, _3097_ };

  always @(\t3.t0.s0.out or fangyuan25) begin
    casez (fangyuan25)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3096_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3096_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3096_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3096_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3096_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3096_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3096_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3096_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3096_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3096_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3096_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3096_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3096_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3096_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3096_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3096_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3096_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3096_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3096_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3096_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3096_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3096_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3096_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3096_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3096_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3096_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3096_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3096_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3096_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3096_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3096_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3096_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3096_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3096_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3096_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3096_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3096_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3096_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3096_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3096_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3096_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3096_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3096_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3096_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3096_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3096_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3096_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3096_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3096_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3096_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3096_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3096_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3096_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3096_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3096_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3096_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3096_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3096_ = 8'b01100011 ;
      default:
        _3096_ = \t3.t0.s0.out ;
    endcase
  end
  assign _3097_ = state_in[31:24] == 8'b11111111;
  assign _3098_ = state_in[31:24] == 8'b11111110;
  assign _3099_ = state_in[31:24] == 8'b11111101;
  assign _3100_ = state_in[31:24] == 8'b11111100;
  assign _3101_ = state_in[31:24] == 8'b11111011;
  assign _3102_ = state_in[31:24] == 8'b11111010;
  assign _3103_ = state_in[31:24] == 8'b11111001;
  assign _3104_ = state_in[31:24] == 8'b11111000;
  assign _3105_ = state_in[31:24] == 8'b11110111;
  assign _3106_ = state_in[31:24] == 8'b11110110;
  assign _3107_ = state_in[31:24] == 8'b11110101;
  assign _3108_ = state_in[31:24] == 8'b11110100;
  assign _3109_ = state_in[31:24] == 8'b11110011;
  assign _3110_ = state_in[31:24] == 8'b11110010;
  assign _3111_ = state_in[31:24] == 8'b11110001;
  assign _3112_ = state_in[31:24] == 8'b11110000;
  assign _3113_ = state_in[31:24] == 8'b11101111;
  assign _3114_ = state_in[31:24] == 8'b11101110;
  assign _3115_ = state_in[31:24] == 8'b11101101;
  assign _3116_ = state_in[31:24] == 8'b11101100;
  assign _3117_ = state_in[31:24] == 8'b11101011;
  assign _3118_ = state_in[31:24] == 8'b11101010;
  assign _3119_ = state_in[31:24] == 8'b11101001;
  assign _3120_ = state_in[31:24] == 8'b11101000;
  assign _3121_ = state_in[31:24] == 8'b11100111;
  assign _3122_ = state_in[31:24] == 8'b11100110;
  assign _3123_ = state_in[31:24] == 8'b11100101;
  assign _3124_ = state_in[31:24] == 8'b11100100;
  assign _3125_ = state_in[31:24] == 8'b11100011;
  assign _3126_ = state_in[31:24] == 8'b11100010;
  assign _3127_ = state_in[31:24] == 8'b11100001;
  assign _3128_ = state_in[31:24] == 8'b11100000;
  assign _3129_ = state_in[31:24] == 8'b11011111;
  assign _3130_ = state_in[31:24] == 8'b11011110;
  assign _3131_ = state_in[31:24] == 8'b11011101;
  assign _3132_ = state_in[31:24] == 8'b11011100;
  assign _3133_ = state_in[31:24] == 8'b11011011;
  assign _3134_ = state_in[31:24] == 8'b11011010;
  assign _3135_ = state_in[31:24] == 8'b11011001;
  assign _3136_ = state_in[31:24] == 8'b11011000;
  assign _3137_ = state_in[31:24] == 8'b11010111;
  assign _3138_ = state_in[31:24] == 8'b11010110;
  assign _3139_ = state_in[31:24] == 8'b11010101;
  assign _3140_ = state_in[31:24] == 8'b11010100;
  assign _3141_ = state_in[31:24] == 8'b11010011;
  assign _3142_ = state_in[31:24] == 8'b11010010;
  assign _3143_ = state_in[31:24] == 8'b11010001;
  assign _3144_ = state_in[31:24] == 8'b11010000;
  assign _3145_ = state_in[31:24] == 8'b11001111;
  assign _3146_ = state_in[31:24] == 8'b11001110;
  assign _3147_ = state_in[31:24] == 8'b11001101;
  assign _3148_ = state_in[31:24] == 8'b11001100;
  assign _3149_ = state_in[31:24] == 8'b11001011;
  assign _3150_ = state_in[31:24] == 8'b11001010;
  assign _3151_ = state_in[31:24] == 8'b11001001;
  assign _3152_ = state_in[31:24] == 8'b11001000;
  assign _3153_ = state_in[31:24] == 8'b11000111;
  assign _3154_ = state_in[31:24] == 8'b11000110;
  assign _3155_ = state_in[31:24] == 8'b11000101;
  assign _3156_ = state_in[31:24] == 8'b11000100;
  assign _3157_ = state_in[31:24] == 8'b11000011;
  assign _3158_ = state_in[31:24] == 8'b11000010;
  assign _3159_ = state_in[31:24] == 8'b11000001;
  assign _3160_ = state_in[31:24] == 8'b11000000;
  assign _3161_ = state_in[31:24] == 8'b10111111;
  assign _3162_ = state_in[31:24] == 8'b10111110;
  assign _3163_ = state_in[31:24] == 8'b10111101;
  assign _3164_ = state_in[31:24] == 8'b10111100;
  assign _3165_ = state_in[31:24] == 8'b10111011;
  assign _3166_ = state_in[31:24] == 8'b10111010;
  assign _3167_ = state_in[31:24] == 8'b10111001;
  assign _3168_ = state_in[31:24] == 8'b10111000;
  assign _3169_ = state_in[31:24] == 8'b10110111;
  assign _3170_ = state_in[31:24] == 8'b10110110;
  assign _3171_ = state_in[31:24] == 8'b10110101;
  assign _3172_ = state_in[31:24] == 8'b10110100;
  assign _3173_ = state_in[31:24] == 8'b10110011;
  assign _3174_ = state_in[31:24] == 8'b10110010;
  assign _3175_ = state_in[31:24] == 8'b10110001;
  assign _3176_ = state_in[31:24] == 8'b10110000;
  assign _3177_ = state_in[31:24] == 8'b10101111;
  assign _3178_ = state_in[31:24] == 8'b10101110;
  assign _3179_ = state_in[31:24] == 8'b10101101;
  assign _3180_ = state_in[31:24] == 8'b10101100;
  assign _3181_ = state_in[31:24] == 8'b10101011;
  assign _3182_ = state_in[31:24] == 8'b10101010;
  assign _3183_ = state_in[31:24] == 8'b10101001;
  assign _3184_ = state_in[31:24] == 8'b10101000;
  assign _3185_ = state_in[31:24] == 8'b10100111;
  assign _3186_ = state_in[31:24] == 8'b10100110;
  assign _3187_ = state_in[31:24] == 8'b10100101;
  assign _3188_ = state_in[31:24] == 8'b10100100;
  assign _3189_ = state_in[31:24] == 8'b10100011;
  assign _3190_ = state_in[31:24] == 8'b10100010;
  assign _3191_ = state_in[31:24] == 8'b10100001;
  assign _3192_ = state_in[31:24] == 8'b10100000;
  assign _3193_ = state_in[31:24] == 8'b10011111;
  assign _3194_ = state_in[31:24] == 8'b10011110;
  assign _3195_ = state_in[31:24] == 8'b10011101;
  assign _3196_ = state_in[31:24] == 8'b10011100;
  assign _3197_ = state_in[31:24] == 8'b10011011;
  assign _3198_ = state_in[31:24] == 8'b10011010;
  assign _3199_ = state_in[31:24] == 8'b10011001;
  assign _3200_ = state_in[31:24] == 8'b10011000;
  assign _3201_ = state_in[31:24] == 8'b10010111;
  assign _3202_ = state_in[31:24] == 8'b10010110;
  assign _3203_ = state_in[31:24] == 8'b10010101;
  assign _3204_ = state_in[31:24] == 8'b10010100;
  assign _3205_ = state_in[31:24] == 8'b10010011;
  assign _3206_ = state_in[31:24] == 8'b10010010;
  assign _3207_ = state_in[31:24] == 8'b10010001;
  assign _3208_ = state_in[31:24] == 8'b10010000;
  assign _3209_ = state_in[31:24] == 8'b10001111;
  assign _3210_ = state_in[31:24] == 8'b10001110;
  assign _3211_ = state_in[31:24] == 8'b10001101;
  assign _3212_ = state_in[31:24] == 8'b10001100;
  assign _3213_ = state_in[31:24] == 8'b10001011;
  assign _3214_ = state_in[31:24] == 8'b10001010;
  assign _3215_ = state_in[31:24] == 8'b10001001;
  assign _3216_ = state_in[31:24] == 8'b10001000;
  assign _3217_ = state_in[31:24] == 8'b10000111;
  assign _3218_ = state_in[31:24] == 8'b10000110;
  assign _3219_ = state_in[31:24] == 8'b10000101;
  assign _3220_ = state_in[31:24] == 8'b10000100;
  assign _3221_ = state_in[31:24] == 8'b10000011;
  assign _3222_ = state_in[31:24] == 8'b10000010;
  assign _3223_ = state_in[31:24] == 8'b10000001;
  assign _3224_ = state_in[31:24] == 8'b10000000;
  assign _3225_ = state_in[31:24] == 7'b1111111;
  assign _3226_ = state_in[31:24] == 7'b1111110;
  assign _3227_ = state_in[31:24] == 7'b1111101;
  assign _3228_ = state_in[31:24] == 7'b1111100;
  assign _3229_ = state_in[31:24] == 7'b1111011;
  assign _3230_ = state_in[31:24] == 7'b1111010;
  assign _3231_ = state_in[31:24] == 7'b1111001;
  assign _3232_ = state_in[31:24] == 7'b1111000;
  assign _3233_ = state_in[31:24] == 7'b1110111;
  assign _3234_ = state_in[31:24] == 7'b1110110;
  assign _3235_ = state_in[31:24] == 7'b1110101;
  assign _3236_ = state_in[31:24] == 7'b1110100;
  assign _3237_ = state_in[31:24] == 7'b1110011;
  assign _3238_ = state_in[31:24] == 7'b1110010;
  assign _3239_ = state_in[31:24] == 7'b1110001;
  assign _3240_ = state_in[31:24] == 7'b1110000;
  assign _3241_ = state_in[31:24] == 7'b1101111;
  assign _3242_ = state_in[31:24] == 7'b1101110;
  assign _3243_ = state_in[31:24] == 7'b1101101;
  assign _3244_ = state_in[31:24] == 7'b1101100;
  assign _3245_ = state_in[31:24] == 7'b1101011;
  assign _3246_ = state_in[31:24] == 7'b1101010;
  assign _3247_ = state_in[31:24] == 7'b1101001;
  assign _3248_ = state_in[31:24] == 7'b1101000;
  assign _3249_ = state_in[31:24] == 7'b1100111;
  assign _3250_ = state_in[31:24] == 7'b1100110;
  assign _3251_ = state_in[31:24] == 7'b1100101;
  assign _3252_ = state_in[31:24] == 7'b1100100;
  assign _3253_ = state_in[31:24] == 7'b1100011;
  assign _3254_ = state_in[31:24] == 7'b1100010;
  assign _3255_ = state_in[31:24] == 7'b1100001;
  assign _3256_ = state_in[31:24] == 7'b1100000;
  assign _3257_ = state_in[31:24] == 7'b1011111;
  assign _3258_ = state_in[31:24] == 7'b1011110;
  assign _3259_ = state_in[31:24] == 7'b1011101;
  assign _3260_ = state_in[31:24] == 7'b1011100;
  assign _3261_ = state_in[31:24] == 7'b1011011;
  assign _3262_ = state_in[31:24] == 7'b1011010;
  assign _3263_ = state_in[31:24] == 7'b1011001;
  assign _3264_ = state_in[31:24] == 7'b1011000;
  assign _3265_ = state_in[31:24] == 7'b1010111;
  assign _3266_ = state_in[31:24] == 7'b1010110;
  assign _3267_ = state_in[31:24] == 7'b1010101;
  assign _3268_ = state_in[31:24] == 7'b1010100;
  assign _3269_ = state_in[31:24] == 7'b1010011;
  assign _3270_ = state_in[31:24] == 7'b1010010;
  assign _3271_ = state_in[31:24] == 7'b1010001;
  assign _3272_ = state_in[31:24] == 7'b1010000;
  assign _3273_ = state_in[31:24] == 7'b1001111;
  assign _3274_ = state_in[31:24] == 7'b1001110;
  assign _3275_ = state_in[31:24] == 7'b1001101;
  assign _3276_ = state_in[31:24] == 7'b1001100;
  assign _3277_ = state_in[31:24] == 7'b1001011;
  assign _3278_ = state_in[31:24] == 7'b1001010;
  assign _3279_ = state_in[31:24] == 7'b1001001;
  assign _3280_ = state_in[31:24] == 7'b1001000;
  assign _3281_ = state_in[31:24] == 7'b1000111;
  assign _3282_ = state_in[31:24] == 7'b1000110;
  assign _3283_ = state_in[31:24] == 7'b1000101;
  assign _3284_ = state_in[31:24] == 7'b1000100;
  assign _3285_ = state_in[31:24] == 7'b1000011;
  assign _3286_ = state_in[31:24] == 7'b1000010;
  assign _3287_ = state_in[31:24] == 7'b1000001;
  assign _3288_ = state_in[31:24] == 7'b1000000;
  assign _3289_ = state_in[31:24] == 6'b111111;
  assign _3290_ = state_in[31:24] == 6'b111110;
  assign _3291_ = state_in[31:24] == 6'b111101;
  assign _3292_ = state_in[31:24] == 6'b111100;
  assign _3293_ = state_in[31:24] == 6'b111011;
  assign _3294_ = state_in[31:24] == 6'b111010;
  assign _3295_ = state_in[31:24] == 6'b111001;
  assign _3296_ = state_in[31:24] == 6'b111000;
  assign _3297_ = state_in[31:24] == 6'b110111;
  assign _3298_ = state_in[31:24] == 6'b110110;
  assign _3299_ = state_in[31:24] == 6'b110101;
  assign _3300_ = state_in[31:24] == 6'b110100;
  assign _3301_ = state_in[31:24] == 6'b110011;
  assign _3302_ = state_in[31:24] == 6'b110010;
  assign _3303_ = state_in[31:24] == 6'b110001;
  assign _3304_ = state_in[31:24] == 6'b110000;
  assign _3305_ = state_in[31:24] == 6'b101111;
  assign _3306_ = state_in[31:24] == 6'b101110;
  assign _3307_ = state_in[31:24] == 6'b101101;
  assign _3308_ = state_in[31:24] == 6'b101100;
  assign _3309_ = state_in[31:24] == 6'b101011;
  assign _3310_ = state_in[31:24] == 6'b101010;
  assign _3311_ = state_in[31:24] == 6'b101001;
  assign _3312_ = state_in[31:24] == 6'b101000;
  assign _3313_ = state_in[31:24] == 6'b100111;
  assign _3314_ = state_in[31:24] == 6'b100110;
  assign _3315_ = state_in[31:24] == 6'b100101;
  assign _3316_ = state_in[31:24] == 6'b100100;
  assign _3317_ = state_in[31:24] == 6'b100011;
  assign _3318_ = state_in[31:24] == 6'b100010;
  assign _3319_ = state_in[31:24] == 6'b100001;
  assign _3320_ = state_in[31:24] == 6'b100000;
  assign _3321_ = state_in[31:24] == 5'b11111;
  assign _3322_ = state_in[31:24] == 5'b11110;
  assign _3323_ = state_in[31:24] == 5'b11101;
  assign _3324_ = state_in[31:24] == 5'b11100;
  assign _3325_ = state_in[31:24] == 5'b11011;
  assign _3326_ = state_in[31:24] == 5'b11010;
  assign _3327_ = state_in[31:24] == 5'b11001;
  assign _3328_ = state_in[31:24] == 5'b11000;
  assign _3329_ = state_in[31:24] == 5'b10111;
  assign _3330_ = state_in[31:24] == 5'b10110;
  assign _3331_ = state_in[31:24] == 5'b10101;
  assign _3332_ = state_in[31:24] == 5'b10100;
  assign _3333_ = state_in[31:24] == 5'b10011;
  assign _3334_ = state_in[31:24] == 5'b10010;
  assign _3335_ = state_in[31:24] == 5'b10001;
  assign _3336_ = state_in[31:24] == 5'b10000;
  assign _3337_ = state_in[31:24] == 4'b1111;
  assign _3338_ = state_in[31:24] == 4'b1110;
  assign _3339_ = state_in[31:24] == 4'b1101;
  assign _3340_ = state_in[31:24] == 4'b1100;
  assign _3341_ = state_in[31:24] == 4'b1011;
  assign _3342_ = state_in[31:24] == 4'b1010;
  assign _3343_ = state_in[31:24] == 4'b1001;
  assign _3344_ = state_in[31:24] == 4'b1000;
  assign _3345_ = state_in[31:24] == 3'b111;
  assign _3346_ = state_in[31:24] == 3'b110;
  assign _3347_ = state_in[31:24] == 3'b101;
  assign _3348_ = state_in[31:24] == 3'b100;
  assign _3349_ = state_in[31:24] == 2'b11;
  assign _3350_ = state_in[31:24] == 2'b10;
  assign _3351_ = state_in[31:24] == 1'b1;
  assign _3352_ = ! state_in[31:24];
  always @(posedge clk)
      \t3.t0.s4.out <= _3353_;
  logic [255:0] fangyuan26;
  assign fangyuan26 = { _3352_, _3351_, _3350_, _3349_, _3348_, _3347_, _3346_, _3345_, _3344_, _3343_, _3342_, _3341_, _3340_, _3339_, _3338_, _3337_, _3336_, _3335_, _3334_, _3333_, _3332_, _3331_, _3330_, _3329_, _3328_, _3327_, _3326_, _3325_, _3324_, _3323_, _3322_, _3321_, _3320_, _3319_, _3318_, _3317_, _3316_, _3315_, _3314_, _3313_, _3312_, _3311_, _3310_, _3309_, _3308_, _3307_, _3306_, _3305_, _3304_, _3303_, _3302_, _3301_, _3300_, _3299_, _3298_, _3297_, _3296_, _3295_, _3294_, _3293_, _3292_, _3291_, _3290_, _3289_, _3288_, _3287_, _3286_, _3285_, _3284_, _3283_, _3282_, _3281_, _3280_, _3279_, _3278_, _3277_, _3276_, _3275_, _3274_, _3273_, _3272_, _3271_, _3270_, _3269_, _3268_, _3267_, _3266_, _3265_, _3264_, _3263_, _3262_, _3261_, _3260_, _3259_, _3258_, _3257_, _3256_, _3255_, _3254_, _3253_, _3252_, _3251_, _3250_, _3249_, _3248_, _3247_, _3246_, _3245_, _3244_, _3243_, _3242_, _3241_, _3240_, _3239_, _3238_, _3237_, _3236_, _3235_, _3234_, _3233_, _3232_, _3231_, _3230_, _3229_, _3228_, _3227_, _3226_, _3225_, _3224_, _3223_, _3222_, _3221_, _3220_, _3219_, _3218_, _3217_, _3216_, _3215_, _3214_, _3213_, _3212_, _3211_, _3210_, _3209_, _3208_, _3207_, _3206_, _3205_, _3204_, _3203_, _3202_, _3201_, _3200_, _3199_, _3198_, _3197_, _3196_, _3195_, _3194_, _3193_, _3192_, _3191_, _3190_, _3189_, _3188_, _3187_, _3186_, _3185_, _3184_, _3183_, _3182_, _3181_, _3180_, _3179_, _3178_, _3177_, _3176_, _3175_, _3174_, _3173_, _3172_, _3171_, _3170_, _3169_, _3168_, _3167_, _3166_, _3165_, _3164_, _3163_, _3162_, _3161_, _3160_, _3159_, _3158_, _3157_, _3156_, _3155_, _3154_, _3153_, _3152_, _3151_, _3150_, _3149_, _3148_, _3147_, _3146_, _3145_, _3144_, _3143_, _3142_, _3141_, _3140_, _3139_, _3138_, _3137_, _3136_, _3135_, _3134_, _3133_, _3132_, _3131_, _3130_, _3129_, _3128_, _3127_, _3126_, _3125_, _3124_, _3123_, _3122_, _3121_, _3120_, _3119_, _3118_, _3117_, _3116_, _3115_, _3114_, _3113_, _3112_, _3111_, _3110_, _3109_, _3108_, _3107_, _3106_, _3105_, _3104_, _3103_, _3102_, _3101_, _3100_, _3099_, _3098_, _3097_ };

  always @(\t3.t0.s4.out or fangyuan26) begin
    casez (fangyuan26)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3353_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3353_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3353_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3353_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3353_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3353_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3353_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3353_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3353_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3353_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3353_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3353_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3353_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3353_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3353_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3353_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3353_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3353_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3353_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3353_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3353_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3353_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3353_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3353_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3353_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3353_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3353_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3353_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3353_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3353_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3353_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3353_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3353_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3353_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3353_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3353_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3353_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3353_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3353_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3353_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3353_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3353_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3353_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3353_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3353_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3353_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3353_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3353_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3353_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3353_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3353_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3353_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3353_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3353_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3353_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3353_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3353_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3353_ = 8'b11000110 ;
      default:
        _3353_ = \t3.t0.s4.out ;
    endcase
  end
  assign p31[31:24] = \t3.t1.s0.out ^ \t3.t1.s4.out ;
  always @(posedge clk)
      \t3.t1.s0.out <= _3354_;
  logic [255:0] fangyuan27;
  assign fangyuan27 = { _3610_, _3609_, _3608_, _3607_, _3606_, _3605_, _3604_, _3603_, _3602_, _3601_, _3600_, _3599_, _3598_, _3597_, _3596_, _3595_, _3594_, _3593_, _3592_, _3591_, _3590_, _3589_, _3588_, _3587_, _3586_, _3585_, _3584_, _3583_, _3582_, _3581_, _3580_, _3579_, _3578_, _3577_, _3576_, _3575_, _3574_, _3573_, _3572_, _3571_, _3570_, _3569_, _3568_, _3567_, _3566_, _3565_, _3564_, _3563_, _3562_, _3561_, _3560_, _3559_, _3558_, _3557_, _3556_, _3555_, _3554_, _3553_, _3552_, _3551_, _3550_, _3549_, _3548_, _3547_, _3546_, _3545_, _3544_, _3543_, _3542_, _3541_, _3540_, _3539_, _3538_, _3537_, _3536_, _3535_, _3534_, _3533_, _3532_, _3531_, _3530_, _3529_, _3528_, _3527_, _3526_, _3525_, _3524_, _3523_, _3522_, _3521_, _3520_, _3519_, _3518_, _3517_, _3516_, _3515_, _3514_, _3513_, _3512_, _3511_, _3510_, _3509_, _3508_, _3507_, _3506_, _3505_, _3504_, _3503_, _3502_, _3501_, _3500_, _3499_, _3498_, _3497_, _3496_, _3495_, _3494_, _3493_, _3492_, _3491_, _3490_, _3489_, _3488_, _3487_, _3486_, _3485_, _3484_, _3483_, _3482_, _3481_, _3480_, _3479_, _3478_, _3477_, _3476_, _3475_, _3474_, _3473_, _3472_, _3471_, _3470_, _3469_, _3468_, _3467_, _3466_, _3465_, _3464_, _3463_, _3462_, _3461_, _3460_, _3459_, _3458_, _3457_, _3456_, _3455_, _3454_, _3453_, _3452_, _3451_, _3450_, _3449_, _3448_, _3447_, _3446_, _3445_, _3444_, _3443_, _3442_, _3441_, _3440_, _3439_, _3438_, _3437_, _3436_, _3435_, _3434_, _3433_, _3432_, _3431_, _3430_, _3429_, _3428_, _3427_, _3426_, _3425_, _3424_, _3423_, _3422_, _3421_, _3420_, _3419_, _3418_, _3417_, _3416_, _3415_, _3414_, _3413_, _3412_, _3411_, _3410_, _3409_, _3408_, _3407_, _3406_, _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_, _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_ };

  always @(\t3.t1.s0.out or fangyuan27) begin
    casez (fangyuan27)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3354_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3354_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3354_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3354_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3354_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3354_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3354_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3354_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3354_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3354_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3354_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3354_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3354_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3354_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3354_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3354_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3354_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3354_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3354_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3354_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3354_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3354_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3354_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3354_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3354_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3354_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3354_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3354_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3354_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3354_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3354_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3354_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3354_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3354_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3354_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3354_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3354_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3354_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3354_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3354_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3354_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3354_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3354_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3354_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3354_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3354_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3354_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3354_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3354_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3354_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3354_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3354_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3354_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3354_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3354_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3354_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3354_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3354_ = 8'b01100011 ;
      default:
        _3354_ = \t3.t1.s0.out ;
    endcase
  end
  assign _3355_ = state_in[23:16] == 8'b11111111;
  assign _3356_ = state_in[23:16] == 8'b11111110;
  assign _3357_ = state_in[23:16] == 8'b11111101;
  assign _3358_ = state_in[23:16] == 8'b11111100;
  assign _3359_ = state_in[23:16] == 8'b11111011;
  assign _3360_ = state_in[23:16] == 8'b11111010;
  assign _3361_ = state_in[23:16] == 8'b11111001;
  assign _3362_ = state_in[23:16] == 8'b11111000;
  assign _3363_ = state_in[23:16] == 8'b11110111;
  assign _3364_ = state_in[23:16] == 8'b11110110;
  assign _3365_ = state_in[23:16] == 8'b11110101;
  assign _3366_ = state_in[23:16] == 8'b11110100;
  assign _3367_ = state_in[23:16] == 8'b11110011;
  assign _3368_ = state_in[23:16] == 8'b11110010;
  assign _3369_ = state_in[23:16] == 8'b11110001;
  assign _3370_ = state_in[23:16] == 8'b11110000;
  assign _3371_ = state_in[23:16] == 8'b11101111;
  assign _3372_ = state_in[23:16] == 8'b11101110;
  assign _3373_ = state_in[23:16] == 8'b11101101;
  assign _3374_ = state_in[23:16] == 8'b11101100;
  assign _3375_ = state_in[23:16] == 8'b11101011;
  assign _3376_ = state_in[23:16] == 8'b11101010;
  assign _3377_ = state_in[23:16] == 8'b11101001;
  assign _3378_ = state_in[23:16] == 8'b11101000;
  assign _3379_ = state_in[23:16] == 8'b11100111;
  assign _3380_ = state_in[23:16] == 8'b11100110;
  assign _3381_ = state_in[23:16] == 8'b11100101;
  assign _3382_ = state_in[23:16] == 8'b11100100;
  assign _3383_ = state_in[23:16] == 8'b11100011;
  assign _3384_ = state_in[23:16] == 8'b11100010;
  assign _3385_ = state_in[23:16] == 8'b11100001;
  assign _3386_ = state_in[23:16] == 8'b11100000;
  assign _3387_ = state_in[23:16] == 8'b11011111;
  assign _3388_ = state_in[23:16] == 8'b11011110;
  assign _3389_ = state_in[23:16] == 8'b11011101;
  assign _3390_ = state_in[23:16] == 8'b11011100;
  assign _3391_ = state_in[23:16] == 8'b11011011;
  assign _3392_ = state_in[23:16] == 8'b11011010;
  assign _3393_ = state_in[23:16] == 8'b11011001;
  assign _3394_ = state_in[23:16] == 8'b11011000;
  assign _3395_ = state_in[23:16] == 8'b11010111;
  assign _3396_ = state_in[23:16] == 8'b11010110;
  assign _3397_ = state_in[23:16] == 8'b11010101;
  assign _3398_ = state_in[23:16] == 8'b11010100;
  assign _3399_ = state_in[23:16] == 8'b11010011;
  assign _3400_ = state_in[23:16] == 8'b11010010;
  assign _3401_ = state_in[23:16] == 8'b11010001;
  assign _3402_ = state_in[23:16] == 8'b11010000;
  assign _3403_ = state_in[23:16] == 8'b11001111;
  assign _3404_ = state_in[23:16] == 8'b11001110;
  assign _3405_ = state_in[23:16] == 8'b11001101;
  assign _3406_ = state_in[23:16] == 8'b11001100;
  assign _3407_ = state_in[23:16] == 8'b11001011;
  assign _3408_ = state_in[23:16] == 8'b11001010;
  assign _3409_ = state_in[23:16] == 8'b11001001;
  assign _3410_ = state_in[23:16] == 8'b11001000;
  assign _3411_ = state_in[23:16] == 8'b11000111;
  assign _3412_ = state_in[23:16] == 8'b11000110;
  assign _3413_ = state_in[23:16] == 8'b11000101;
  assign _3414_ = state_in[23:16] == 8'b11000100;
  assign _3415_ = state_in[23:16] == 8'b11000011;
  assign _3416_ = state_in[23:16] == 8'b11000010;
  assign _3417_ = state_in[23:16] == 8'b11000001;
  assign _3418_ = state_in[23:16] == 8'b11000000;
  assign _3419_ = state_in[23:16] == 8'b10111111;
  assign _3420_ = state_in[23:16] == 8'b10111110;
  assign _3421_ = state_in[23:16] == 8'b10111101;
  assign _3422_ = state_in[23:16] == 8'b10111100;
  assign _3423_ = state_in[23:16] == 8'b10111011;
  assign _3424_ = state_in[23:16] == 8'b10111010;
  assign _3425_ = state_in[23:16] == 8'b10111001;
  assign _3426_ = state_in[23:16] == 8'b10111000;
  assign _3427_ = state_in[23:16] == 8'b10110111;
  assign _3428_ = state_in[23:16] == 8'b10110110;
  assign _3429_ = state_in[23:16] == 8'b10110101;
  assign _3430_ = state_in[23:16] == 8'b10110100;
  assign _3431_ = state_in[23:16] == 8'b10110011;
  assign _3432_ = state_in[23:16] == 8'b10110010;
  assign _3433_ = state_in[23:16] == 8'b10110001;
  assign _3434_ = state_in[23:16] == 8'b10110000;
  assign _3435_ = state_in[23:16] == 8'b10101111;
  assign _3436_ = state_in[23:16] == 8'b10101110;
  assign _3437_ = state_in[23:16] == 8'b10101101;
  assign _3438_ = state_in[23:16] == 8'b10101100;
  assign _3439_ = state_in[23:16] == 8'b10101011;
  assign _3440_ = state_in[23:16] == 8'b10101010;
  assign _3441_ = state_in[23:16] == 8'b10101001;
  assign _3442_ = state_in[23:16] == 8'b10101000;
  assign _3443_ = state_in[23:16] == 8'b10100111;
  assign _3444_ = state_in[23:16] == 8'b10100110;
  assign _3445_ = state_in[23:16] == 8'b10100101;
  assign _3446_ = state_in[23:16] == 8'b10100100;
  assign _3447_ = state_in[23:16] == 8'b10100011;
  assign _3448_ = state_in[23:16] == 8'b10100010;
  assign _3449_ = state_in[23:16] == 8'b10100001;
  assign _3450_ = state_in[23:16] == 8'b10100000;
  assign _3451_ = state_in[23:16] == 8'b10011111;
  assign _3452_ = state_in[23:16] == 8'b10011110;
  assign _3453_ = state_in[23:16] == 8'b10011101;
  assign _3454_ = state_in[23:16] == 8'b10011100;
  assign _3455_ = state_in[23:16] == 8'b10011011;
  assign _3456_ = state_in[23:16] == 8'b10011010;
  assign _3457_ = state_in[23:16] == 8'b10011001;
  assign _3458_ = state_in[23:16] == 8'b10011000;
  assign _3459_ = state_in[23:16] == 8'b10010111;
  assign _3460_ = state_in[23:16] == 8'b10010110;
  assign _3461_ = state_in[23:16] == 8'b10010101;
  assign _3462_ = state_in[23:16] == 8'b10010100;
  assign _3463_ = state_in[23:16] == 8'b10010011;
  assign _3464_ = state_in[23:16] == 8'b10010010;
  assign _3465_ = state_in[23:16] == 8'b10010001;
  assign _3466_ = state_in[23:16] == 8'b10010000;
  assign _3467_ = state_in[23:16] == 8'b10001111;
  assign _3468_ = state_in[23:16] == 8'b10001110;
  assign _3469_ = state_in[23:16] == 8'b10001101;
  assign _3470_ = state_in[23:16] == 8'b10001100;
  assign _3471_ = state_in[23:16] == 8'b10001011;
  assign _3472_ = state_in[23:16] == 8'b10001010;
  assign _3473_ = state_in[23:16] == 8'b10001001;
  assign _3474_ = state_in[23:16] == 8'b10001000;
  assign _3475_ = state_in[23:16] == 8'b10000111;
  assign _3476_ = state_in[23:16] == 8'b10000110;
  assign _3477_ = state_in[23:16] == 8'b10000101;
  assign _3478_ = state_in[23:16] == 8'b10000100;
  assign _3479_ = state_in[23:16] == 8'b10000011;
  assign _3480_ = state_in[23:16] == 8'b10000010;
  assign _3481_ = state_in[23:16] == 8'b10000001;
  assign _3482_ = state_in[23:16] == 8'b10000000;
  assign _3483_ = state_in[23:16] == 7'b1111111;
  assign _3484_ = state_in[23:16] == 7'b1111110;
  assign _3485_ = state_in[23:16] == 7'b1111101;
  assign _3486_ = state_in[23:16] == 7'b1111100;
  assign _3487_ = state_in[23:16] == 7'b1111011;
  assign _3488_ = state_in[23:16] == 7'b1111010;
  assign _3489_ = state_in[23:16] == 7'b1111001;
  assign _3490_ = state_in[23:16] == 7'b1111000;
  assign _3491_ = state_in[23:16] == 7'b1110111;
  assign _3492_ = state_in[23:16] == 7'b1110110;
  assign _3493_ = state_in[23:16] == 7'b1110101;
  assign _3494_ = state_in[23:16] == 7'b1110100;
  assign _3495_ = state_in[23:16] == 7'b1110011;
  assign _3496_ = state_in[23:16] == 7'b1110010;
  assign _3497_ = state_in[23:16] == 7'b1110001;
  assign _3498_ = state_in[23:16] == 7'b1110000;
  assign _3499_ = state_in[23:16] == 7'b1101111;
  assign _3500_ = state_in[23:16] == 7'b1101110;
  assign _3501_ = state_in[23:16] == 7'b1101101;
  assign _3502_ = state_in[23:16] == 7'b1101100;
  assign _3503_ = state_in[23:16] == 7'b1101011;
  assign _3504_ = state_in[23:16] == 7'b1101010;
  assign _3505_ = state_in[23:16] == 7'b1101001;
  assign _3506_ = state_in[23:16] == 7'b1101000;
  assign _3507_ = state_in[23:16] == 7'b1100111;
  assign _3508_ = state_in[23:16] == 7'b1100110;
  assign _3509_ = state_in[23:16] == 7'b1100101;
  assign _3510_ = state_in[23:16] == 7'b1100100;
  assign _3511_ = state_in[23:16] == 7'b1100011;
  assign _3512_ = state_in[23:16] == 7'b1100010;
  assign _3513_ = state_in[23:16] == 7'b1100001;
  assign _3514_ = state_in[23:16] == 7'b1100000;
  assign _3515_ = state_in[23:16] == 7'b1011111;
  assign _3516_ = state_in[23:16] == 7'b1011110;
  assign _3517_ = state_in[23:16] == 7'b1011101;
  assign _3518_ = state_in[23:16] == 7'b1011100;
  assign _3519_ = state_in[23:16] == 7'b1011011;
  assign _3520_ = state_in[23:16] == 7'b1011010;
  assign _3521_ = state_in[23:16] == 7'b1011001;
  assign _3522_ = state_in[23:16] == 7'b1011000;
  assign _3523_ = state_in[23:16] == 7'b1010111;
  assign _3524_ = state_in[23:16] == 7'b1010110;
  assign _3525_ = state_in[23:16] == 7'b1010101;
  assign _3526_ = state_in[23:16] == 7'b1010100;
  assign _3527_ = state_in[23:16] == 7'b1010011;
  assign _3528_ = state_in[23:16] == 7'b1010010;
  assign _3529_ = state_in[23:16] == 7'b1010001;
  assign _3530_ = state_in[23:16] == 7'b1010000;
  assign _3531_ = state_in[23:16] == 7'b1001111;
  assign _3532_ = state_in[23:16] == 7'b1001110;
  assign _3533_ = state_in[23:16] == 7'b1001101;
  assign _3534_ = state_in[23:16] == 7'b1001100;
  assign _3535_ = state_in[23:16] == 7'b1001011;
  assign _3536_ = state_in[23:16] == 7'b1001010;
  assign _3537_ = state_in[23:16] == 7'b1001001;
  assign _3538_ = state_in[23:16] == 7'b1001000;
  assign _3539_ = state_in[23:16] == 7'b1000111;
  assign _3540_ = state_in[23:16] == 7'b1000110;
  assign _3541_ = state_in[23:16] == 7'b1000101;
  assign _3542_ = state_in[23:16] == 7'b1000100;
  assign _3543_ = state_in[23:16] == 7'b1000011;
  assign _3544_ = state_in[23:16] == 7'b1000010;
  assign _3545_ = state_in[23:16] == 7'b1000001;
  assign _3546_ = state_in[23:16] == 7'b1000000;
  assign _3547_ = state_in[23:16] == 6'b111111;
  assign _3548_ = state_in[23:16] == 6'b111110;
  assign _3549_ = state_in[23:16] == 6'b111101;
  assign _3550_ = state_in[23:16] == 6'b111100;
  assign _3551_ = state_in[23:16] == 6'b111011;
  assign _3552_ = state_in[23:16] == 6'b111010;
  assign _3553_ = state_in[23:16] == 6'b111001;
  assign _3554_ = state_in[23:16] == 6'b111000;
  assign _3555_ = state_in[23:16] == 6'b110111;
  assign _3556_ = state_in[23:16] == 6'b110110;
  assign _3557_ = state_in[23:16] == 6'b110101;
  assign _3558_ = state_in[23:16] == 6'b110100;
  assign _3559_ = state_in[23:16] == 6'b110011;
  assign _3560_ = state_in[23:16] == 6'b110010;
  assign _3561_ = state_in[23:16] == 6'b110001;
  assign _3562_ = state_in[23:16] == 6'b110000;
  assign _3563_ = state_in[23:16] == 6'b101111;
  assign _3564_ = state_in[23:16] == 6'b101110;
  assign _3565_ = state_in[23:16] == 6'b101101;
  assign _3566_ = state_in[23:16] == 6'b101100;
  assign _3567_ = state_in[23:16] == 6'b101011;
  assign _3568_ = state_in[23:16] == 6'b101010;
  assign _3569_ = state_in[23:16] == 6'b101001;
  assign _3570_ = state_in[23:16] == 6'b101000;
  assign _3571_ = state_in[23:16] == 6'b100111;
  assign _3572_ = state_in[23:16] == 6'b100110;
  assign _3573_ = state_in[23:16] == 6'b100101;
  assign _3574_ = state_in[23:16] == 6'b100100;
  assign _3575_ = state_in[23:16] == 6'b100011;
  assign _3576_ = state_in[23:16] == 6'b100010;
  assign _3577_ = state_in[23:16] == 6'b100001;
  assign _3578_ = state_in[23:16] == 6'b100000;
  assign _3579_ = state_in[23:16] == 5'b11111;
  assign _3580_ = state_in[23:16] == 5'b11110;
  assign _3581_ = state_in[23:16] == 5'b11101;
  assign _3582_ = state_in[23:16] == 5'b11100;
  assign _3583_ = state_in[23:16] == 5'b11011;
  assign _3584_ = state_in[23:16] == 5'b11010;
  assign _3585_ = state_in[23:16] == 5'b11001;
  assign _3586_ = state_in[23:16] == 5'b11000;
  assign _3587_ = state_in[23:16] == 5'b10111;
  assign _3588_ = state_in[23:16] == 5'b10110;
  assign _3589_ = state_in[23:16] == 5'b10101;
  assign _3590_ = state_in[23:16] == 5'b10100;
  assign _3591_ = state_in[23:16] == 5'b10011;
  assign _3592_ = state_in[23:16] == 5'b10010;
  assign _3593_ = state_in[23:16] == 5'b10001;
  assign _3594_ = state_in[23:16] == 5'b10000;
  assign _3595_ = state_in[23:16] == 4'b1111;
  assign _3596_ = state_in[23:16] == 4'b1110;
  assign _3597_ = state_in[23:16] == 4'b1101;
  assign _3598_ = state_in[23:16] == 4'b1100;
  assign _3599_ = state_in[23:16] == 4'b1011;
  assign _3600_ = state_in[23:16] == 4'b1010;
  assign _3601_ = state_in[23:16] == 4'b1001;
  assign _3602_ = state_in[23:16] == 4'b1000;
  assign _3603_ = state_in[23:16] == 3'b111;
  assign _3604_ = state_in[23:16] == 3'b110;
  assign _3605_ = state_in[23:16] == 3'b101;
  assign _3606_ = state_in[23:16] == 3'b100;
  assign _3607_ = state_in[23:16] == 2'b11;
  assign _3608_ = state_in[23:16] == 2'b10;
  assign _3609_ = state_in[23:16] == 1'b1;
  assign _3610_ = ! state_in[23:16];
  always @(posedge clk)
      \t3.t1.s4.out <= _3611_;
  logic [255:0] fangyuan28;
  assign fangyuan28 = { _3610_, _3609_, _3608_, _3607_, _3606_, _3605_, _3604_, _3603_, _3602_, _3601_, _3600_, _3599_, _3598_, _3597_, _3596_, _3595_, _3594_, _3593_, _3592_, _3591_, _3590_, _3589_, _3588_, _3587_, _3586_, _3585_, _3584_, _3583_, _3582_, _3581_, _3580_, _3579_, _3578_, _3577_, _3576_, _3575_, _3574_, _3573_, _3572_, _3571_, _3570_, _3569_, _3568_, _3567_, _3566_, _3565_, _3564_, _3563_, _3562_, _3561_, _3560_, _3559_, _3558_, _3557_, _3556_, _3555_, _3554_, _3553_, _3552_, _3551_, _3550_, _3549_, _3548_, _3547_, _3546_, _3545_, _3544_, _3543_, _3542_, _3541_, _3540_, _3539_, _3538_, _3537_, _3536_, _3535_, _3534_, _3533_, _3532_, _3531_, _3530_, _3529_, _3528_, _3527_, _3526_, _3525_, _3524_, _3523_, _3522_, _3521_, _3520_, _3519_, _3518_, _3517_, _3516_, _3515_, _3514_, _3513_, _3512_, _3511_, _3510_, _3509_, _3508_, _3507_, _3506_, _3505_, _3504_, _3503_, _3502_, _3501_, _3500_, _3499_, _3498_, _3497_, _3496_, _3495_, _3494_, _3493_, _3492_, _3491_, _3490_, _3489_, _3488_, _3487_, _3486_, _3485_, _3484_, _3483_, _3482_, _3481_, _3480_, _3479_, _3478_, _3477_, _3476_, _3475_, _3474_, _3473_, _3472_, _3471_, _3470_, _3469_, _3468_, _3467_, _3466_, _3465_, _3464_, _3463_, _3462_, _3461_, _3460_, _3459_, _3458_, _3457_, _3456_, _3455_, _3454_, _3453_, _3452_, _3451_, _3450_, _3449_, _3448_, _3447_, _3446_, _3445_, _3444_, _3443_, _3442_, _3441_, _3440_, _3439_, _3438_, _3437_, _3436_, _3435_, _3434_, _3433_, _3432_, _3431_, _3430_, _3429_, _3428_, _3427_, _3426_, _3425_, _3424_, _3423_, _3422_, _3421_, _3420_, _3419_, _3418_, _3417_, _3416_, _3415_, _3414_, _3413_, _3412_, _3411_, _3410_, _3409_, _3408_, _3407_, _3406_, _3405_, _3404_, _3403_, _3402_, _3401_, _3400_, _3399_, _3398_, _3397_, _3396_, _3395_, _3394_, _3393_, _3392_, _3391_, _3390_, _3389_, _3388_, _3387_, _3386_, _3385_, _3384_, _3383_, _3382_, _3381_, _3380_, _3379_, _3378_, _3377_, _3376_, _3375_, _3374_, _3373_, _3372_, _3371_, _3370_, _3369_, _3368_, _3367_, _3366_, _3365_, _3364_, _3363_, _3362_, _3361_, _3360_, _3359_, _3358_, _3357_, _3356_, _3355_ };

  always @(\t3.t1.s4.out or fangyuan28) begin
    casez (fangyuan28)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3611_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3611_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3611_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3611_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3611_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3611_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3611_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3611_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3611_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3611_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3611_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3611_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3611_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3611_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3611_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3611_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3611_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3611_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3611_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3611_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3611_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3611_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3611_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3611_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3611_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3611_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3611_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3611_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3611_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3611_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3611_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3611_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3611_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3611_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3611_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3611_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3611_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3611_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3611_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3611_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3611_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3611_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3611_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3611_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3611_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3611_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3611_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3611_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3611_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3611_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3611_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3611_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3611_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3611_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3611_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3611_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3611_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3611_ = 8'b11000110 ;
      default:
        _3611_ = \t3.t1.s4.out ;
    endcase
  end
  assign p32[23:16] = \t3.t2.s0.out ^ \t3.t2.s4.out ;
  always @(posedge clk)
      \t3.t2.s0.out <= _3612_;
  logic [255:0] fangyuan29;
  assign fangyuan29 = { _3868_, _3867_, _3866_, _3865_, _3864_, _3863_, _3862_, _3861_, _3860_, _3859_, _3858_, _3857_, _3856_, _3855_, _3854_, _3853_, _3852_, _3851_, _3850_, _3849_, _3848_, _3847_, _3846_, _3845_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3838_, _3837_, _3836_, _3835_, _3834_, _3833_, _3832_, _3831_, _3830_, _3829_, _3828_, _3827_, _3826_, _3825_, _3824_, _3823_, _3822_, _3821_, _3820_, _3819_, _3818_, _3817_, _3816_, _3815_, _3814_, _3813_, _3812_, _3811_, _3810_, _3809_, _3808_, _3807_, _3806_, _3805_, _3804_, _3803_, _3802_, _3801_, _3800_, _3799_, _3798_, _3797_, _3796_, _3795_, _3794_, _3793_, _3792_, _3791_, _3790_, _3789_, _3788_, _3787_, _3786_, _3785_, _3784_, _3783_, _3782_, _3781_, _3780_, _3779_, _3778_, _3777_, _3776_, _3775_, _3774_, _3773_, _3772_, _3771_, _3770_, _3769_, _3768_, _3767_, _3766_, _3765_, _3764_, _3763_, _3762_, _3761_, _3760_, _3759_, _3758_, _3757_, _3756_, _3755_, _3754_, _3753_, _3752_, _3751_, _3750_, _3749_, _3748_, _3747_, _3746_, _3745_, _3744_, _3743_, _3742_, _3741_, _3740_, _3739_, _3738_, _3737_, _3736_, _3735_, _3734_, _3733_, _3732_, _3731_, _3730_, _3729_, _3728_, _3727_, _3726_, _3725_, _3724_, _3723_, _3722_, _3721_, _3720_, _3719_, _3718_, _3717_, _3716_, _3715_, _3714_, _3713_, _3712_, _3711_, _3710_, _3709_, _3708_, _3707_, _3706_, _3705_, _3704_, _3703_, _3702_, _3701_, _3700_, _3699_, _3698_, _3697_, _3696_, _3695_, _3694_, _3693_, _3692_, _3691_, _3690_, _3689_, _3688_, _3687_, _3686_, _3685_, _3684_, _3683_, _3682_, _3681_, _3680_, _3679_, _3678_, _3677_, _3676_, _3675_, _3674_, _3673_, _3672_, _3671_, _3670_, _3669_, _3668_, _3667_, _3666_, _3665_, _3664_, _3663_, _3662_, _3661_, _3660_, _3659_, _3658_, _3657_, _3656_, _3655_, _3654_, _3653_, _3652_, _3651_, _3650_, _3649_, _3648_, _3647_, _3646_, _3645_, _3644_, _3643_, _3642_, _3641_, _3640_, _3639_, _3638_, _3637_, _3636_, _3635_, _3634_, _3633_, _3632_, _3631_, _3630_, _3629_, _3628_, _3627_, _3626_, _3625_, _3624_, _3623_, _3622_, _3621_, _3620_, _3619_, _3618_, _3617_, _3616_, _3615_, _3614_, _3613_ };

  always @(\t3.t2.s0.out or fangyuan29) begin
    casez (fangyuan29)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3612_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3612_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3612_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3612_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3612_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3612_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3612_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3612_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3612_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3612_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3612_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3612_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3612_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3612_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3612_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3612_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3612_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3612_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3612_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3612_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3612_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3612_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3612_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3612_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3612_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3612_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3612_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3612_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3612_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3612_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3612_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3612_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3612_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3612_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3612_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3612_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3612_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3612_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3612_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3612_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3612_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3612_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3612_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3612_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3612_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3612_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3612_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3612_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3612_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3612_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3612_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3612_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3612_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3612_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3612_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3612_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3612_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3612_ = 8'b01100011 ;
      default:
        _3612_ = \t3.t2.s0.out ;
    endcase
  end
  assign _3613_ = state_in[15:8] == 8'b11111111;
  assign _3614_ = state_in[15:8] == 8'b11111110;
  assign _3615_ = state_in[15:8] == 8'b11111101;
  assign _3616_ = state_in[15:8] == 8'b11111100;
  assign _3617_ = state_in[15:8] == 8'b11111011;
  assign _3618_ = state_in[15:8] == 8'b11111010;
  assign _3619_ = state_in[15:8] == 8'b11111001;
  assign _3620_ = state_in[15:8] == 8'b11111000;
  assign _3621_ = state_in[15:8] == 8'b11110111;
  assign _3622_ = state_in[15:8] == 8'b11110110;
  assign _3623_ = state_in[15:8] == 8'b11110101;
  assign _3624_ = state_in[15:8] == 8'b11110100;
  assign _3625_ = state_in[15:8] == 8'b11110011;
  assign _3626_ = state_in[15:8] == 8'b11110010;
  assign _3627_ = state_in[15:8] == 8'b11110001;
  assign _3628_ = state_in[15:8] == 8'b11110000;
  assign _3629_ = state_in[15:8] == 8'b11101111;
  assign _3630_ = state_in[15:8] == 8'b11101110;
  assign _3631_ = state_in[15:8] == 8'b11101101;
  assign _3632_ = state_in[15:8] == 8'b11101100;
  assign _3633_ = state_in[15:8] == 8'b11101011;
  assign _3634_ = state_in[15:8] == 8'b11101010;
  assign _3635_ = state_in[15:8] == 8'b11101001;
  assign _3636_ = state_in[15:8] == 8'b11101000;
  assign _3637_ = state_in[15:8] == 8'b11100111;
  assign _3638_ = state_in[15:8] == 8'b11100110;
  assign _3639_ = state_in[15:8] == 8'b11100101;
  assign _3640_ = state_in[15:8] == 8'b11100100;
  assign _3641_ = state_in[15:8] == 8'b11100011;
  assign _3642_ = state_in[15:8] == 8'b11100010;
  assign _3643_ = state_in[15:8] == 8'b11100001;
  assign _3644_ = state_in[15:8] == 8'b11100000;
  assign _3645_ = state_in[15:8] == 8'b11011111;
  assign _3646_ = state_in[15:8] == 8'b11011110;
  assign _3647_ = state_in[15:8] == 8'b11011101;
  assign _3648_ = state_in[15:8] == 8'b11011100;
  assign _3649_ = state_in[15:8] == 8'b11011011;
  assign _3650_ = state_in[15:8] == 8'b11011010;
  assign _3651_ = state_in[15:8] == 8'b11011001;
  assign _3652_ = state_in[15:8] == 8'b11011000;
  assign _3653_ = state_in[15:8] == 8'b11010111;
  assign _3654_ = state_in[15:8] == 8'b11010110;
  assign _3655_ = state_in[15:8] == 8'b11010101;
  assign _3656_ = state_in[15:8] == 8'b11010100;
  assign _3657_ = state_in[15:8] == 8'b11010011;
  assign _3658_ = state_in[15:8] == 8'b11010010;
  assign _3659_ = state_in[15:8] == 8'b11010001;
  assign _3660_ = state_in[15:8] == 8'b11010000;
  assign _3661_ = state_in[15:8] == 8'b11001111;
  assign _3662_ = state_in[15:8] == 8'b11001110;
  assign _3663_ = state_in[15:8] == 8'b11001101;
  assign _3664_ = state_in[15:8] == 8'b11001100;
  assign _3665_ = state_in[15:8] == 8'b11001011;
  assign _3666_ = state_in[15:8] == 8'b11001010;
  assign _3667_ = state_in[15:8] == 8'b11001001;
  assign _3668_ = state_in[15:8] == 8'b11001000;
  assign _3669_ = state_in[15:8] == 8'b11000111;
  assign _3670_ = state_in[15:8] == 8'b11000110;
  assign _3671_ = state_in[15:8] == 8'b11000101;
  assign _3672_ = state_in[15:8] == 8'b11000100;
  assign _3673_ = state_in[15:8] == 8'b11000011;
  assign _3674_ = state_in[15:8] == 8'b11000010;
  assign _3675_ = state_in[15:8] == 8'b11000001;
  assign _3676_ = state_in[15:8] == 8'b11000000;
  assign _3677_ = state_in[15:8] == 8'b10111111;
  assign _3678_ = state_in[15:8] == 8'b10111110;
  assign _3679_ = state_in[15:8] == 8'b10111101;
  assign _3680_ = state_in[15:8] == 8'b10111100;
  assign _3681_ = state_in[15:8] == 8'b10111011;
  assign _3682_ = state_in[15:8] == 8'b10111010;
  assign _3683_ = state_in[15:8] == 8'b10111001;
  assign _3684_ = state_in[15:8] == 8'b10111000;
  assign _3685_ = state_in[15:8] == 8'b10110111;
  assign _3686_ = state_in[15:8] == 8'b10110110;
  assign _3687_ = state_in[15:8] == 8'b10110101;
  assign _3688_ = state_in[15:8] == 8'b10110100;
  assign _3689_ = state_in[15:8] == 8'b10110011;
  assign _3690_ = state_in[15:8] == 8'b10110010;
  assign _3691_ = state_in[15:8] == 8'b10110001;
  assign _3692_ = state_in[15:8] == 8'b10110000;
  assign _3693_ = state_in[15:8] == 8'b10101111;
  assign _3694_ = state_in[15:8] == 8'b10101110;
  assign _3695_ = state_in[15:8] == 8'b10101101;
  assign _3696_ = state_in[15:8] == 8'b10101100;
  assign _3697_ = state_in[15:8] == 8'b10101011;
  assign _3698_ = state_in[15:8] == 8'b10101010;
  assign _3699_ = state_in[15:8] == 8'b10101001;
  assign _3700_ = state_in[15:8] == 8'b10101000;
  assign _3701_ = state_in[15:8] == 8'b10100111;
  assign _3702_ = state_in[15:8] == 8'b10100110;
  assign _3703_ = state_in[15:8] == 8'b10100101;
  assign _3704_ = state_in[15:8] == 8'b10100100;
  assign _3705_ = state_in[15:8] == 8'b10100011;
  assign _3706_ = state_in[15:8] == 8'b10100010;
  assign _3707_ = state_in[15:8] == 8'b10100001;
  assign _3708_ = state_in[15:8] == 8'b10100000;
  assign _3709_ = state_in[15:8] == 8'b10011111;
  assign _3710_ = state_in[15:8] == 8'b10011110;
  assign _3711_ = state_in[15:8] == 8'b10011101;
  assign _3712_ = state_in[15:8] == 8'b10011100;
  assign _3713_ = state_in[15:8] == 8'b10011011;
  assign _3714_ = state_in[15:8] == 8'b10011010;
  assign _3715_ = state_in[15:8] == 8'b10011001;
  assign _3716_ = state_in[15:8] == 8'b10011000;
  assign _3717_ = state_in[15:8] == 8'b10010111;
  assign _3718_ = state_in[15:8] == 8'b10010110;
  assign _3719_ = state_in[15:8] == 8'b10010101;
  assign _3720_ = state_in[15:8] == 8'b10010100;
  assign _3721_ = state_in[15:8] == 8'b10010011;
  assign _3722_ = state_in[15:8] == 8'b10010010;
  assign _3723_ = state_in[15:8] == 8'b10010001;
  assign _3724_ = state_in[15:8] == 8'b10010000;
  assign _3725_ = state_in[15:8] == 8'b10001111;
  assign _3726_ = state_in[15:8] == 8'b10001110;
  assign _3727_ = state_in[15:8] == 8'b10001101;
  assign _3728_ = state_in[15:8] == 8'b10001100;
  assign _3729_ = state_in[15:8] == 8'b10001011;
  assign _3730_ = state_in[15:8] == 8'b10001010;
  assign _3731_ = state_in[15:8] == 8'b10001001;
  assign _3732_ = state_in[15:8] == 8'b10001000;
  assign _3733_ = state_in[15:8] == 8'b10000111;
  assign _3734_ = state_in[15:8] == 8'b10000110;
  assign _3735_ = state_in[15:8] == 8'b10000101;
  assign _3736_ = state_in[15:8] == 8'b10000100;
  assign _3737_ = state_in[15:8] == 8'b10000011;
  assign _3738_ = state_in[15:8] == 8'b10000010;
  assign _3739_ = state_in[15:8] == 8'b10000001;
  assign _3740_ = state_in[15:8] == 8'b10000000;
  assign _3741_ = state_in[15:8] == 7'b1111111;
  assign _3742_ = state_in[15:8] == 7'b1111110;
  assign _3743_ = state_in[15:8] == 7'b1111101;
  assign _3744_ = state_in[15:8] == 7'b1111100;
  assign _3745_ = state_in[15:8] == 7'b1111011;
  assign _3746_ = state_in[15:8] == 7'b1111010;
  assign _3747_ = state_in[15:8] == 7'b1111001;
  assign _3748_ = state_in[15:8] == 7'b1111000;
  assign _3749_ = state_in[15:8] == 7'b1110111;
  assign _3750_ = state_in[15:8] == 7'b1110110;
  assign _3751_ = state_in[15:8] == 7'b1110101;
  assign _3752_ = state_in[15:8] == 7'b1110100;
  assign _3753_ = state_in[15:8] == 7'b1110011;
  assign _3754_ = state_in[15:8] == 7'b1110010;
  assign _3755_ = state_in[15:8] == 7'b1110001;
  assign _3756_ = state_in[15:8] == 7'b1110000;
  assign _3757_ = state_in[15:8] == 7'b1101111;
  assign _3758_ = state_in[15:8] == 7'b1101110;
  assign _3759_ = state_in[15:8] == 7'b1101101;
  assign _3760_ = state_in[15:8] == 7'b1101100;
  assign _3761_ = state_in[15:8] == 7'b1101011;
  assign _3762_ = state_in[15:8] == 7'b1101010;
  assign _3763_ = state_in[15:8] == 7'b1101001;
  assign _3764_ = state_in[15:8] == 7'b1101000;
  assign _3765_ = state_in[15:8] == 7'b1100111;
  assign _3766_ = state_in[15:8] == 7'b1100110;
  assign _3767_ = state_in[15:8] == 7'b1100101;
  assign _3768_ = state_in[15:8] == 7'b1100100;
  assign _3769_ = state_in[15:8] == 7'b1100011;
  assign _3770_ = state_in[15:8] == 7'b1100010;
  assign _3771_ = state_in[15:8] == 7'b1100001;
  assign _3772_ = state_in[15:8] == 7'b1100000;
  assign _3773_ = state_in[15:8] == 7'b1011111;
  assign _3774_ = state_in[15:8] == 7'b1011110;
  assign _3775_ = state_in[15:8] == 7'b1011101;
  assign _3776_ = state_in[15:8] == 7'b1011100;
  assign _3777_ = state_in[15:8] == 7'b1011011;
  assign _3778_ = state_in[15:8] == 7'b1011010;
  assign _3779_ = state_in[15:8] == 7'b1011001;
  assign _3780_ = state_in[15:8] == 7'b1011000;
  assign _3781_ = state_in[15:8] == 7'b1010111;
  assign _3782_ = state_in[15:8] == 7'b1010110;
  assign _3783_ = state_in[15:8] == 7'b1010101;
  assign _3784_ = state_in[15:8] == 7'b1010100;
  assign _3785_ = state_in[15:8] == 7'b1010011;
  assign _3786_ = state_in[15:8] == 7'b1010010;
  assign _3787_ = state_in[15:8] == 7'b1010001;
  assign _3788_ = state_in[15:8] == 7'b1010000;
  assign _3789_ = state_in[15:8] == 7'b1001111;
  assign _3790_ = state_in[15:8] == 7'b1001110;
  assign _3791_ = state_in[15:8] == 7'b1001101;
  assign _3792_ = state_in[15:8] == 7'b1001100;
  assign _3793_ = state_in[15:8] == 7'b1001011;
  assign _3794_ = state_in[15:8] == 7'b1001010;
  assign _3795_ = state_in[15:8] == 7'b1001001;
  assign _3796_ = state_in[15:8] == 7'b1001000;
  assign _3797_ = state_in[15:8] == 7'b1000111;
  assign _3798_ = state_in[15:8] == 7'b1000110;
  assign _3799_ = state_in[15:8] == 7'b1000101;
  assign _3800_ = state_in[15:8] == 7'b1000100;
  assign _3801_ = state_in[15:8] == 7'b1000011;
  assign _3802_ = state_in[15:8] == 7'b1000010;
  assign _3803_ = state_in[15:8] == 7'b1000001;
  assign _3804_ = state_in[15:8] == 7'b1000000;
  assign _3805_ = state_in[15:8] == 6'b111111;
  assign _3806_ = state_in[15:8] == 6'b111110;
  assign _3807_ = state_in[15:8] == 6'b111101;
  assign _3808_ = state_in[15:8] == 6'b111100;
  assign _3809_ = state_in[15:8] == 6'b111011;
  assign _3810_ = state_in[15:8] == 6'b111010;
  assign _3811_ = state_in[15:8] == 6'b111001;
  assign _3812_ = state_in[15:8] == 6'b111000;
  assign _3813_ = state_in[15:8] == 6'b110111;
  assign _3814_ = state_in[15:8] == 6'b110110;
  assign _3815_ = state_in[15:8] == 6'b110101;
  assign _3816_ = state_in[15:8] == 6'b110100;
  assign _3817_ = state_in[15:8] == 6'b110011;
  assign _3818_ = state_in[15:8] == 6'b110010;
  assign _3819_ = state_in[15:8] == 6'b110001;
  assign _3820_ = state_in[15:8] == 6'b110000;
  assign _3821_ = state_in[15:8] == 6'b101111;
  assign _3822_ = state_in[15:8] == 6'b101110;
  assign _3823_ = state_in[15:8] == 6'b101101;
  assign _3824_ = state_in[15:8] == 6'b101100;
  assign _3825_ = state_in[15:8] == 6'b101011;
  assign _3826_ = state_in[15:8] == 6'b101010;
  assign _3827_ = state_in[15:8] == 6'b101001;
  assign _3828_ = state_in[15:8] == 6'b101000;
  assign _3829_ = state_in[15:8] == 6'b100111;
  assign _3830_ = state_in[15:8] == 6'b100110;
  assign _3831_ = state_in[15:8] == 6'b100101;
  assign _3832_ = state_in[15:8] == 6'b100100;
  assign _3833_ = state_in[15:8] == 6'b100011;
  assign _3834_ = state_in[15:8] == 6'b100010;
  assign _3835_ = state_in[15:8] == 6'b100001;
  assign _3836_ = state_in[15:8] == 6'b100000;
  assign _3837_ = state_in[15:8] == 5'b11111;
  assign _3838_ = state_in[15:8] == 5'b11110;
  assign _3839_ = state_in[15:8] == 5'b11101;
  assign _3840_ = state_in[15:8] == 5'b11100;
  assign _3841_ = state_in[15:8] == 5'b11011;
  assign _3842_ = state_in[15:8] == 5'b11010;
  assign _3843_ = state_in[15:8] == 5'b11001;
  assign _3844_ = state_in[15:8] == 5'b11000;
  assign _3845_ = state_in[15:8] == 5'b10111;
  assign _3846_ = state_in[15:8] == 5'b10110;
  assign _3847_ = state_in[15:8] == 5'b10101;
  assign _3848_ = state_in[15:8] == 5'b10100;
  assign _3849_ = state_in[15:8] == 5'b10011;
  assign _3850_ = state_in[15:8] == 5'b10010;
  assign _3851_ = state_in[15:8] == 5'b10001;
  assign _3852_ = state_in[15:8] == 5'b10000;
  assign _3853_ = state_in[15:8] == 4'b1111;
  assign _3854_ = state_in[15:8] == 4'b1110;
  assign _3855_ = state_in[15:8] == 4'b1101;
  assign _3856_ = state_in[15:8] == 4'b1100;
  assign _3857_ = state_in[15:8] == 4'b1011;
  assign _3858_ = state_in[15:8] == 4'b1010;
  assign _3859_ = state_in[15:8] == 4'b1001;
  assign _3860_ = state_in[15:8] == 4'b1000;
  assign _3861_ = state_in[15:8] == 3'b111;
  assign _3862_ = state_in[15:8] == 3'b110;
  assign _3863_ = state_in[15:8] == 3'b101;
  assign _3864_ = state_in[15:8] == 3'b100;
  assign _3865_ = state_in[15:8] == 2'b11;
  assign _3866_ = state_in[15:8] == 2'b10;
  assign _3867_ = state_in[15:8] == 1'b1;
  assign _3868_ = ! state_in[15:8];
  always @(posedge clk)
      \t3.t2.s4.out <= _3869_;
  logic [255:0] fangyuan30;
  assign fangyuan30 = { _3868_, _3867_, _3866_, _3865_, _3864_, _3863_, _3862_, _3861_, _3860_, _3859_, _3858_, _3857_, _3856_, _3855_, _3854_, _3853_, _3852_, _3851_, _3850_, _3849_, _3848_, _3847_, _3846_, _3845_, _3844_, _3843_, _3842_, _3841_, _3840_, _3839_, _3838_, _3837_, _3836_, _3835_, _3834_, _3833_, _3832_, _3831_, _3830_, _3829_, _3828_, _3827_, _3826_, _3825_, _3824_, _3823_, _3822_, _3821_, _3820_, _3819_, _3818_, _3817_, _3816_, _3815_, _3814_, _3813_, _3812_, _3811_, _3810_, _3809_, _3808_, _3807_, _3806_, _3805_, _3804_, _3803_, _3802_, _3801_, _3800_, _3799_, _3798_, _3797_, _3796_, _3795_, _3794_, _3793_, _3792_, _3791_, _3790_, _3789_, _3788_, _3787_, _3786_, _3785_, _3784_, _3783_, _3782_, _3781_, _3780_, _3779_, _3778_, _3777_, _3776_, _3775_, _3774_, _3773_, _3772_, _3771_, _3770_, _3769_, _3768_, _3767_, _3766_, _3765_, _3764_, _3763_, _3762_, _3761_, _3760_, _3759_, _3758_, _3757_, _3756_, _3755_, _3754_, _3753_, _3752_, _3751_, _3750_, _3749_, _3748_, _3747_, _3746_, _3745_, _3744_, _3743_, _3742_, _3741_, _3740_, _3739_, _3738_, _3737_, _3736_, _3735_, _3734_, _3733_, _3732_, _3731_, _3730_, _3729_, _3728_, _3727_, _3726_, _3725_, _3724_, _3723_, _3722_, _3721_, _3720_, _3719_, _3718_, _3717_, _3716_, _3715_, _3714_, _3713_, _3712_, _3711_, _3710_, _3709_, _3708_, _3707_, _3706_, _3705_, _3704_, _3703_, _3702_, _3701_, _3700_, _3699_, _3698_, _3697_, _3696_, _3695_, _3694_, _3693_, _3692_, _3691_, _3690_, _3689_, _3688_, _3687_, _3686_, _3685_, _3684_, _3683_, _3682_, _3681_, _3680_, _3679_, _3678_, _3677_, _3676_, _3675_, _3674_, _3673_, _3672_, _3671_, _3670_, _3669_, _3668_, _3667_, _3666_, _3665_, _3664_, _3663_, _3662_, _3661_, _3660_, _3659_, _3658_, _3657_, _3656_, _3655_, _3654_, _3653_, _3652_, _3651_, _3650_, _3649_, _3648_, _3647_, _3646_, _3645_, _3644_, _3643_, _3642_, _3641_, _3640_, _3639_, _3638_, _3637_, _3636_, _3635_, _3634_, _3633_, _3632_, _3631_, _3630_, _3629_, _3628_, _3627_, _3626_, _3625_, _3624_, _3623_, _3622_, _3621_, _3620_, _3619_, _3618_, _3617_, _3616_, _3615_, _3614_, _3613_ };

  always @(\t3.t2.s4.out or fangyuan30) begin
    casez (fangyuan30)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3869_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3869_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3869_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3869_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3869_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3869_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3869_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3869_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3869_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3869_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3869_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3869_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3869_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3869_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3869_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3869_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3869_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3869_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3869_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3869_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3869_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3869_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3869_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3869_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3869_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3869_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3869_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3869_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3869_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3869_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3869_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3869_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3869_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3869_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3869_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3869_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3869_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3869_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3869_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3869_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3869_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3869_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3869_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3869_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3869_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3869_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3869_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3869_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3869_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3869_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3869_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3869_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3869_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3869_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3869_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3869_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3869_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3869_ = 8'b11000110 ;
      default:
        _3869_ = \t3.t2.s4.out ;
    endcase
  end
  assign p33[15:8] = \t3.t3.s0.out ^ \t3.t3.s4.out ;
  always @(posedge clk)
      \t3.t3.s0.out <= _3870_;
  logic [255:0] fangyuan31;
  assign fangyuan31 = { _4126_, _4125_, _4124_, _4123_, _4122_, _4121_, _4120_, _4119_, _4118_, _4117_, _4116_, _4115_, _4114_, _4113_, _4112_, _4111_, _4110_, _4109_, _4108_, _4107_, _4106_, _4105_, _4104_, _4103_, _4102_, _4101_, _4100_, _4099_, _4098_, _4097_, _4096_, _4095_, _4094_, _4093_, _4092_, _4091_, _4090_, _4089_, _4088_, _4087_, _4086_, _4085_, _4084_, _4083_, _4082_, _4081_, _4080_, _4079_, _4078_, _4077_, _4076_, _4075_, _4074_, _4073_, _4072_, _4071_, _4070_, _4069_, _4068_, _4067_, _4066_, _4065_, _4064_, _4063_, _4062_, _4061_, _4060_, _4059_, _4058_, _4057_, _4056_, _4055_, _4054_, _4053_, _4052_, _4051_, _4050_, _4049_, _4048_, _4047_, _4046_, _4045_, _4044_, _4043_, _4042_, _4041_, _4040_, _4039_, _4038_, _4037_, _4036_, _4035_, _4034_, _4033_, _4032_, _4031_, _4030_, _4029_, _4028_, _4027_, _4026_, _4025_, _4024_, _4023_, _4022_, _4021_, _4020_, _4019_, _4018_, _4017_, _4016_, _4015_, _4014_, _4013_, _4012_, _4011_, _4010_, _4009_, _4008_, _4007_, _4006_, _4005_, _4004_, _4003_, _4002_, _4001_, _4000_, _3999_, _3998_, _3997_, _3996_, _3995_, _3994_, _3993_, _3992_, _3991_, _3990_, _3989_, _3988_, _3987_, _3986_, _3985_, _3984_, _3983_, _3982_, _3981_, _3980_, _3979_, _3978_, _3977_, _3976_, _3975_, _3974_, _3973_, _3972_, _3971_, _3970_, _3969_, _3968_, _3967_, _3966_, _3965_, _3964_, _3963_, _3962_, _3961_, _3960_, _3959_, _3958_, _3957_, _3956_, _3955_, _3954_, _3953_, _3952_, _3951_, _3950_, _3949_, _3948_, _3947_, _3946_, _3945_, _3944_, _3943_, _3942_, _3941_, _3940_, _3939_, _3938_, _3937_, _3936_, _3935_, _3934_, _3933_, _3932_, _3931_, _3930_, _3929_, _3928_, _3927_, _3926_, _3925_, _3924_, _3923_, _3922_, _3921_, _3920_, _3919_, _3918_, _3917_, _3916_, _3915_, _3914_, _3913_, _3912_, _3911_, _3910_, _3909_, _3908_, _3907_, _3906_, _3905_, _3904_, _3903_, _3902_, _3901_, _3900_, _3899_, _3898_, _3897_, _3896_, _3895_, _3894_, _3893_, _3892_, _3891_, _3890_, _3889_, _3888_, _3887_, _3886_, _3885_, _3884_, _3883_, _3882_, _3881_, _3880_, _3879_, _3878_, _3877_, _3876_, _3875_, _3874_, _3873_, _3872_, _3871_ };

  always @(\t3.t3.s0.out or fangyuan31) begin
    casez (fangyuan31)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _3870_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _3870_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _3870_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _3870_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _3870_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _3870_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _3870_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _3870_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _3870_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _3870_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _3870_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _3870_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _3870_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _3870_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _3870_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _3870_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _3870_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _3870_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _3870_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _3870_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _3870_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _3870_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _3870_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _3870_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _3870_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _3870_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _3870_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _3870_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _3870_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _3870_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _3870_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _3870_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _3870_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _3870_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _3870_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _3870_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _3870_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _3870_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _3870_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _3870_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _3870_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _3870_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _3870_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _3870_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _3870_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _3870_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _3870_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _3870_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _3870_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _3870_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _3870_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _3870_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _3870_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _3870_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _3870_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _3870_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _3870_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _3870_ = 8'b01100011 ;
      default:
        _3870_ = \t3.t3.s0.out ;
    endcase
  end
  assign _3871_ = state_in[7:0] == 8'b11111111;
  assign _3872_ = state_in[7:0] == 8'b11111110;
  assign _3873_ = state_in[7:0] == 8'b11111101;
  assign _3874_ = state_in[7:0] == 8'b11111100;
  assign _3875_ = state_in[7:0] == 8'b11111011;
  assign _3876_ = state_in[7:0] == 8'b11111010;
  assign _3877_ = state_in[7:0] == 8'b11111001;
  assign _3878_ = state_in[7:0] == 8'b11111000;
  assign _3879_ = state_in[7:0] == 8'b11110111;
  assign _3880_ = state_in[7:0] == 8'b11110110;
  assign _3881_ = state_in[7:0] == 8'b11110101;
  assign _3882_ = state_in[7:0] == 8'b11110100;
  assign _3883_ = state_in[7:0] == 8'b11110011;
  assign _3884_ = state_in[7:0] == 8'b11110010;
  assign _3885_ = state_in[7:0] == 8'b11110001;
  assign _3886_ = state_in[7:0] == 8'b11110000;
  assign _3887_ = state_in[7:0] == 8'b11101111;
  assign _3888_ = state_in[7:0] == 8'b11101110;
  assign _3889_ = state_in[7:0] == 8'b11101101;
  assign _3890_ = state_in[7:0] == 8'b11101100;
  assign _3891_ = state_in[7:0] == 8'b11101011;
  assign _3892_ = state_in[7:0] == 8'b11101010;
  assign _3893_ = state_in[7:0] == 8'b11101001;
  assign _3894_ = state_in[7:0] == 8'b11101000;
  assign _3895_ = state_in[7:0] == 8'b11100111;
  assign _3896_ = state_in[7:0] == 8'b11100110;
  assign _3897_ = state_in[7:0] == 8'b11100101;
  assign _3898_ = state_in[7:0] == 8'b11100100;
  assign _3899_ = state_in[7:0] == 8'b11100011;
  assign _3900_ = state_in[7:0] == 8'b11100010;
  assign _3901_ = state_in[7:0] == 8'b11100001;
  assign _3902_ = state_in[7:0] == 8'b11100000;
  assign _3903_ = state_in[7:0] == 8'b11011111;
  assign _3904_ = state_in[7:0] == 8'b11011110;
  assign _3905_ = state_in[7:0] == 8'b11011101;
  assign _3906_ = state_in[7:0] == 8'b11011100;
  assign _3907_ = state_in[7:0] == 8'b11011011;
  assign _3908_ = state_in[7:0] == 8'b11011010;
  assign _3909_ = state_in[7:0] == 8'b11011001;
  assign _3910_ = state_in[7:0] == 8'b11011000;
  assign _3911_ = state_in[7:0] == 8'b11010111;
  assign _3912_ = state_in[7:0] == 8'b11010110;
  assign _3913_ = state_in[7:0] == 8'b11010101;
  assign _3914_ = state_in[7:0] == 8'b11010100;
  assign _3915_ = state_in[7:0] == 8'b11010011;
  assign _3916_ = state_in[7:0] == 8'b11010010;
  assign _3917_ = state_in[7:0] == 8'b11010001;
  assign _3918_ = state_in[7:0] == 8'b11010000;
  assign _3919_ = state_in[7:0] == 8'b11001111;
  assign _3920_ = state_in[7:0] == 8'b11001110;
  assign _3921_ = state_in[7:0] == 8'b11001101;
  assign _3922_ = state_in[7:0] == 8'b11001100;
  assign _3923_ = state_in[7:0] == 8'b11001011;
  assign _3924_ = state_in[7:0] == 8'b11001010;
  assign _3925_ = state_in[7:0] == 8'b11001001;
  assign _3926_ = state_in[7:0] == 8'b11001000;
  assign _3927_ = state_in[7:0] == 8'b11000111;
  assign _3928_ = state_in[7:0] == 8'b11000110;
  assign _3929_ = state_in[7:0] == 8'b11000101;
  assign _3930_ = state_in[7:0] == 8'b11000100;
  assign _3931_ = state_in[7:0] == 8'b11000011;
  assign _3932_ = state_in[7:0] == 8'b11000010;
  assign _3933_ = state_in[7:0] == 8'b11000001;
  assign _3934_ = state_in[7:0] == 8'b11000000;
  assign _3935_ = state_in[7:0] == 8'b10111111;
  assign _3936_ = state_in[7:0] == 8'b10111110;
  assign _3937_ = state_in[7:0] == 8'b10111101;
  assign _3938_ = state_in[7:0] == 8'b10111100;
  assign _3939_ = state_in[7:0] == 8'b10111011;
  assign _3940_ = state_in[7:0] == 8'b10111010;
  assign _3941_ = state_in[7:0] == 8'b10111001;
  assign _3942_ = state_in[7:0] == 8'b10111000;
  assign _3943_ = state_in[7:0] == 8'b10110111;
  assign _3944_ = state_in[7:0] == 8'b10110110;
  assign _3945_ = state_in[7:0] == 8'b10110101;
  assign _3946_ = state_in[7:0] == 8'b10110100;
  assign _3947_ = state_in[7:0] == 8'b10110011;
  assign _3948_ = state_in[7:0] == 8'b10110010;
  assign _3949_ = state_in[7:0] == 8'b10110001;
  assign _3950_ = state_in[7:0] == 8'b10110000;
  assign _3951_ = state_in[7:0] == 8'b10101111;
  assign _3952_ = state_in[7:0] == 8'b10101110;
  assign _3953_ = state_in[7:0] == 8'b10101101;
  assign _3954_ = state_in[7:0] == 8'b10101100;
  assign _3955_ = state_in[7:0] == 8'b10101011;
  assign _3956_ = state_in[7:0] == 8'b10101010;
  assign _3957_ = state_in[7:0] == 8'b10101001;
  assign _3958_ = state_in[7:0] == 8'b10101000;
  assign _3959_ = state_in[7:0] == 8'b10100111;
  assign _3960_ = state_in[7:0] == 8'b10100110;
  assign _3961_ = state_in[7:0] == 8'b10100101;
  assign _3962_ = state_in[7:0] == 8'b10100100;
  assign _3963_ = state_in[7:0] == 8'b10100011;
  assign _3964_ = state_in[7:0] == 8'b10100010;
  assign _3965_ = state_in[7:0] == 8'b10100001;
  assign _3966_ = state_in[7:0] == 8'b10100000;
  assign _3967_ = state_in[7:0] == 8'b10011111;
  assign _3968_ = state_in[7:0] == 8'b10011110;
  assign _3969_ = state_in[7:0] == 8'b10011101;
  assign _3970_ = state_in[7:0] == 8'b10011100;
  assign _3971_ = state_in[7:0] == 8'b10011011;
  assign _3972_ = state_in[7:0] == 8'b10011010;
  assign _3973_ = state_in[7:0] == 8'b10011001;
  assign _3974_ = state_in[7:0] == 8'b10011000;
  assign _3975_ = state_in[7:0] == 8'b10010111;
  assign _3976_ = state_in[7:0] == 8'b10010110;
  assign _3977_ = state_in[7:0] == 8'b10010101;
  assign _3978_ = state_in[7:0] == 8'b10010100;
  assign _3979_ = state_in[7:0] == 8'b10010011;
  assign _3980_ = state_in[7:0] == 8'b10010010;
  assign _3981_ = state_in[7:0] == 8'b10010001;
  assign _3982_ = state_in[7:0] == 8'b10010000;
  assign _3983_ = state_in[7:0] == 8'b10001111;
  assign _3984_ = state_in[7:0] == 8'b10001110;
  assign _3985_ = state_in[7:0] == 8'b10001101;
  assign _3986_ = state_in[7:0] == 8'b10001100;
  assign _3987_ = state_in[7:0] == 8'b10001011;
  assign _3988_ = state_in[7:0] == 8'b10001010;
  assign _3989_ = state_in[7:0] == 8'b10001001;
  assign _3990_ = state_in[7:0] == 8'b10001000;
  assign _3991_ = state_in[7:0] == 8'b10000111;
  assign _3992_ = state_in[7:0] == 8'b10000110;
  assign _3993_ = state_in[7:0] == 8'b10000101;
  assign _3994_ = state_in[7:0] == 8'b10000100;
  assign _3995_ = state_in[7:0] == 8'b10000011;
  assign _3996_ = state_in[7:0] == 8'b10000010;
  assign _3997_ = state_in[7:0] == 8'b10000001;
  assign _3998_ = state_in[7:0] == 8'b10000000;
  assign _3999_ = state_in[7:0] == 7'b1111111;
  assign _4000_ = state_in[7:0] == 7'b1111110;
  assign _4001_ = state_in[7:0] == 7'b1111101;
  assign _4002_ = state_in[7:0] == 7'b1111100;
  assign _4003_ = state_in[7:0] == 7'b1111011;
  assign _4004_ = state_in[7:0] == 7'b1111010;
  assign _4005_ = state_in[7:0] == 7'b1111001;
  assign _4006_ = state_in[7:0] == 7'b1111000;
  assign _4007_ = state_in[7:0] == 7'b1110111;
  assign _4008_ = state_in[7:0] == 7'b1110110;
  assign _4009_ = state_in[7:0] == 7'b1110101;
  assign _4010_ = state_in[7:0] == 7'b1110100;
  assign _4011_ = state_in[7:0] == 7'b1110011;
  assign _4012_ = state_in[7:0] == 7'b1110010;
  assign _4013_ = state_in[7:0] == 7'b1110001;
  assign _4014_ = state_in[7:0] == 7'b1110000;
  assign _4015_ = state_in[7:0] == 7'b1101111;
  assign _4016_ = state_in[7:0] == 7'b1101110;
  assign _4017_ = state_in[7:0] == 7'b1101101;
  assign _4018_ = state_in[7:0] == 7'b1101100;
  assign _4019_ = state_in[7:0] == 7'b1101011;
  assign _4020_ = state_in[7:0] == 7'b1101010;
  assign _4021_ = state_in[7:0] == 7'b1101001;
  assign _4022_ = state_in[7:0] == 7'b1101000;
  assign _4023_ = state_in[7:0] == 7'b1100111;
  assign _4024_ = state_in[7:0] == 7'b1100110;
  assign _4025_ = state_in[7:0] == 7'b1100101;
  assign _4026_ = state_in[7:0] == 7'b1100100;
  assign _4027_ = state_in[7:0] == 7'b1100011;
  assign _4028_ = state_in[7:0] == 7'b1100010;
  assign _4029_ = state_in[7:0] == 7'b1100001;
  assign _4030_ = state_in[7:0] == 7'b1100000;
  assign _4031_ = state_in[7:0] == 7'b1011111;
  assign _4032_ = state_in[7:0] == 7'b1011110;
  assign _4033_ = state_in[7:0] == 7'b1011101;
  assign _4034_ = state_in[7:0] == 7'b1011100;
  assign _4035_ = state_in[7:0] == 7'b1011011;
  assign _4036_ = state_in[7:0] == 7'b1011010;
  assign _4037_ = state_in[7:0] == 7'b1011001;
  assign _4038_ = state_in[7:0] == 7'b1011000;
  assign _4039_ = state_in[7:0] == 7'b1010111;
  assign _4040_ = state_in[7:0] == 7'b1010110;
  assign _4041_ = state_in[7:0] == 7'b1010101;
  assign _4042_ = state_in[7:0] == 7'b1010100;
  assign _4043_ = state_in[7:0] == 7'b1010011;
  assign _4044_ = state_in[7:0] == 7'b1010010;
  assign _4045_ = state_in[7:0] == 7'b1010001;
  assign _4046_ = state_in[7:0] == 7'b1010000;
  assign _4047_ = state_in[7:0] == 7'b1001111;
  assign _4048_ = state_in[7:0] == 7'b1001110;
  assign _4049_ = state_in[7:0] == 7'b1001101;
  assign _4050_ = state_in[7:0] == 7'b1001100;
  assign _4051_ = state_in[7:0] == 7'b1001011;
  assign _4052_ = state_in[7:0] == 7'b1001010;
  assign _4053_ = state_in[7:0] == 7'b1001001;
  assign _4054_ = state_in[7:0] == 7'b1001000;
  assign _4055_ = state_in[7:0] == 7'b1000111;
  assign _4056_ = state_in[7:0] == 7'b1000110;
  assign _4057_ = state_in[7:0] == 7'b1000101;
  assign _4058_ = state_in[7:0] == 7'b1000100;
  assign _4059_ = state_in[7:0] == 7'b1000011;
  assign _4060_ = state_in[7:0] == 7'b1000010;
  assign _4061_ = state_in[7:0] == 7'b1000001;
  assign _4062_ = state_in[7:0] == 7'b1000000;
  assign _4063_ = state_in[7:0] == 6'b111111;
  assign _4064_ = state_in[7:0] == 6'b111110;
  assign _4065_ = state_in[7:0] == 6'b111101;
  assign _4066_ = state_in[7:0] == 6'b111100;
  assign _4067_ = state_in[7:0] == 6'b111011;
  assign _4068_ = state_in[7:0] == 6'b111010;
  assign _4069_ = state_in[7:0] == 6'b111001;
  assign _4070_ = state_in[7:0] == 6'b111000;
  assign _4071_ = state_in[7:0] == 6'b110111;
  assign _4072_ = state_in[7:0] == 6'b110110;
  assign _4073_ = state_in[7:0] == 6'b110101;
  assign _4074_ = state_in[7:0] == 6'b110100;
  assign _4075_ = state_in[7:0] == 6'b110011;
  assign _4076_ = state_in[7:0] == 6'b110010;
  assign _4077_ = state_in[7:0] == 6'b110001;
  assign _4078_ = state_in[7:0] == 6'b110000;
  assign _4079_ = state_in[7:0] == 6'b101111;
  assign _4080_ = state_in[7:0] == 6'b101110;
  assign _4081_ = state_in[7:0] == 6'b101101;
  assign _4082_ = state_in[7:0] == 6'b101100;
  assign _4083_ = state_in[7:0] == 6'b101011;
  assign _4084_ = state_in[7:0] == 6'b101010;
  assign _4085_ = state_in[7:0] == 6'b101001;
  assign _4086_ = state_in[7:0] == 6'b101000;
  assign _4087_ = state_in[7:0] == 6'b100111;
  assign _4088_ = state_in[7:0] == 6'b100110;
  assign _4089_ = state_in[7:0] == 6'b100101;
  assign _4090_ = state_in[7:0] == 6'b100100;
  assign _4091_ = state_in[7:0] == 6'b100011;
  assign _4092_ = state_in[7:0] == 6'b100010;
  assign _4093_ = state_in[7:0] == 6'b100001;
  assign _4094_ = state_in[7:0] == 6'b100000;
  assign _4095_ = state_in[7:0] == 5'b11111;
  assign _4096_ = state_in[7:0] == 5'b11110;
  assign _4097_ = state_in[7:0] == 5'b11101;
  assign _4098_ = state_in[7:0] == 5'b11100;
  assign _4099_ = state_in[7:0] == 5'b11011;
  assign _4100_ = state_in[7:0] == 5'b11010;
  assign _4101_ = state_in[7:0] == 5'b11001;
  assign _4102_ = state_in[7:0] == 5'b11000;
  assign _4103_ = state_in[7:0] == 5'b10111;
  assign _4104_ = state_in[7:0] == 5'b10110;
  assign _4105_ = state_in[7:0] == 5'b10101;
  assign _4106_ = state_in[7:0] == 5'b10100;
  assign _4107_ = state_in[7:0] == 5'b10011;
  assign _4108_ = state_in[7:0] == 5'b10010;
  assign _4109_ = state_in[7:0] == 5'b10001;
  assign _4110_ = state_in[7:0] == 5'b10000;
  assign _4111_ = state_in[7:0] == 4'b1111;
  assign _4112_ = state_in[7:0] == 4'b1110;
  assign _4113_ = state_in[7:0] == 4'b1101;
  assign _4114_ = state_in[7:0] == 4'b1100;
  assign _4115_ = state_in[7:0] == 4'b1011;
  assign _4116_ = state_in[7:0] == 4'b1010;
  assign _4117_ = state_in[7:0] == 4'b1001;
  assign _4118_ = state_in[7:0] == 4'b1000;
  assign _4119_ = state_in[7:0] == 3'b111;
  assign _4120_ = state_in[7:0] == 3'b110;
  assign _4121_ = state_in[7:0] == 3'b101;
  assign _4122_ = state_in[7:0] == 3'b100;
  assign _4123_ = state_in[7:0] == 2'b11;
  assign _4124_ = state_in[7:0] == 2'b10;
  assign _4125_ = state_in[7:0] == 1'b1;
  assign _4126_ = ! state_in[7:0];
  always @(posedge clk)
      \t3.t3.s4.out <= _4127_;
  logic [255:0] fangyuan32;
  assign fangyuan32 = { _4126_, _4125_, _4124_, _4123_, _4122_, _4121_, _4120_, _4119_, _4118_, _4117_, _4116_, _4115_, _4114_, _4113_, _4112_, _4111_, _4110_, _4109_, _4108_, _4107_, _4106_, _4105_, _4104_, _4103_, _4102_, _4101_, _4100_, _4099_, _4098_, _4097_, _4096_, _4095_, _4094_, _4093_, _4092_, _4091_, _4090_, _4089_, _4088_, _4087_, _4086_, _4085_, _4084_, _4083_, _4082_, _4081_, _4080_, _4079_, _4078_, _4077_, _4076_, _4075_, _4074_, _4073_, _4072_, _4071_, _4070_, _4069_, _4068_, _4067_, _4066_, _4065_, _4064_, _4063_, _4062_, _4061_, _4060_, _4059_, _4058_, _4057_, _4056_, _4055_, _4054_, _4053_, _4052_, _4051_, _4050_, _4049_, _4048_, _4047_, _4046_, _4045_, _4044_, _4043_, _4042_, _4041_, _4040_, _4039_, _4038_, _4037_, _4036_, _4035_, _4034_, _4033_, _4032_, _4031_, _4030_, _4029_, _4028_, _4027_, _4026_, _4025_, _4024_, _4023_, _4022_, _4021_, _4020_, _4019_, _4018_, _4017_, _4016_, _4015_, _4014_, _4013_, _4012_, _4011_, _4010_, _4009_, _4008_, _4007_, _4006_, _4005_, _4004_, _4003_, _4002_, _4001_, _4000_, _3999_, _3998_, _3997_, _3996_, _3995_, _3994_, _3993_, _3992_, _3991_, _3990_, _3989_, _3988_, _3987_, _3986_, _3985_, _3984_, _3983_, _3982_, _3981_, _3980_, _3979_, _3978_, _3977_, _3976_, _3975_, _3974_, _3973_, _3972_, _3971_, _3970_, _3969_, _3968_, _3967_, _3966_, _3965_, _3964_, _3963_, _3962_, _3961_, _3960_, _3959_, _3958_, _3957_, _3956_, _3955_, _3954_, _3953_, _3952_, _3951_, _3950_, _3949_, _3948_, _3947_, _3946_, _3945_, _3944_, _3943_, _3942_, _3941_, _3940_, _3939_, _3938_, _3937_, _3936_, _3935_, _3934_, _3933_, _3932_, _3931_, _3930_, _3929_, _3928_, _3927_, _3926_, _3925_, _3924_, _3923_, _3922_, _3921_, _3920_, _3919_, _3918_, _3917_, _3916_, _3915_, _3914_, _3913_, _3912_, _3911_, _3910_, _3909_, _3908_, _3907_, _3906_, _3905_, _3904_, _3903_, _3902_, _3901_, _3900_, _3899_, _3898_, _3897_, _3896_, _3895_, _3894_, _3893_, _3892_, _3891_, _3890_, _3889_, _3888_, _3887_, _3886_, _3885_, _3884_, _3883_, _3882_, _3881_, _3880_, _3879_, _3878_, _3877_, _3876_, _3875_, _3874_, _3873_, _3872_, _3871_ };

  always @(\t3.t3.s4.out or fangyuan32) begin
    casez (fangyuan32)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _4127_ = 8'b00101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _4127_ = 8'b01101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _4127_ = 8'b10101000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _4127_ = 8'b01111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _4127_ = 8'b00011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _4127_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _4127_ = 8'b00101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _4127_ = 8'b10000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _4127_ = 8'b11010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _4127_ = 8'b10000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _4127_ = 8'b11010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _4127_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _4127_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _4127_ = 8'b00001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _4127_ = 8'b01011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _4127_ = 8'b00000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _4127_ = 8'b10100101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _4127_ = 8'b01010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _4127_ = 8'b10101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _4127_ = 8'b10000111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _4127_ = 8'b11001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _4127_ = 8'b00010101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _4127_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _4127_ = 8'b00101101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _4127_ = 8'b00110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _4127_ = 8'b00000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _4127_ = 8'b10101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _4127_ = 8'b11010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _4127_ = 8'b00100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _4127_ = 8'b00101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _4127_ = 8'b11101011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _4127_ = 8'b11011001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _4127_ = 8'b00100111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _4127_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _4127_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _4127_ = 8'b00010111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _4127_ = 8'b01101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _4127_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _4127_ = 8'b01101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _4127_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _4127_ = 8'b00011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _4127_ = 8'b11110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _4127_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _4127_ = 8'b10010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _4127_ = 8'b11001100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _4127_ = 8'b01110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _4127_ = 8'b01111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _4127_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _4127_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _4127_ = 8'b00001101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _4127_ = 8'b01100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _4127_ = 8'b10010110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _4127_ = 8'b00111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _4127_ = 8'b11101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _4127_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _4127_ = 8'b11001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _4127_ = 8'b10010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100110 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010011 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011110 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111101 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110111 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110110 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10100100 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011100 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110110 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110100 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011101 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00010010 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111111 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001110 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011011 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100100 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001110 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101111 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001010 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110111 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00110000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011101 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000110 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00001000 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00101010 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100010 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10101011 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100010 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010001 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010001 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101000 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10000011 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110101 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01111110 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01101100 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001100 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00111101 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100001 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01110101 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10011011 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100100 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010011 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00100011 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000101 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01011111 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110011 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01000001 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111011 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001110 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110010 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101111 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111010 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00011111 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10001111 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101100 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01001101 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10110101 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11100111 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01010110 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11001110 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b00000010 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b01100000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b10010001 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11011110 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11010110 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111111 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11110110 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11101110 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11111000 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _4127_ = 8'b11000110 ;
      default:
        _4127_ = \t3.t3.s4.out ;
    endcase
  end
  logic [31:0] fangyuan33;
  assign fangyuan33 = { \t0.t0.s4.out , \t0.t0.s0.out , \t0.t0.s0.out , p00[7:0] };
  logic [31:0] fangyuan34;
  assign fangyuan34 = { p11[31:24], \t1.t1.s4.out , \t1.t1.s0.out , \t1.t1.s0.out };

  assign _4128_ = fangyuan33 ^ fangyuan34;
  logic [31:0] fangyuan35;
  assign fangyuan35 = { \t2.t2.s0.out , p22[23:16], \t2.t2.s4.out , \t2.t2.s0.out };

  assign _4129_ = _4128_ ^ fangyuan35;
  logic [31:0] fangyuan36;
  assign fangyuan36 = { \t3.t3.s0.out , \t3.t3.s0.out , p33[15:8], \t3.t3.s4.out };

  assign _4130_ = _4129_ ^ fangyuan36;
  assign z0 = _4130_ ^ key[127:96];
  logic [31:0] fangyuan37;
  assign fangyuan37 = { \t0.t3.s0.out , \t0.t3.s0.out , p03[15:8], \t0.t3.s4.out };
  logic [31:0] fangyuan38;
  assign fangyuan38 = { \t1.t0.s4.out , \t1.t0.s0.out , \t1.t0.s0.out , p10[7:0] };

  assign _4131_ = fangyuan37 ^ fangyuan38;
  logic [31:0] fangyuan39;
  assign fangyuan39 = { p21[31:24], \t2.t1.s4.out , \t2.t1.s0.out , \t2.t1.s0.out };

  assign _4132_ = _4131_ ^ fangyuan39;
  logic [31:0] fangyuan40;
  assign fangyuan40 = { \t3.t2.s0.out , p32[23:16], \t3.t2.s4.out , \t3.t2.s0.out };

  assign _4133_ = _4132_ ^ fangyuan40;
  assign z1 = _4133_ ^ key[95:64];
  logic [31:0] fangyuan41;
  assign fangyuan41 = { \t2.t0.s4.out , \t2.t0.s0.out , \t2.t0.s0.out , p20[7:0] };

  assign _4134_ = _4136_ ^ fangyuan41;
  logic [31:0] fangyuan42;
  assign fangyuan42 = { p31[31:24], \t3.t1.s4.out , \t3.t1.s0.out , \t3.t1.s0.out };

  assign _4135_ = _4134_ ^ fangyuan42;
  assign z2 = _4135_ ^ key[63:32];
  logic [31:0] fangyuan43;
  assign fangyuan43 = { \t0.t2.s0.out , p02[23:16], \t0.t2.s4.out , \t0.t2.s0.out };
  logic [31:0] fangyuan44;
  assign fangyuan44 = { \t1.t3.s0.out , \t1.t3.s0.out , p13[15:8], \t1.t3.s4.out };

  assign _4136_ = fangyuan43 ^ fangyuan44;
  logic [31:0] fangyuan45;
  assign fangyuan45 = { p01[31:24], \t0.t1.s4.out , \t0.t1.s0.out , \t0.t1.s0.out };
  logic [31:0] fangyuan46;
  assign fangyuan46 = { \t1.t2.s0.out , p12[23:16], \t1.t2.s4.out , \t1.t2.s0.out };

  assign _4137_ = fangyuan45 ^ fangyuan46;
  logic [31:0] fangyuan47;
  assign fangyuan47 = { \t2.t3.s0.out , \t2.t3.s0.out , p23[15:8], \t2.t3.s4.out };

  assign _4138_ = _4137_ ^ fangyuan47;
  logic [31:0] fangyuan48;
  assign fangyuan48 = { \t3.t0.s4.out , \t3.t0.s0.out , \t3.t0.s0.out , p30[7:0] };

  assign _4139_ = _4138_ ^ fangyuan48;
  assign z3 = _4139_ ^ key[31:0];
  assign k0 = key[127:96];
  assign k1 = key[95:64];
  assign k2 = key[63:32];
  assign k3 = key[31:0];
  assign p00[31:8] = { \t0.t0.s4.out , \t0.t0.s0.out , \t0.t0.s0.out };
  assign p01[23:0] = { \t0.t1.s4.out , \t0.t1.s0.out , \t0.t1.s0.out };
  assign p02[31:24] = { \t0.t2.s0.out };
  assign p02[15:0] = { \t0.t2.s4.out, \t0.t2.s0.out };
  assign p03[31:16] = { \t0.t3.s0.out, \t0.t3.s0.out };
  assign p03[7:0] = { \t0.t3.s4.out };
  assign p10[31:8] = { \t1.t0.s4.out , \t1.t0.s0.out , \t1.t0.s0.out };
  assign p11[23:0] = { \t1.t1.s4.out , \t1.t1.s0.out , \t1.t1.s0.out };
  assign p12[31:24] = { \t1.t2.s0.out };
  assign p12[15:0] = { \t1.t2.s4.out, \t1.t2.s0.out };
  assign p13[31:16] = { \t1.t3.s0.out, \t1.t3.s0.out };
  assign p13[7:0] = { \t1.t3.s4.out };
  assign p20[31:8] = { \t2.t0.s4.out , \t2.t0.s0.out , \t2.t0.s0.out };
  assign p21[23:0] = { \t2.t1.s4.out , \t2.t1.s0.out , \t2.t1.s0.out };
  assign p22[31:24] = { \t2.t2.s0.out };
  assign p22[15:0] = { \t2.t2.s4.out, \t2.t2.s0.out };
  assign p23[31:16] = { \t2.t3.s0.out, \t2.t3.s0.out };
  assign p23[7:0] = { \t2.t3.s4.out };
  assign p30[31:8] = { \t3.t0.s4.out , \t3.t0.s0.out , \t3.t0.s0.out };
  assign p31[23:0] = { \t3.t1.s4.out , \t3.t1.s0.out , \t3.t1.s0.out };
  assign p32[31:24] = { \t3.t2.s0.out };
  assign p32[15:0] = { \t3.t2.s4.out, \t3.t2.s0.out };
  assign p33[31:16] = { \t3.t3.s0.out, \t3.t3.s0.out };
  assign p33[7:0] = { \t3.t3.s4.out };
  assign s0 = state_in[127:96];
  assign s1 = state_in[95:64];
  assign s2 = state_in[63:32];
  assign s3 = state_in[31:0];
  assign \t0.b0 = state_in[127:120];
  assign \t0.b1 = state_in[119:112];
  assign \t0.b2 = state_in[111:104];
  assign \t0.b3 = state_in[103:96];
  assign \t0.clk = clk;
  assign \t0.p0 = { \t0.t0.s4.out , \t0.t0.s0.out , \t0.t0.s0.out , p00[7:0] };
  assign \t0.p1 = { p01[31:24], \t0.t1.s4.out , \t0.t1.s0.out , \t0.t1.s0.out };
  assign \t0.p2 = { \t0.t2.s0.out , p02[23:16], \t0.t2.s4.out , \t0.t2.s0.out };
  assign \t0.p3 = { \t0.t3.s0.out , \t0.t3.s0.out , p03[15:8], \t0.t3.s4.out };
  assign \t0.state = state_in[127:96];
  assign \t0.t0.clk = clk;
  assign \t0.t0.in = state_in[127:120];
  assign \t0.t0.out = { \t0.t0.s0.out , \t0.t0.s0.out , p00[7:0], \t0.t0.s4.out };
  assign \t0.t0.s0.clk = clk;
  assign \t0.t0.s0.in = state_in[127:120];
  assign \t0.t0.s4.clk = clk;
  assign \t0.t0.s4.in = state_in[127:120];
  assign \t0.t1.clk = clk;
  assign \t0.t1.in = state_in[119:112];
  assign \t0.t1.out = { \t0.t1.s0.out , \t0.t1.s0.out , p01[31:24], \t0.t1.s4.out };
  assign \t0.t1.s0.clk = clk;
  assign \t0.t1.s0.in = state_in[119:112];
  assign \t0.t1.s4.clk = clk;
  assign \t0.t1.s4.in = state_in[119:112];
  assign \t0.t2.clk = clk;
  assign \t0.t2.in = state_in[111:104];
  assign \t0.t2.out = { \t0.t2.s0.out , \t0.t2.s0.out , p02[23:16], \t0.t2.s4.out };
  assign \t0.t2.s0.clk = clk;
  assign \t0.t2.s0.in = state_in[111:104];
  assign \t0.t2.s4.clk = clk;
  assign \t0.t2.s4.in = state_in[111:104];
  assign \t0.t3.clk = clk;
  assign \t0.t3.in = state_in[103:96];
  assign \t0.t3.out = { \t0.t3.s0.out , \t0.t3.s0.out , p03[15:8], \t0.t3.s4.out };
  assign \t0.t3.s0.clk = clk;
  assign \t0.t3.s0.in = state_in[103:96];
  assign \t0.t3.s4.clk = clk;
  assign \t0.t3.s4.in = state_in[103:96];
  assign \t1.b0 = state_in[95:88];
  assign \t1.b1 = state_in[87:80];
  assign \t1.b2 = state_in[79:72];
  assign \t1.b3 = state_in[71:64];
  assign \t1.clk = clk;
  assign \t1.p0 = { \t1.t0.s4.out , \t1.t0.s0.out , \t1.t0.s0.out , p10[7:0] };
  assign \t1.p1 = { p11[31:24], \t1.t1.s4.out , \t1.t1.s0.out , \t1.t1.s0.out };
  assign \t1.p2 = { \t1.t2.s0.out , p12[23:16], \t1.t2.s4.out , \t1.t2.s0.out };
  assign \t1.p3 = { \t1.t3.s0.out , \t1.t3.s0.out , p13[15:8], \t1.t3.s4.out };
  assign \t1.state = state_in[95:64];
  assign \t1.t0.clk = clk;
  assign \t1.t0.in = state_in[95:88];
  assign \t1.t0.out = { \t1.t0.s0.out , \t1.t0.s0.out , p10[7:0], \t1.t0.s4.out };
  assign \t1.t0.s0.clk = clk;
  assign \t1.t0.s0.in = state_in[95:88];
  assign \t1.t0.s4.clk = clk;
  assign \t1.t0.s4.in = state_in[95:88];
  assign \t1.t1.clk = clk;
  assign \t1.t1.in = state_in[87:80];
  assign \t1.t1.out = { \t1.t1.s0.out , \t1.t1.s0.out , p11[31:24], \t1.t1.s4.out };
  assign \t1.t1.s0.clk = clk;
  assign \t1.t1.s0.in = state_in[87:80];
  assign \t1.t1.s4.clk = clk;
  assign \t1.t1.s4.in = state_in[87:80];
  assign \t1.t2.clk = clk;
  assign \t1.t2.in = state_in[79:72];
  assign \t1.t2.out = { \t1.t2.s0.out , \t1.t2.s0.out , p12[23:16], \t1.t2.s4.out };
  assign \t1.t2.s0.clk = clk;
  assign \t1.t2.s0.in = state_in[79:72];
  assign \t1.t2.s4.clk = clk;
  assign \t1.t2.s4.in = state_in[79:72];
  assign \t1.t3.clk = clk;
  assign \t1.t3.in = state_in[71:64];
  assign \t1.t3.out = { \t1.t3.s0.out , \t1.t3.s0.out , p13[15:8], \t1.t3.s4.out };
  assign \t1.t3.s0.clk = clk;
  assign \t1.t3.s0.in = state_in[71:64];
  assign \t1.t3.s4.clk = clk;
  assign \t1.t3.s4.in = state_in[71:64];
  assign \t2.b0 = state_in[63:56];
  assign \t2.b1 = state_in[55:48];
  assign \t2.b2 = state_in[47:40];
  assign \t2.b3 = state_in[39:32];
  assign \t2.clk = clk;
  assign \t2.p0 = { \t2.t0.s4.out , \t2.t0.s0.out , \t2.t0.s0.out , p20[7:0] };
  assign \t2.p1 = { p21[31:24], \t2.t1.s4.out , \t2.t1.s0.out , \t2.t1.s0.out };
  assign \t2.p2 = { \t2.t2.s0.out , p22[23:16], \t2.t2.s4.out , \t2.t2.s0.out };
  assign \t2.p3 = { \t2.t3.s0.out , \t2.t3.s0.out , p23[15:8], \t2.t3.s4.out };
  assign \t2.state = state_in[63:32];
  assign \t2.t0.clk = clk;
  assign \t2.t0.in = state_in[63:56];
  assign \t2.t0.out = { \t2.t0.s0.out , \t2.t0.s0.out , p20[7:0], \t2.t0.s4.out };
  assign \t2.t0.s0.clk = clk;
  assign \t2.t0.s0.in = state_in[63:56];
  assign \t2.t0.s4.clk = clk;
  assign \t2.t0.s4.in = state_in[63:56];
  assign \t2.t1.clk = clk;
  assign \t2.t1.in = state_in[55:48];
  assign \t2.t1.out = { \t2.t1.s0.out , \t2.t1.s0.out , p21[31:24], \t2.t1.s4.out };
  assign \t2.t1.s0.clk = clk;
  assign \t2.t1.s0.in = state_in[55:48];
  assign \t2.t1.s4.clk = clk;
  assign \t2.t1.s4.in = state_in[55:48];
  assign \t2.t2.clk = clk;
  assign \t2.t2.in = state_in[47:40];
  assign \t2.t2.out = { \t2.t2.s0.out , \t2.t2.s0.out , p22[23:16], \t2.t2.s4.out };
  assign \t2.t2.s0.clk = clk;
  assign \t2.t2.s0.in = state_in[47:40];
  assign \t2.t2.s4.clk = clk;
  assign \t2.t2.s4.in = state_in[47:40];
  assign \t2.t3.clk = clk;
  assign \t2.t3.in = state_in[39:32];
  assign \t2.t3.out = { \t2.t3.s0.out , \t2.t3.s0.out , p23[15:8], \t2.t3.s4.out };
  assign \t2.t3.s0.clk = clk;
  assign \t2.t3.s0.in = state_in[39:32];
  assign \t2.t3.s4.clk = clk;
  assign \t2.t3.s4.in = state_in[39:32];
  assign \t3.b0 = state_in[31:24];
  assign \t3.b1 = state_in[23:16];
  assign \t3.b2 = state_in[15:8];
  assign \t3.b3 = state_in[7:0];
  assign \t3.clk = clk;
  assign \t3.p0 = { \t3.t0.s4.out , \t3.t0.s0.out , \t3.t0.s0.out , p30[7:0] };
  assign \t3.p1 = { p31[31:24], \t3.t1.s4.out , \t3.t1.s0.out , \t3.t1.s0.out };
  assign \t3.p2 = { \t3.t2.s0.out , p32[23:16], \t3.t2.s4.out , \t3.t2.s0.out };
  assign \t3.p3 = { \t3.t3.s0.out , \t3.t3.s0.out , p33[15:8], \t3.t3.s4.out };
  assign \t3.state = state_in[31:0];
  assign \t3.t0.clk = clk;
  assign \t3.t0.in = state_in[31:24];
  assign \t3.t0.out = { \t3.t0.s0.out , \t3.t0.s0.out , p30[7:0], \t3.t0.s4.out };
  assign \t3.t0.s0.clk = clk;
  assign \t3.t0.s0.in = state_in[31:24];
  assign \t3.t0.s4.clk = clk;
  assign \t3.t0.s4.in = state_in[31:24];
  assign \t3.t1.clk = clk;
  assign \t3.t1.in = state_in[23:16];
  assign \t3.t1.out = { \t3.t1.s0.out , \t3.t1.s0.out , p31[31:24], \t3.t1.s4.out };
  assign \t3.t1.s0.clk = clk;
  assign \t3.t1.s0.in = state_in[23:16];
  assign \t3.t1.s4.clk = clk;
  assign \t3.t1.s4.in = state_in[23:16];
  assign \t3.t2.clk = clk;
  assign \t3.t2.in = state_in[15:8];
  assign \t3.t2.out = { \t3.t2.s0.out , \t3.t2.s0.out , p32[23:16], \t3.t2.s4.out };
  assign \t3.t2.s0.clk = clk;
  assign \t3.t2.s0.in = state_in[15:8];
  assign \t3.t2.s4.clk = clk;
  assign \t3.t2.s4.in = state_in[15:8];
  assign \t3.t3.clk = clk;
  assign \t3.t3.in = state_in[7:0];
  assign \t3.t3.out = { \t3.t3.s0.out , \t3.t3.s0.out , p33[15:8], \t3.t3.s4.out };
  assign \t3.t3.s0.clk = clk;
  assign \t3.t3.s0.in = state_in[7:0];
  assign \t3.t3.s4.clk = clk;
  assign \t3.t3.s4.in = state_in[7:0];
endmodule
