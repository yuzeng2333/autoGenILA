module \$paramod\SDP_Y_IDX_mgc_in_wire_v1\rscid=3\width=32 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:78" *)
  output [31:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_idx.v:79" *)
  input [31:0] z;
  assign d = z;
endmodule
