module bar__DOT__i1(
__START__,
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
in,
rcon,
out_1,
__COUNTER_start__n0
);
input            __START__;
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg    [127:0] in;
output reg      [7:0] rcon;
output reg    [127:0] out_1;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire            __START__;
wire      [7:0] bv_8_0_n582;
wire      [7:0] bv_8_100_n416;
wire      [7:0] bv_8_101_n260;
wire      [7:0] bv_8_102_n175;
wire      [7:0] bv_8_103_n524;
wire      [7:0] bv_8_104_n38;
wire      [7:0] bv_8_105_n112;
wire      [7:0] bv_8_106_n515;
wire      [7:0] bv_8_107_n512;
wire      [7:0] bv_8_108_n271;
wire      [7:0] bv_8_109_n288;
wire      [7:0] bv_8_10_n342;
wire      [7:0] bv_8_110_n503;
wire      [7:0] bv_8_111_n500;
wire      [7:0] bv_8_112_n187;
wire      [7:0] bv_8_113_n494;
wire      [7:0] bv_8_114_n490;
wire      [7:0] bv_8_115_n407;
wire      [7:0] bv_8_116_n210;
wire      [7:0] bv_8_117_n483;
wire      [7:0] bv_8_118_n479;
wire      [7:0] bv_8_119_n476;
wire      [7:0] bv_8_11_n358;
wire      [7:0] bv_8_120_n242;
wire      [7:0] bv_8_121_n301;
wire      [7:0] bv_8_122_n256;
wire      [7:0] bv_8_123_n466;
wire      [7:0] bv_8_124_n462;
wire      [7:0] bv_8_125_n459;
wire      [7:0] bv_8_126_n422;
wire      [7:0] bv_8_127_n454;
wire      [7:0] bv_8_128_n451;
wire      [7:0] bv_8_129_n400;
wire      [7:0] bv_8_12_n449;
wire      [7:0] bv_8_130_n444;
wire      [7:0] bv_8_131_n441;
wire      [7:0] bv_8_132_n437;
wire      [7:0] bv_8_133_n434;
wire      [7:0] bv_8_134_n141;
wire      [7:0] bv_8_135_n90;
wire      [7:0] bv_8_136_n380;
wire      [7:0] bv_8_137_n58;
wire      [7:0] bv_8_138_n191;
wire      [7:0] bv_8_139_n194;
wire      [7:0] bv_8_13_n54;
wire      [7:0] bv_8_140_n66;
wire      [7:0] bv_8_141_n284;
wire      [7:0] bv_8_142_n104;
wire      [7:0] bv_8_143_n405;
wire      [7:0] bv_8_144_n384;
wire      [7:0] bv_8_145_n311;
wire      [7:0] bv_8_146_n395;
wire      [7:0] bv_8_147_n392;
wire      [7:0] bv_8_148_n101;
wire      [7:0] bv_8_149_n307;
wire      [7:0] bv_8_14_n160;
wire      [7:0] bv_8_150_n382;
wire      [7:0] bv_8_151_n378;
wire      [7:0] bv_8_152_n120;
wire      [7:0] bv_8_153_n30;
wire      [7:0] bv_8_154_n370;
wire      [7:0] bv_8_155_n97;
wire      [7:0] bv_8_156_n364;
wire      [7:0] bv_8_157_n360;
wire      [7:0] bv_8_158_n129;
wire      [7:0] bv_8_159_n354;
wire      [7:0] bv_8_15_n22;
wire      [7:0] bv_8_160_n351;
wire      [7:0] bv_8_161_n62;
wire      [7:0] bv_8_162_n344;
wire      [7:0] bv_8_163_n340;
wire      [7:0] bv_8_164_n336;
wire      [7:0] bv_8_165_n332;
wire      [7:0] bv_8_166_n227;
wire      [7:0] bv_8_167_n325;
wire      [7:0] bv_8_168_n322;
wire      [7:0] bv_8_169_n275;
wire      [7:0] bv_8_16_n464;
wire      [7:0] bv_8_170_n317;
wire      [7:0] bv_8_171_n313;
wire      [7:0] bv_8_172_n309;
wire      [7:0] bv_8_173_n305;
wire      [7:0] bv_8_174_n253;
wire      [7:0] bv_8_175_n299;
wire      [7:0] bv_8_176_n18;
wire      [7:0] bv_8_177_n294;
wire      [7:0] bv_8_178_n290;
wire      [7:0] bv_8_179_n286;
wire      [7:0] bv_8_17_n116;
wire      [7:0] bv_8_180_n223;
wire      [7:0] bv_8_181_n179;
wire      [7:0] bv_8_182_n277;
wire      [7:0] bv_8_183_n273;
wire      [7:0] bv_8_184_n269;
wire      [7:0] bv_8_185_n145;
wire      [7:0] bv_8_186_n246;
wire      [7:0] bv_8_187_n10;
wire      [7:0] bv_8_188_n258;
wire      [7:0] bv_8_189_n198;
wire      [7:0] bv_8_18_n643;
wire      [7:0] bv_8_190_n251;
wire      [7:0] bv_8_191_n50;
wire      [7:0] bv_8_192_n244;
wire      [7:0] bv_8_193_n137;
wire      [7:0] bv_8_194_n237;
wire      [7:0] bv_8_195_n233;
wire      [7:0] bv_8_196_n229;
wire      [7:0] bv_8_197_n225;
wire      [7:0] bv_8_198_n220;
wire      [7:0] bv_8_199_n218;
wire      [7:0] bv_8_19_n446;
wire      [7:0] bv_8_1_n752;
wire      [7:0] bv_8_200_n215;
wire      [7:0] bv_8_201_n212;
wire      [7:0] bv_8_202_n208;
wire      [7:0] bv_8_203_n204;
wire      [7:0] bv_8_204_n200;
wire      [7:0] bv_8_205_n196;
wire      [7:0] bv_8_206_n82;
wire      [7:0] bv_8_207_n189;
wire      [7:0] bv_8_208_n185;
wire      [7:0] bv_8_209_n181;
wire      [7:0] bv_8_20_n368;
wire      [7:0] bv_8_210_n177;
wire      [7:0] bv_8_211_n173;
wire      [7:0] bv_8_212_n169;
wire      [7:0] bv_8_213_n165;
wire      [7:0] bv_8_214_n162;
wire      [7:0] bv_8_215_n158;
wire      [7:0] bv_8_216_n154;
wire      [7:0] bv_8_217_n108;
wire      [7:0] bv_8_218_n147;
wire      [7:0] bv_8_219_n143;
wire      [7:0] bv_8_21_n673;
wire      [7:0] bv_8_220_n139;
wire      [7:0] bv_8_221_n135;
wire      [7:0] bv_8_222_n131;
wire      [7:0] bv_8_223_n70;
wire      [7:0] bv_8_224_n125;
wire      [7:0] bv_8_225_n122;
wire      [7:0] bv_8_226_n118;
wire      [7:0] bv_8_227_n114;
wire      [7:0] bv_8_228_n110;
wire      [7:0] bv_8_229_n106;
wire      [7:0] bv_8_22_n6;
wire      [7:0] bv_8_230_n46;
wire      [7:0] bv_8_231_n99;
wire      [7:0] bv_8_232_n95;
wire      [7:0] bv_8_233_n86;
wire      [7:0] bv_8_234_n88;
wire      [7:0] bv_8_235_n84;
wire      [7:0] bv_8_236_n80;
wire      [7:0] bv_8_237_n76;
wire      [7:0] bv_8_238_n72;
wire      [7:0] bv_8_239_n68;
wire      [7:0] bv_8_23_n429;
wire      [7:0] bv_8_240_n64;
wire      [7:0] bv_8_241_n60;
wire      [7:0] bv_8_242_n56;
wire      [7:0] bv_8_243_n52;
wire      [7:0] bv_8_244_n48;
wire      [7:0] bv_8_245_n44;
wire      [7:0] bv_8_246_n40;
wire      [7:0] bv_8_247_n36;
wire      [7:0] bv_8_248_n32;
wire      [7:0] bv_8_249_n28;
wire      [7:0] bv_8_24_n658;
wire      [7:0] bv_8_250_n24;
wire      [7:0] bv_8_251_n20;
wire      [7:0] bv_8_252_n16;
wire      [7:0] bv_8_253_n12;
wire      [7:0] bv_8_254_n8;
wire      [7:0] bv_8_255_n4;
wire      [7:0] bv_8_25_n410;
wire      [7:0] bv_8_26_n618;
wire      [7:0] bv_8_27_n615;
wire      [7:0] bv_8_28_n231;
wire      [7:0] bv_8_29_n133;
wire      [7:0] bv_8_2_n517;
wire      [7:0] bv_8_30_n93;
wire      [7:0] bv_8_31_n206;
wire      [7:0] bv_8_32_n575;
wire      [7:0] bv_8_33_n468;
wire      [7:0] bv_8_34_n390;
wire      [7:0] bv_8_35_n663;
wire      [7:0] bv_8_36_n330;
wire      [7:0] bv_8_37_n239;
wire      [7:0] bv_8_38_n692;
wire      [7:0] bv_8_39_n634;
wire      [7:0] bv_8_3_n167;
wire      [7:0] bv_8_40_n74;
wire      [7:0] bv_8_41_n596;
wire      [7:0] bv_8_42_n387;
wire      [7:0] bv_8_43_n681;
wire      [7:0] bv_8_44_n621;
wire      [7:0] bv_8_45_n26;
wire      [7:0] bv_8_46_n235;
wire      [7:0] bv_8_47_n591;
wire      [7:0] bv_8_48_n668;
wire      [7:0] bv_8_49_n665;
wire      [7:0] bv_8_4_n670;
wire      [7:0] bv_8_50_n349;
wire      [7:0] bv_8_51_n528;
wire      [7:0] bv_8_52_n656;
wire      [7:0] bv_8_53_n152;
wire      [7:0] bv_8_54_n650;
wire      [7:0] bv_8_55_n292;
wire      [7:0] bv_8_56_n481;
wire      [7:0] bv_8_57_n558;
wire      [7:0] bv_8_58_n346;
wire      [7:0] bv_8_59_n603;
wire      [7:0] bv_8_5_n652;
wire      [7:0] bv_8_60_n507;
wire      [7:0] bv_8_61_n419;
wire      [7:0] bv_8_62_n183;
wire      [7:0] bv_8_63_n628;
wire      [7:0] bv_8_64_n492;
wire      [7:0] bv_8_65_n34;
wire      [7:0] bv_8_66_n42;
wire      [7:0] bv_8_67_n534;
wire      [7:0] bv_8_68_n432;
wire      [7:0] bv_8_69_n522;
wire      [7:0] bv_8_6_n334;
wire      [7:0] bv_8_70_n376;
wire      [7:0] bv_8_71_n607;
wire      [7:0] bv_8_72_n171;
wire      [7:0] bv_8_73_n338;
wire      [7:0] bv_8_74_n554;
wire      [7:0] bv_8_75_n202;
wire      [7:0] bv_8_76_n551;
wire      [7:0] bv_8_77_n531;
wire      [7:0] bv_8_78_n279;
wire      [7:0] bv_8_79_n397;
wire      [7:0] bv_8_7_n646;
wire      [7:0] bv_8_80_n510;
wire      [7:0] bv_8_81_n498;
wire      [7:0] bv_8_82_n580;
wire      [7:0] bv_8_83_n577;
wire      [7:0] bv_8_84_n14;
wire      [7:0] bv_8_85_n78;
wire      [7:0] bv_8_86_n267;
wire      [7:0] bv_8_87_n149;
wire      [7:0] bv_8_88_n548;
wire      [7:0] bv_8_89_n563;
wire      [7:0] bv_8_8_n249;
wire      [7:0] bv_8_90_n560;
wire      [7:0] bv_8_91_n556;
wire      [7:0] bv_8_92_n327;
wire      [7:0] bv_8_93_n413;
wire      [7:0] bv_8_94_n362;
wire      [7:0] bv_8_95_n439;
wire      [7:0] bv_8_96_n403;
wire      [7:0] bv_8_97_n156;
wire      [7:0] bv_8_98_n315;
wire      [7:0] bv_8_99_n536;
wire      [7:0] bv_8_9_n626;
wire            clk;
(* keep *) wire    [127:0] in_randinit;
wire      [7:0] n1;
wire            n100;
wire      [7:0] n1000;
wire      [7:0] n1001;
wire      [7:0] n1002;
wire      [7:0] n1003;
wire      [7:0] n1004;
wire      [7:0] n1005;
wire      [7:0] n1006;
wire      [7:0] n1007;
wire      [7:0] n1008;
wire      [7:0] n1009;
wire      [7:0] n1010;
wire      [7:0] n1011;
wire      [7:0] n1012;
wire      [7:0] n1013;
wire      [7:0] n1014;
wire      [7:0] n1015;
wire      [7:0] n1016;
wire      [7:0] n1017;
wire      [7:0] n1018;
wire      [7:0] n1019;
wire      [7:0] n102;
wire      [7:0] n1020;
wire      [7:0] n1021;
wire      [7:0] n1022;
wire      [7:0] n1023;
wire      [7:0] n1024;
wire      [7:0] n1025;
wire      [7:0] n1026;
wire      [7:0] n1027;
wire      [7:0] n1028;
wire      [7:0] n1029;
wire            n103;
wire            n1030;
wire      [7:0] n1031;
wire            n1032;
wire      [7:0] n1033;
wire            n1034;
wire      [7:0] n1035;
wire            n1036;
wire      [7:0] n1037;
wire            n1038;
wire      [7:0] n1039;
wire            n1040;
wire      [7:0] n1041;
wire            n1042;
wire      [7:0] n1043;
wire            n1044;
wire      [7:0] n1045;
wire            n1046;
wire      [7:0] n1047;
wire            n1048;
wire      [7:0] n1049;
wire      [7:0] n105;
wire            n1050;
wire      [7:0] n1051;
wire            n1052;
wire      [7:0] n1053;
wire            n1054;
wire      [7:0] n1055;
wire            n1056;
wire      [7:0] n1057;
wire            n1058;
wire      [7:0] n1059;
wire            n1060;
wire      [7:0] n1061;
wire            n1062;
wire      [7:0] n1063;
wire            n1064;
wire      [7:0] n1065;
wire            n1066;
wire      [7:0] n1067;
wire            n1068;
wire      [7:0] n1069;
wire            n107;
wire            n1070;
wire      [7:0] n1071;
wire            n1072;
wire      [7:0] n1073;
wire            n1074;
wire      [7:0] n1075;
wire            n1076;
wire      [7:0] n1077;
wire            n1078;
wire      [7:0] n1079;
wire            n1080;
wire      [7:0] n1081;
wire            n1082;
wire      [7:0] n1083;
wire            n1084;
wire      [7:0] n1085;
wire            n1086;
wire      [7:0] n1087;
wire            n1088;
wire      [7:0] n1089;
wire      [7:0] n109;
wire            n1090;
wire      [7:0] n1091;
wire            n1092;
wire      [7:0] n1093;
wire            n1094;
wire      [7:0] n1095;
wire            n1096;
wire      [7:0] n1097;
wire            n1098;
wire      [7:0] n1099;
wire      [7:0] n11;
wire            n1100;
wire      [7:0] n1101;
wire            n1102;
wire      [7:0] n1103;
wire            n1104;
wire      [7:0] n1105;
wire            n1106;
wire      [7:0] n1107;
wire            n1108;
wire      [7:0] n1109;
wire            n111;
wire            n1110;
wire      [7:0] n1111;
wire            n1112;
wire      [7:0] n1113;
wire            n1114;
wire      [7:0] n1115;
wire            n1116;
wire      [7:0] n1117;
wire            n1118;
wire      [7:0] n1119;
wire            n1120;
wire      [7:0] n1121;
wire            n1122;
wire      [7:0] n1123;
wire            n1124;
wire      [7:0] n1125;
wire            n1126;
wire      [7:0] n1127;
wire            n1128;
wire      [7:0] n1129;
wire      [7:0] n113;
wire            n1130;
wire      [7:0] n1131;
wire            n1132;
wire      [7:0] n1133;
wire            n1134;
wire      [7:0] n1135;
wire            n1136;
wire      [7:0] n1137;
wire            n1138;
wire      [7:0] n1139;
wire            n1140;
wire      [7:0] n1141;
wire            n1142;
wire      [7:0] n1143;
wire            n1144;
wire      [7:0] n1145;
wire            n1146;
wire      [7:0] n1147;
wire            n1148;
wire      [7:0] n1149;
wire            n115;
wire            n1150;
wire      [7:0] n1151;
wire            n1152;
wire      [7:0] n1153;
wire            n1154;
wire      [7:0] n1155;
wire            n1156;
wire      [7:0] n1157;
wire            n1158;
wire      [7:0] n1159;
wire            n1160;
wire      [7:0] n1161;
wire            n1162;
wire      [7:0] n1163;
wire            n1164;
wire      [7:0] n1165;
wire            n1166;
wire      [7:0] n1167;
wire            n1168;
wire      [7:0] n1169;
wire      [7:0] n117;
wire            n1170;
wire      [7:0] n1171;
wire            n1172;
wire      [7:0] n1173;
wire            n1174;
wire      [7:0] n1175;
wire            n1176;
wire      [7:0] n1177;
wire            n1178;
wire      [7:0] n1179;
wire            n1180;
wire      [7:0] n1181;
wire            n1182;
wire      [7:0] n1183;
wire            n1184;
wire      [7:0] n1185;
wire            n1186;
wire      [7:0] n1187;
wire            n1188;
wire      [7:0] n1189;
wire            n119;
wire            n1190;
wire      [7:0] n1191;
wire            n1192;
wire      [7:0] n1193;
wire            n1194;
wire      [7:0] n1195;
wire            n1196;
wire      [7:0] n1197;
wire            n1198;
wire      [7:0] n1199;
wire            n1200;
wire      [7:0] n1201;
wire            n1202;
wire      [7:0] n1203;
wire            n1204;
wire      [7:0] n1205;
wire            n1206;
wire      [7:0] n1207;
wire            n1208;
wire      [7:0] n1209;
wire      [7:0] n121;
wire            n1210;
wire      [7:0] n1211;
wire            n1212;
wire      [7:0] n1213;
wire            n1214;
wire      [7:0] n1215;
wire            n1216;
wire      [7:0] n1217;
wire            n1218;
wire      [7:0] n1219;
wire            n1220;
wire      [7:0] n1221;
wire            n1222;
wire      [7:0] n1223;
wire            n1224;
wire      [7:0] n1225;
wire            n1226;
wire      [7:0] n1227;
wire            n1228;
wire      [7:0] n1229;
wire            n123;
wire            n1230;
wire      [7:0] n1231;
wire            n1232;
wire      [7:0] n1233;
wire            n1234;
wire      [7:0] n1235;
wire            n1236;
wire      [7:0] n1237;
wire            n1238;
wire      [7:0] n1239;
wire      [7:0] n124;
wire            n1240;
wire      [7:0] n1241;
wire            n1242;
wire      [7:0] n1243;
wire            n1244;
wire      [7:0] n1245;
wire            n1246;
wire      [7:0] n1247;
wire            n1248;
wire      [7:0] n1249;
wire            n1250;
wire      [7:0] n1251;
wire            n1252;
wire      [7:0] n1253;
wire            n1254;
wire      [7:0] n1255;
wire            n1256;
wire      [7:0] n1257;
wire            n1258;
wire      [7:0] n1259;
wire            n126;
wire            n1260;
wire      [7:0] n1261;
wire            n1262;
wire      [7:0] n1263;
wire            n1264;
wire      [7:0] n1265;
wire            n1266;
wire      [7:0] n1267;
wire            n1268;
wire      [7:0] n1269;
wire      [7:0] n127;
wire            n1270;
wire      [7:0] n1271;
wire            n1272;
wire      [7:0] n1273;
wire            n1274;
wire      [7:0] n1275;
wire            n1276;
wire      [7:0] n1277;
wire            n1278;
wire      [7:0] n1279;
wire            n128;
wire            n1280;
wire      [7:0] n1281;
wire            n1282;
wire      [7:0] n1283;
wire            n1284;
wire      [7:0] n1285;
wire            n1286;
wire      [7:0] n1287;
wire            n1288;
wire      [7:0] n1289;
wire            n1290;
wire      [7:0] n1291;
wire            n1292;
wire      [7:0] n1293;
wire            n1294;
wire      [7:0] n1295;
wire            n1296;
wire      [7:0] n1297;
wire            n1298;
wire      [7:0] n1299;
wire            n13;
wire      [7:0] n130;
wire            n1300;
wire      [7:0] n1301;
wire            n1302;
wire      [7:0] n1303;
wire            n1304;
wire      [7:0] n1305;
wire            n1306;
wire      [7:0] n1307;
wire            n1308;
wire      [7:0] n1309;
wire            n1310;
wire      [7:0] n1311;
wire            n1312;
wire      [7:0] n1313;
wire            n1314;
wire      [7:0] n1315;
wire            n1316;
wire      [7:0] n1317;
wire            n1318;
wire      [7:0] n1319;
wire            n132;
wire            n1320;
wire      [7:0] n1321;
wire            n1322;
wire      [7:0] n1323;
wire            n1324;
wire      [7:0] n1325;
wire            n1326;
wire      [7:0] n1327;
wire            n1328;
wire      [7:0] n1329;
wire            n1330;
wire      [7:0] n1331;
wire            n1332;
wire      [7:0] n1333;
wire            n1334;
wire      [7:0] n1335;
wire            n1336;
wire      [7:0] n1337;
wire            n1338;
wire      [7:0] n1339;
wire      [7:0] n134;
wire            n1340;
wire      [7:0] n1341;
wire            n1342;
wire      [7:0] n1343;
wire            n1344;
wire      [7:0] n1345;
wire            n1346;
wire      [7:0] n1347;
wire            n1348;
wire      [7:0] n1349;
wire            n1350;
wire      [7:0] n1351;
wire            n1352;
wire      [7:0] n1353;
wire            n1354;
wire      [7:0] n1355;
wire            n1356;
wire      [7:0] n1357;
wire            n1358;
wire      [7:0] n1359;
wire            n136;
wire            n1360;
wire      [7:0] n1361;
wire            n1362;
wire      [7:0] n1363;
wire            n1364;
wire      [7:0] n1365;
wire            n1366;
wire      [7:0] n1367;
wire            n1368;
wire      [7:0] n1369;
wire            n1370;
wire      [7:0] n1371;
wire            n1372;
wire      [7:0] n1373;
wire            n1374;
wire      [7:0] n1375;
wire            n1376;
wire      [7:0] n1377;
wire            n1378;
wire      [7:0] n1379;
wire      [7:0] n138;
wire            n1380;
wire      [7:0] n1381;
wire            n1382;
wire      [7:0] n1383;
wire            n1384;
wire      [7:0] n1385;
wire            n1386;
wire      [7:0] n1387;
wire            n1388;
wire      [7:0] n1389;
wire            n1390;
wire      [7:0] n1391;
wire            n1392;
wire      [7:0] n1393;
wire            n1394;
wire      [7:0] n1395;
wire            n1396;
wire      [7:0] n1397;
wire            n1398;
wire      [7:0] n1399;
wire            n140;
wire            n1400;
wire      [7:0] n1401;
wire            n1402;
wire      [7:0] n1403;
wire            n1404;
wire      [7:0] n1405;
wire            n1406;
wire      [7:0] n1407;
wire            n1408;
wire      [7:0] n1409;
wire            n1410;
wire      [7:0] n1411;
wire            n1412;
wire      [7:0] n1413;
wire            n1414;
wire      [7:0] n1415;
wire            n1416;
wire      [7:0] n1417;
wire            n1418;
wire      [7:0] n1419;
wire      [7:0] n142;
wire            n1420;
wire      [7:0] n1421;
wire            n1422;
wire      [7:0] n1423;
wire            n1424;
wire      [7:0] n1425;
wire            n1426;
wire      [7:0] n1427;
wire            n1428;
wire      [7:0] n1429;
wire            n1430;
wire      [7:0] n1431;
wire            n1432;
wire      [7:0] n1433;
wire            n1434;
wire      [7:0] n1435;
wire            n1436;
wire      [7:0] n1437;
wire            n1438;
wire      [7:0] n1439;
wire            n144;
wire            n1440;
wire      [7:0] n1441;
wire            n1442;
wire      [7:0] n1443;
wire            n1444;
wire      [7:0] n1445;
wire            n1446;
wire      [7:0] n1447;
wire            n1448;
wire      [7:0] n1449;
wire            n1450;
wire      [7:0] n1451;
wire            n1452;
wire      [7:0] n1453;
wire            n1454;
wire      [7:0] n1455;
wire            n1456;
wire      [7:0] n1457;
wire            n1458;
wire      [7:0] n1459;
wire      [7:0] n146;
wire            n1460;
wire      [7:0] n1461;
wire            n1462;
wire      [7:0] n1463;
wire            n1464;
wire      [7:0] n1465;
wire            n1466;
wire      [7:0] n1467;
wire            n1468;
wire      [7:0] n1469;
wire            n1470;
wire      [7:0] n1471;
wire            n1472;
wire      [7:0] n1473;
wire            n1474;
wire      [7:0] n1475;
wire            n1476;
wire      [7:0] n1477;
wire            n1478;
wire      [7:0] n1479;
wire            n148;
wire            n1480;
wire      [7:0] n1481;
wire            n1482;
wire      [7:0] n1483;
wire            n1484;
wire      [7:0] n1485;
wire            n1486;
wire      [7:0] n1487;
wire            n1488;
wire      [7:0] n1489;
wire            n1490;
wire      [7:0] n1491;
wire            n1492;
wire      [7:0] n1493;
wire            n1494;
wire      [7:0] n1495;
wire            n1496;
wire      [7:0] n1497;
wire            n1498;
wire      [7:0] n1499;
wire      [7:0] n15;
wire      [7:0] n150;
wire            n1500;
wire      [7:0] n1501;
wire            n1502;
wire      [7:0] n1503;
wire            n1504;
wire      [7:0] n1505;
wire            n1506;
wire      [7:0] n1507;
wire            n1508;
wire      [7:0] n1509;
wire            n151;
wire            n1510;
wire      [7:0] n1511;
wire            n1512;
wire      [7:0] n1513;
wire            n1514;
wire      [7:0] n1515;
wire            n1516;
wire      [7:0] n1517;
wire            n1518;
wire      [7:0] n1519;
wire            n1520;
wire      [7:0] n1521;
wire            n1522;
wire      [7:0] n1523;
wire            n1524;
wire      [7:0] n1525;
wire            n1526;
wire      [7:0] n1527;
wire            n1528;
wire      [7:0] n1529;
wire      [7:0] n153;
wire            n1530;
wire      [7:0] n1531;
wire            n1532;
wire      [7:0] n1533;
wire            n1534;
wire      [7:0] n1535;
wire            n1536;
wire      [7:0] n1537;
wire            n1538;
wire      [7:0] n1539;
wire            n1540;
wire      [7:0] n1541;
wire      [7:0] n1542;
wire      [7:0] n1543;
wire      [7:0] n1544;
wire      [7:0] n1545;
wire      [7:0] n1546;
wire      [7:0] n1547;
wire      [7:0] n1548;
wire      [7:0] n1549;
wire            n155;
wire      [7:0] n1550;
wire      [7:0] n1551;
wire      [7:0] n1552;
wire      [7:0] n1553;
wire      [7:0] n1554;
wire      [7:0] n1555;
wire      [7:0] n1556;
wire      [7:0] n1557;
wire      [7:0] n1558;
wire      [7:0] n1559;
wire      [7:0] n1560;
wire      [7:0] n1561;
wire      [7:0] n1562;
wire      [7:0] n1563;
wire      [7:0] n1564;
wire      [7:0] n1565;
wire      [7:0] n1566;
wire      [7:0] n1567;
wire      [7:0] n1568;
wire      [7:0] n1569;
wire      [7:0] n157;
wire      [7:0] n1570;
wire      [7:0] n1571;
wire      [7:0] n1572;
wire      [7:0] n1573;
wire      [7:0] n1574;
wire      [7:0] n1575;
wire      [7:0] n1576;
wire      [7:0] n1577;
wire      [7:0] n1578;
wire      [7:0] n1579;
wire      [7:0] n1580;
wire      [7:0] n1581;
wire      [7:0] n1582;
wire      [7:0] n1583;
wire      [7:0] n1584;
wire      [7:0] n1585;
wire      [7:0] n1586;
wire      [7:0] n1587;
wire      [7:0] n1588;
wire      [7:0] n1589;
wire            n159;
wire      [7:0] n1590;
wire      [7:0] n1591;
wire      [7:0] n1592;
wire      [7:0] n1593;
wire      [7:0] n1594;
wire      [7:0] n1595;
wire      [7:0] n1596;
wire      [7:0] n1597;
wire      [7:0] n1598;
wire      [7:0] n1599;
wire      [7:0] n1600;
wire      [7:0] n1601;
wire      [7:0] n1602;
wire      [7:0] n1603;
wire      [7:0] n1604;
wire      [7:0] n1605;
wire      [7:0] n1606;
wire      [7:0] n1607;
wire      [7:0] n1608;
wire      [7:0] n1609;
wire      [7:0] n161;
wire      [7:0] n1610;
wire      [7:0] n1611;
wire      [7:0] n1612;
wire      [7:0] n1613;
wire      [7:0] n1614;
wire      [7:0] n1615;
wire      [7:0] n1616;
wire      [7:0] n1617;
wire      [7:0] n1618;
wire      [7:0] n1619;
wire      [7:0] n1620;
wire      [7:0] n1621;
wire      [7:0] n1622;
wire      [7:0] n1623;
wire      [7:0] n1624;
wire      [7:0] n1625;
wire      [7:0] n1626;
wire      [7:0] n1627;
wire      [7:0] n1628;
wire      [7:0] n1629;
wire            n163;
wire      [7:0] n1630;
wire      [7:0] n1631;
wire      [7:0] n1632;
wire      [7:0] n1633;
wire      [7:0] n1634;
wire      [7:0] n1635;
wire      [7:0] n1636;
wire      [7:0] n1637;
wire      [7:0] n1638;
wire      [7:0] n1639;
wire      [7:0] n164;
wire      [7:0] n1640;
wire      [7:0] n1641;
wire      [7:0] n1642;
wire      [7:0] n1643;
wire      [7:0] n1644;
wire      [7:0] n1645;
wire      [7:0] n1646;
wire      [7:0] n1647;
wire      [7:0] n1648;
wire      [7:0] n1649;
wire      [7:0] n1650;
wire      [7:0] n1651;
wire      [7:0] n1652;
wire      [7:0] n1653;
wire      [7:0] n1654;
wire      [7:0] n1655;
wire      [7:0] n1656;
wire      [7:0] n1657;
wire      [7:0] n1658;
wire      [7:0] n1659;
wire            n166;
wire      [7:0] n1660;
wire      [7:0] n1661;
wire      [7:0] n1662;
wire      [7:0] n1663;
wire      [7:0] n1664;
wire      [7:0] n1665;
wire      [7:0] n1666;
wire      [7:0] n1667;
wire      [7:0] n1668;
wire      [7:0] n1669;
wire      [7:0] n1670;
wire      [7:0] n1671;
wire      [7:0] n1672;
wire      [7:0] n1673;
wire      [7:0] n1674;
wire      [7:0] n1675;
wire      [7:0] n1676;
wire      [7:0] n1677;
wire      [7:0] n1678;
wire      [7:0] n1679;
wire      [7:0] n168;
wire      [7:0] n1680;
wire      [7:0] n1681;
wire      [7:0] n1682;
wire      [7:0] n1683;
wire      [7:0] n1684;
wire      [7:0] n1685;
wire      [7:0] n1686;
wire      [7:0] n1687;
wire      [7:0] n1688;
wire      [7:0] n1689;
wire      [7:0] n1690;
wire      [7:0] n1691;
wire      [7:0] n1692;
wire      [7:0] n1693;
wire      [7:0] n1694;
wire      [7:0] n1695;
wire      [7:0] n1696;
wire      [7:0] n1697;
wire      [7:0] n1698;
wire      [7:0] n1699;
wire            n17;
wire            n170;
wire      [7:0] n1700;
wire      [7:0] n1701;
wire      [7:0] n1702;
wire      [7:0] n1703;
wire      [7:0] n1704;
wire      [7:0] n1705;
wire      [7:0] n1706;
wire      [7:0] n1707;
wire      [7:0] n1708;
wire      [7:0] n1709;
wire      [7:0] n1710;
wire      [7:0] n1711;
wire      [7:0] n1712;
wire      [7:0] n1713;
wire      [7:0] n1714;
wire      [7:0] n1715;
wire      [7:0] n1716;
wire      [7:0] n1717;
wire      [7:0] n1718;
wire      [7:0] n1719;
wire      [7:0] n172;
wire      [7:0] n1720;
wire      [7:0] n1721;
wire      [7:0] n1722;
wire      [7:0] n1723;
wire      [7:0] n1724;
wire      [7:0] n1725;
wire      [7:0] n1726;
wire      [7:0] n1727;
wire      [7:0] n1728;
wire      [7:0] n1729;
wire      [7:0] n1730;
wire      [7:0] n1731;
wire      [7:0] n1732;
wire      [7:0] n1733;
wire      [7:0] n1734;
wire      [7:0] n1735;
wire      [7:0] n1736;
wire      [7:0] n1737;
wire      [7:0] n1738;
wire      [7:0] n1739;
wire            n174;
wire      [7:0] n1740;
wire      [7:0] n1741;
wire      [7:0] n1742;
wire      [7:0] n1743;
wire      [7:0] n1744;
wire      [7:0] n1745;
wire      [7:0] n1746;
wire      [7:0] n1747;
wire      [7:0] n1748;
wire      [7:0] n1749;
wire      [7:0] n1750;
wire      [7:0] n1751;
wire      [7:0] n1752;
wire      [7:0] n1753;
wire      [7:0] n1754;
wire      [7:0] n1755;
wire      [7:0] n1756;
wire      [7:0] n1757;
wire      [7:0] n1758;
wire      [7:0] n1759;
wire      [7:0] n176;
wire      [7:0] n1760;
wire      [7:0] n1761;
wire      [7:0] n1762;
wire      [7:0] n1763;
wire      [7:0] n1764;
wire      [7:0] n1765;
wire      [7:0] n1766;
wire      [7:0] n1767;
wire      [7:0] n1768;
wire      [7:0] n1769;
wire      [7:0] n1770;
wire      [7:0] n1771;
wire      [7:0] n1772;
wire      [7:0] n1773;
wire      [7:0] n1774;
wire      [7:0] n1775;
wire      [7:0] n1776;
wire      [7:0] n1777;
wire      [7:0] n1778;
wire      [7:0] n1779;
wire            n178;
wire      [7:0] n1780;
wire      [7:0] n1781;
wire      [7:0] n1782;
wire      [7:0] n1783;
wire      [7:0] n1784;
wire      [7:0] n1785;
wire      [7:0] n1786;
wire      [7:0] n1787;
wire      [7:0] n1788;
wire      [7:0] n1789;
wire      [7:0] n1790;
wire      [7:0] n1791;
wire      [7:0] n1792;
wire      [7:0] n1793;
wire      [7:0] n1794;
wire      [7:0] n1795;
wire      [7:0] n1796;
wire      [7:0] n1797;
wire     [15:0] n1798;
wire      [7:0] n1799;
wire      [7:0] n180;
wire      [7:0] n1800;
wire            n1801;
wire      [7:0] n1802;
wire            n1803;
wire      [7:0] n1804;
wire            n1805;
wire      [7:0] n1806;
wire            n1807;
wire      [7:0] n1808;
wire            n1809;
wire      [7:0] n1810;
wire            n1811;
wire      [7:0] n1812;
wire            n1813;
wire      [7:0] n1814;
wire            n1815;
wire      [7:0] n1816;
wire            n1817;
wire      [7:0] n1818;
wire            n1819;
wire            n182;
wire      [7:0] n1820;
wire            n1821;
wire      [7:0] n1822;
wire            n1823;
wire      [7:0] n1824;
wire            n1825;
wire      [7:0] n1826;
wire            n1827;
wire      [7:0] n1828;
wire            n1829;
wire      [7:0] n1830;
wire            n1831;
wire      [7:0] n1832;
wire            n1833;
wire      [7:0] n1834;
wire            n1835;
wire      [7:0] n1836;
wire            n1837;
wire      [7:0] n1838;
wire            n1839;
wire      [7:0] n184;
wire      [7:0] n1840;
wire            n1841;
wire      [7:0] n1842;
wire            n1843;
wire      [7:0] n1844;
wire            n1845;
wire      [7:0] n1846;
wire            n1847;
wire      [7:0] n1848;
wire            n1849;
wire      [7:0] n1850;
wire            n1851;
wire      [7:0] n1852;
wire            n1853;
wire      [7:0] n1854;
wire            n1855;
wire      [7:0] n1856;
wire            n1857;
wire      [7:0] n1858;
wire            n1859;
wire            n186;
wire      [7:0] n1860;
wire            n1861;
wire      [7:0] n1862;
wire            n1863;
wire      [7:0] n1864;
wire            n1865;
wire      [7:0] n1866;
wire            n1867;
wire      [7:0] n1868;
wire            n1869;
wire      [7:0] n1870;
wire            n1871;
wire      [7:0] n1872;
wire            n1873;
wire      [7:0] n1874;
wire            n1875;
wire      [7:0] n1876;
wire            n1877;
wire      [7:0] n1878;
wire            n1879;
wire      [7:0] n188;
wire      [7:0] n1880;
wire            n1881;
wire      [7:0] n1882;
wire            n1883;
wire      [7:0] n1884;
wire            n1885;
wire      [7:0] n1886;
wire            n1887;
wire      [7:0] n1888;
wire            n1889;
wire      [7:0] n1890;
wire            n1891;
wire      [7:0] n1892;
wire            n1893;
wire      [7:0] n1894;
wire            n1895;
wire      [7:0] n1896;
wire            n1897;
wire      [7:0] n1898;
wire            n1899;
wire      [7:0] n19;
wire            n190;
wire      [7:0] n1900;
wire            n1901;
wire      [7:0] n1902;
wire            n1903;
wire      [7:0] n1904;
wire            n1905;
wire      [7:0] n1906;
wire            n1907;
wire      [7:0] n1908;
wire            n1909;
wire      [7:0] n1910;
wire            n1911;
wire      [7:0] n1912;
wire            n1913;
wire      [7:0] n1914;
wire            n1915;
wire      [7:0] n1916;
wire            n1917;
wire      [7:0] n1918;
wire            n1919;
wire      [7:0] n192;
wire      [7:0] n1920;
wire            n1921;
wire      [7:0] n1922;
wire            n1923;
wire      [7:0] n1924;
wire            n1925;
wire      [7:0] n1926;
wire            n1927;
wire      [7:0] n1928;
wire            n1929;
wire            n193;
wire      [7:0] n1930;
wire            n1931;
wire      [7:0] n1932;
wire            n1933;
wire      [7:0] n1934;
wire            n1935;
wire      [7:0] n1936;
wire            n1937;
wire      [7:0] n1938;
wire            n1939;
wire      [7:0] n1940;
wire            n1941;
wire      [7:0] n1942;
wire            n1943;
wire      [7:0] n1944;
wire            n1945;
wire      [7:0] n1946;
wire            n1947;
wire      [7:0] n1948;
wire            n1949;
wire      [7:0] n195;
wire      [7:0] n1950;
wire            n1951;
wire      [7:0] n1952;
wire            n1953;
wire      [7:0] n1954;
wire            n1955;
wire      [7:0] n1956;
wire            n1957;
wire      [7:0] n1958;
wire            n1959;
wire      [7:0] n1960;
wire            n1961;
wire      [7:0] n1962;
wire            n1963;
wire      [7:0] n1964;
wire            n1965;
wire      [7:0] n1966;
wire            n1967;
wire      [7:0] n1968;
wire            n1969;
wire            n197;
wire      [7:0] n1970;
wire            n1971;
wire      [7:0] n1972;
wire            n1973;
wire      [7:0] n1974;
wire            n1975;
wire      [7:0] n1976;
wire            n1977;
wire      [7:0] n1978;
wire            n1979;
wire      [7:0] n1980;
wire            n1981;
wire      [7:0] n1982;
wire            n1983;
wire      [7:0] n1984;
wire            n1985;
wire      [7:0] n1986;
wire            n1987;
wire      [7:0] n1988;
wire            n1989;
wire      [7:0] n199;
wire      [7:0] n1990;
wire            n1991;
wire      [7:0] n1992;
wire            n1993;
wire      [7:0] n1994;
wire            n1995;
wire      [7:0] n1996;
wire            n1997;
wire      [7:0] n1998;
wire            n1999;
wire      [7:0] n2;
wire      [7:0] n2000;
wire            n2001;
wire      [7:0] n2002;
wire            n2003;
wire      [7:0] n2004;
wire            n2005;
wire      [7:0] n2006;
wire            n2007;
wire      [7:0] n2008;
wire            n2009;
wire            n201;
wire      [7:0] n2010;
wire            n2011;
wire      [7:0] n2012;
wire            n2013;
wire      [7:0] n2014;
wire            n2015;
wire      [7:0] n2016;
wire            n2017;
wire      [7:0] n2018;
wire            n2019;
wire      [7:0] n2020;
wire            n2021;
wire      [7:0] n2022;
wire            n2023;
wire      [7:0] n2024;
wire            n2025;
wire      [7:0] n2026;
wire            n2027;
wire      [7:0] n2028;
wire            n2029;
wire      [7:0] n203;
wire      [7:0] n2030;
wire            n2031;
wire      [7:0] n2032;
wire            n2033;
wire      [7:0] n2034;
wire            n2035;
wire      [7:0] n2036;
wire            n2037;
wire      [7:0] n2038;
wire            n2039;
wire      [7:0] n2040;
wire            n2041;
wire      [7:0] n2042;
wire            n2043;
wire      [7:0] n2044;
wire            n2045;
wire      [7:0] n2046;
wire            n2047;
wire      [7:0] n2048;
wire            n2049;
wire            n205;
wire      [7:0] n2050;
wire            n2051;
wire      [7:0] n2052;
wire            n2053;
wire      [7:0] n2054;
wire            n2055;
wire      [7:0] n2056;
wire            n2057;
wire      [7:0] n2058;
wire            n2059;
wire      [7:0] n2060;
wire            n2061;
wire      [7:0] n2062;
wire            n2063;
wire      [7:0] n2064;
wire            n2065;
wire      [7:0] n2066;
wire            n2067;
wire      [7:0] n2068;
wire            n2069;
wire      [7:0] n207;
wire      [7:0] n2070;
wire            n2071;
wire      [7:0] n2072;
wire            n2073;
wire      [7:0] n2074;
wire            n2075;
wire      [7:0] n2076;
wire            n2077;
wire      [7:0] n2078;
wire            n2079;
wire      [7:0] n2080;
wire            n2081;
wire      [7:0] n2082;
wire            n2083;
wire      [7:0] n2084;
wire            n2085;
wire      [7:0] n2086;
wire            n2087;
wire      [7:0] n2088;
wire            n2089;
wire            n209;
wire      [7:0] n2090;
wire            n2091;
wire      [7:0] n2092;
wire            n2093;
wire      [7:0] n2094;
wire            n2095;
wire      [7:0] n2096;
wire            n2097;
wire      [7:0] n2098;
wire            n2099;
wire            n21;
wire      [7:0] n2100;
wire            n2101;
wire      [7:0] n2102;
wire            n2103;
wire      [7:0] n2104;
wire            n2105;
wire      [7:0] n2106;
wire            n2107;
wire      [7:0] n2108;
wire            n2109;
wire      [7:0] n211;
wire      [7:0] n2110;
wire            n2111;
wire      [7:0] n2112;
wire            n2113;
wire      [7:0] n2114;
wire            n2115;
wire      [7:0] n2116;
wire            n2117;
wire      [7:0] n2118;
wire            n2119;
wire      [7:0] n2120;
wire            n2121;
wire      [7:0] n2122;
wire            n2123;
wire      [7:0] n2124;
wire            n2125;
wire      [7:0] n2126;
wire            n2127;
wire      [7:0] n2128;
wire            n2129;
wire            n213;
wire      [7:0] n2130;
wire            n2131;
wire      [7:0] n2132;
wire            n2133;
wire      [7:0] n2134;
wire            n2135;
wire      [7:0] n2136;
wire            n2137;
wire      [7:0] n2138;
wire            n2139;
wire      [7:0] n214;
wire      [7:0] n2140;
wire            n2141;
wire      [7:0] n2142;
wire            n2143;
wire      [7:0] n2144;
wire            n2145;
wire      [7:0] n2146;
wire            n2147;
wire      [7:0] n2148;
wire            n2149;
wire      [7:0] n2150;
wire            n2151;
wire      [7:0] n2152;
wire            n2153;
wire      [7:0] n2154;
wire            n2155;
wire      [7:0] n2156;
wire            n2157;
wire      [7:0] n2158;
wire            n2159;
wire            n216;
wire      [7:0] n2160;
wire            n2161;
wire      [7:0] n2162;
wire            n2163;
wire      [7:0] n2164;
wire            n2165;
wire      [7:0] n2166;
wire            n2167;
wire      [7:0] n2168;
wire            n2169;
wire      [7:0] n217;
wire      [7:0] n2170;
wire            n2171;
wire      [7:0] n2172;
wire            n2173;
wire      [7:0] n2174;
wire            n2175;
wire      [7:0] n2176;
wire            n2177;
wire      [7:0] n2178;
wire            n2179;
wire      [7:0] n2180;
wire            n2181;
wire      [7:0] n2182;
wire            n2183;
wire      [7:0] n2184;
wire            n2185;
wire      [7:0] n2186;
wire            n2187;
wire      [7:0] n2188;
wire            n2189;
wire            n219;
wire      [7:0] n2190;
wire            n2191;
wire      [7:0] n2192;
wire            n2193;
wire      [7:0] n2194;
wire            n2195;
wire      [7:0] n2196;
wire            n2197;
wire      [7:0] n2198;
wire            n2199;
wire      [7:0] n2200;
wire            n2201;
wire      [7:0] n2202;
wire            n2203;
wire      [7:0] n2204;
wire            n2205;
wire      [7:0] n2206;
wire            n2207;
wire      [7:0] n2208;
wire            n2209;
wire      [7:0] n221;
wire      [7:0] n2210;
wire            n2211;
wire      [7:0] n2212;
wire            n2213;
wire      [7:0] n2214;
wire            n2215;
wire      [7:0] n2216;
wire            n2217;
wire      [7:0] n2218;
wire            n2219;
wire            n222;
wire      [7:0] n2220;
wire            n2221;
wire      [7:0] n2222;
wire            n2223;
wire      [7:0] n2224;
wire            n2225;
wire      [7:0] n2226;
wire            n2227;
wire      [7:0] n2228;
wire            n2229;
wire      [7:0] n2230;
wire            n2231;
wire      [7:0] n2232;
wire            n2233;
wire      [7:0] n2234;
wire            n2235;
wire      [7:0] n2236;
wire            n2237;
wire      [7:0] n2238;
wire            n2239;
wire      [7:0] n224;
wire      [7:0] n2240;
wire            n2241;
wire      [7:0] n2242;
wire            n2243;
wire      [7:0] n2244;
wire            n2245;
wire      [7:0] n2246;
wire            n2247;
wire      [7:0] n2248;
wire            n2249;
wire      [7:0] n2250;
wire            n2251;
wire      [7:0] n2252;
wire            n2253;
wire      [7:0] n2254;
wire            n2255;
wire      [7:0] n2256;
wire            n2257;
wire      [7:0] n2258;
wire            n2259;
wire            n226;
wire      [7:0] n2260;
wire            n2261;
wire      [7:0] n2262;
wire            n2263;
wire      [7:0] n2264;
wire            n2265;
wire      [7:0] n2266;
wire            n2267;
wire      [7:0] n2268;
wire            n2269;
wire      [7:0] n2270;
wire            n2271;
wire      [7:0] n2272;
wire            n2273;
wire      [7:0] n2274;
wire            n2275;
wire      [7:0] n2276;
wire            n2277;
wire      [7:0] n2278;
wire            n2279;
wire      [7:0] n228;
wire      [7:0] n2280;
wire            n2281;
wire      [7:0] n2282;
wire            n2283;
wire      [7:0] n2284;
wire            n2285;
wire      [7:0] n2286;
wire            n2287;
wire      [7:0] n2288;
wire            n2289;
wire      [7:0] n2290;
wire            n2291;
wire      [7:0] n2292;
wire            n2293;
wire      [7:0] n2294;
wire            n2295;
wire      [7:0] n2296;
wire            n2297;
wire      [7:0] n2298;
wire            n2299;
wire      [7:0] n23;
wire            n230;
wire      [7:0] n2300;
wire            n2301;
wire      [7:0] n2302;
wire            n2303;
wire      [7:0] n2304;
wire            n2305;
wire      [7:0] n2306;
wire            n2307;
wire      [7:0] n2308;
wire            n2309;
wire      [7:0] n2310;
wire            n2311;
wire      [7:0] n2312;
wire      [7:0] n2313;
wire      [7:0] n2314;
wire      [7:0] n2315;
wire      [7:0] n2316;
wire      [7:0] n2317;
wire      [7:0] n2318;
wire      [7:0] n2319;
wire      [7:0] n232;
wire      [7:0] n2320;
wire      [7:0] n2321;
wire      [7:0] n2322;
wire      [7:0] n2323;
wire      [7:0] n2324;
wire      [7:0] n2325;
wire      [7:0] n2326;
wire      [7:0] n2327;
wire      [7:0] n2328;
wire      [7:0] n2329;
wire      [7:0] n2330;
wire      [7:0] n2331;
wire      [7:0] n2332;
wire      [7:0] n2333;
wire      [7:0] n2334;
wire      [7:0] n2335;
wire      [7:0] n2336;
wire      [7:0] n2337;
wire      [7:0] n2338;
wire      [7:0] n2339;
wire            n234;
wire      [7:0] n2340;
wire      [7:0] n2341;
wire      [7:0] n2342;
wire      [7:0] n2343;
wire      [7:0] n2344;
wire      [7:0] n2345;
wire      [7:0] n2346;
wire      [7:0] n2347;
wire      [7:0] n2348;
wire      [7:0] n2349;
wire      [7:0] n2350;
wire      [7:0] n2351;
wire      [7:0] n2352;
wire      [7:0] n2353;
wire      [7:0] n2354;
wire      [7:0] n2355;
wire      [7:0] n2356;
wire      [7:0] n2357;
wire      [7:0] n2358;
wire      [7:0] n2359;
wire      [7:0] n236;
wire      [7:0] n2360;
wire      [7:0] n2361;
wire      [7:0] n2362;
wire      [7:0] n2363;
wire      [7:0] n2364;
wire      [7:0] n2365;
wire      [7:0] n2366;
wire      [7:0] n2367;
wire      [7:0] n2368;
wire      [7:0] n2369;
wire      [7:0] n2370;
wire      [7:0] n2371;
wire      [7:0] n2372;
wire      [7:0] n2373;
wire      [7:0] n2374;
wire      [7:0] n2375;
wire      [7:0] n2376;
wire      [7:0] n2377;
wire      [7:0] n2378;
wire      [7:0] n2379;
wire            n238;
wire      [7:0] n2380;
wire      [7:0] n2381;
wire      [7:0] n2382;
wire      [7:0] n2383;
wire      [7:0] n2384;
wire      [7:0] n2385;
wire      [7:0] n2386;
wire      [7:0] n2387;
wire      [7:0] n2388;
wire      [7:0] n2389;
wire      [7:0] n2390;
wire      [7:0] n2391;
wire      [7:0] n2392;
wire      [7:0] n2393;
wire      [7:0] n2394;
wire      [7:0] n2395;
wire      [7:0] n2396;
wire      [7:0] n2397;
wire      [7:0] n2398;
wire      [7:0] n2399;
wire      [7:0] n240;
wire      [7:0] n2400;
wire      [7:0] n2401;
wire      [7:0] n2402;
wire      [7:0] n2403;
wire      [7:0] n2404;
wire      [7:0] n2405;
wire      [7:0] n2406;
wire      [7:0] n2407;
wire      [7:0] n2408;
wire      [7:0] n2409;
wire            n241;
wire      [7:0] n2410;
wire      [7:0] n2411;
wire      [7:0] n2412;
wire      [7:0] n2413;
wire      [7:0] n2414;
wire      [7:0] n2415;
wire      [7:0] n2416;
wire      [7:0] n2417;
wire      [7:0] n2418;
wire      [7:0] n2419;
wire      [7:0] n2420;
wire      [7:0] n2421;
wire      [7:0] n2422;
wire      [7:0] n2423;
wire      [7:0] n2424;
wire      [7:0] n2425;
wire      [7:0] n2426;
wire      [7:0] n2427;
wire      [7:0] n2428;
wire      [7:0] n2429;
wire      [7:0] n243;
wire      [7:0] n2430;
wire      [7:0] n2431;
wire      [7:0] n2432;
wire      [7:0] n2433;
wire      [7:0] n2434;
wire      [7:0] n2435;
wire      [7:0] n2436;
wire      [7:0] n2437;
wire      [7:0] n2438;
wire      [7:0] n2439;
wire      [7:0] n2440;
wire      [7:0] n2441;
wire      [7:0] n2442;
wire      [7:0] n2443;
wire      [7:0] n2444;
wire      [7:0] n2445;
wire      [7:0] n2446;
wire      [7:0] n2447;
wire      [7:0] n2448;
wire      [7:0] n2449;
wire            n245;
wire      [7:0] n2450;
wire      [7:0] n2451;
wire      [7:0] n2452;
wire      [7:0] n2453;
wire      [7:0] n2454;
wire      [7:0] n2455;
wire      [7:0] n2456;
wire      [7:0] n2457;
wire      [7:0] n2458;
wire      [7:0] n2459;
wire      [7:0] n2460;
wire      [7:0] n2461;
wire      [7:0] n2462;
wire      [7:0] n2463;
wire      [7:0] n2464;
wire      [7:0] n2465;
wire      [7:0] n2466;
wire      [7:0] n2467;
wire      [7:0] n2468;
wire      [7:0] n2469;
wire      [7:0] n247;
wire      [7:0] n2470;
wire      [7:0] n2471;
wire      [7:0] n2472;
wire      [7:0] n2473;
wire      [7:0] n2474;
wire      [7:0] n2475;
wire      [7:0] n2476;
wire      [7:0] n2477;
wire      [7:0] n2478;
wire      [7:0] n2479;
wire            n248;
wire      [7:0] n2480;
wire      [7:0] n2481;
wire      [7:0] n2482;
wire      [7:0] n2483;
wire      [7:0] n2484;
wire      [7:0] n2485;
wire      [7:0] n2486;
wire      [7:0] n2487;
wire      [7:0] n2488;
wire      [7:0] n2489;
wire      [7:0] n2490;
wire      [7:0] n2491;
wire      [7:0] n2492;
wire      [7:0] n2493;
wire      [7:0] n2494;
wire      [7:0] n2495;
wire      [7:0] n2496;
wire      [7:0] n2497;
wire      [7:0] n2498;
wire      [7:0] n2499;
wire            n25;
wire      [7:0] n250;
wire      [7:0] n2500;
wire      [7:0] n2501;
wire      [7:0] n2502;
wire      [7:0] n2503;
wire      [7:0] n2504;
wire      [7:0] n2505;
wire      [7:0] n2506;
wire      [7:0] n2507;
wire      [7:0] n2508;
wire      [7:0] n2509;
wire      [7:0] n2510;
wire      [7:0] n2511;
wire      [7:0] n2512;
wire      [7:0] n2513;
wire      [7:0] n2514;
wire      [7:0] n2515;
wire      [7:0] n2516;
wire      [7:0] n2517;
wire      [7:0] n2518;
wire      [7:0] n2519;
wire            n252;
wire      [7:0] n2520;
wire      [7:0] n2521;
wire      [7:0] n2522;
wire      [7:0] n2523;
wire      [7:0] n2524;
wire      [7:0] n2525;
wire      [7:0] n2526;
wire      [7:0] n2527;
wire      [7:0] n2528;
wire      [7:0] n2529;
wire      [7:0] n2530;
wire      [7:0] n2531;
wire      [7:0] n2532;
wire      [7:0] n2533;
wire      [7:0] n2534;
wire      [7:0] n2535;
wire      [7:0] n2536;
wire      [7:0] n2537;
wire      [7:0] n2538;
wire      [7:0] n2539;
wire      [7:0] n254;
wire      [7:0] n2540;
wire      [7:0] n2541;
wire      [7:0] n2542;
wire      [7:0] n2543;
wire      [7:0] n2544;
wire      [7:0] n2545;
wire      [7:0] n2546;
wire      [7:0] n2547;
wire      [7:0] n2548;
wire      [7:0] n2549;
wire            n255;
wire      [7:0] n2550;
wire      [7:0] n2551;
wire      [7:0] n2552;
wire      [7:0] n2553;
wire      [7:0] n2554;
wire      [7:0] n2555;
wire      [7:0] n2556;
wire      [7:0] n2557;
wire      [7:0] n2558;
wire      [7:0] n2559;
wire      [7:0] n2560;
wire      [7:0] n2561;
wire      [7:0] n2562;
wire      [7:0] n2563;
wire      [7:0] n2564;
wire      [7:0] n2565;
wire      [7:0] n2566;
wire      [7:0] n2567;
wire      [7:0] n2568;
wire     [23:0] n2569;
wire      [7:0] n257;
wire      [7:0] n2570;
wire      [7:0] n2571;
wire            n2572;
wire      [7:0] n2573;
wire            n2574;
wire      [7:0] n2575;
wire            n2576;
wire      [7:0] n2577;
wire            n2578;
wire      [7:0] n2579;
wire            n2580;
wire      [7:0] n2581;
wire            n2582;
wire      [7:0] n2583;
wire            n2584;
wire      [7:0] n2585;
wire            n2586;
wire      [7:0] n2587;
wire            n2588;
wire      [7:0] n2589;
wire            n259;
wire            n2590;
wire      [7:0] n2591;
wire            n2592;
wire      [7:0] n2593;
wire            n2594;
wire      [7:0] n2595;
wire            n2596;
wire      [7:0] n2597;
wire            n2598;
wire      [7:0] n2599;
wire            n2600;
wire      [7:0] n2601;
wire            n2602;
wire      [7:0] n2603;
wire            n2604;
wire      [7:0] n2605;
wire            n2606;
wire      [7:0] n2607;
wire            n2608;
wire      [7:0] n2609;
wire      [7:0] n261;
wire            n2610;
wire      [7:0] n2611;
wire            n2612;
wire      [7:0] n2613;
wire            n2614;
wire      [7:0] n2615;
wire            n2616;
wire      [7:0] n2617;
wire            n2618;
wire      [7:0] n2619;
wire            n262;
wire            n2620;
wire      [7:0] n2621;
wire            n2622;
wire      [7:0] n2623;
wire            n2624;
wire      [7:0] n2625;
wire            n2626;
wire      [7:0] n2627;
wire            n2628;
wire      [7:0] n2629;
wire      [7:0] n263;
wire            n2630;
wire      [7:0] n2631;
wire            n2632;
wire      [7:0] n2633;
wire            n2634;
wire      [7:0] n2635;
wire            n2636;
wire      [7:0] n2637;
wire            n2638;
wire      [7:0] n2639;
wire            n264;
wire            n2640;
wire      [7:0] n2641;
wire            n2642;
wire      [7:0] n2643;
wire            n2644;
wire      [7:0] n2645;
wire            n2646;
wire      [7:0] n2647;
wire            n2648;
wire      [7:0] n2649;
wire      [7:0] n265;
wire            n2650;
wire      [7:0] n2651;
wire            n2652;
wire      [7:0] n2653;
wire            n2654;
wire      [7:0] n2655;
wire            n2656;
wire      [7:0] n2657;
wire            n2658;
wire      [7:0] n2659;
wire            n266;
wire            n2660;
wire      [7:0] n2661;
wire            n2662;
wire      [7:0] n2663;
wire            n2664;
wire      [7:0] n2665;
wire            n2666;
wire      [7:0] n2667;
wire            n2668;
wire      [7:0] n2669;
wire            n2670;
wire      [7:0] n2671;
wire            n2672;
wire      [7:0] n2673;
wire            n2674;
wire      [7:0] n2675;
wire            n2676;
wire      [7:0] n2677;
wire            n2678;
wire      [7:0] n2679;
wire      [7:0] n268;
wire            n2680;
wire      [7:0] n2681;
wire            n2682;
wire      [7:0] n2683;
wire            n2684;
wire      [7:0] n2685;
wire            n2686;
wire      [7:0] n2687;
wire            n2688;
wire      [7:0] n2689;
wire            n2690;
wire      [7:0] n2691;
wire            n2692;
wire      [7:0] n2693;
wire            n2694;
wire      [7:0] n2695;
wire            n2696;
wire      [7:0] n2697;
wire            n2698;
wire      [7:0] n2699;
wire      [7:0] n27;
wire            n270;
wire            n2700;
wire      [7:0] n2701;
wire            n2702;
wire      [7:0] n2703;
wire            n2704;
wire      [7:0] n2705;
wire            n2706;
wire      [7:0] n2707;
wire            n2708;
wire      [7:0] n2709;
wire            n2710;
wire      [7:0] n2711;
wire            n2712;
wire      [7:0] n2713;
wire            n2714;
wire      [7:0] n2715;
wire            n2716;
wire      [7:0] n2717;
wire            n2718;
wire      [7:0] n2719;
wire      [7:0] n272;
wire            n2720;
wire      [7:0] n2721;
wire            n2722;
wire      [7:0] n2723;
wire            n2724;
wire      [7:0] n2725;
wire            n2726;
wire      [7:0] n2727;
wire            n2728;
wire      [7:0] n2729;
wire            n2730;
wire      [7:0] n2731;
wire            n2732;
wire      [7:0] n2733;
wire            n2734;
wire      [7:0] n2735;
wire            n2736;
wire      [7:0] n2737;
wire            n2738;
wire      [7:0] n2739;
wire            n274;
wire            n2740;
wire      [7:0] n2741;
wire            n2742;
wire      [7:0] n2743;
wire            n2744;
wire      [7:0] n2745;
wire            n2746;
wire      [7:0] n2747;
wire            n2748;
wire      [7:0] n2749;
wire            n2750;
wire      [7:0] n2751;
wire            n2752;
wire      [7:0] n2753;
wire            n2754;
wire      [7:0] n2755;
wire            n2756;
wire      [7:0] n2757;
wire            n2758;
wire      [7:0] n2759;
wire      [7:0] n276;
wire            n2760;
wire      [7:0] n2761;
wire            n2762;
wire      [7:0] n2763;
wire            n2764;
wire      [7:0] n2765;
wire            n2766;
wire      [7:0] n2767;
wire            n2768;
wire      [7:0] n2769;
wire            n2770;
wire      [7:0] n2771;
wire            n2772;
wire      [7:0] n2773;
wire            n2774;
wire      [7:0] n2775;
wire            n2776;
wire      [7:0] n2777;
wire            n2778;
wire      [7:0] n2779;
wire            n278;
wire            n2780;
wire      [7:0] n2781;
wire            n2782;
wire      [7:0] n2783;
wire            n2784;
wire      [7:0] n2785;
wire            n2786;
wire      [7:0] n2787;
wire            n2788;
wire      [7:0] n2789;
wire            n2790;
wire      [7:0] n2791;
wire            n2792;
wire      [7:0] n2793;
wire            n2794;
wire      [7:0] n2795;
wire            n2796;
wire      [7:0] n2797;
wire            n2798;
wire      [7:0] n2799;
wire      [7:0] n280;
wire            n2800;
wire      [7:0] n2801;
wire            n2802;
wire      [7:0] n2803;
wire            n2804;
wire      [7:0] n2805;
wire            n2806;
wire      [7:0] n2807;
wire            n2808;
wire      [7:0] n2809;
wire            n281;
wire            n2810;
wire      [7:0] n2811;
wire            n2812;
wire      [7:0] n2813;
wire            n2814;
wire      [7:0] n2815;
wire            n2816;
wire      [7:0] n2817;
wire            n2818;
wire      [7:0] n2819;
wire      [7:0] n282;
wire            n2820;
wire      [7:0] n2821;
wire            n2822;
wire      [7:0] n2823;
wire            n2824;
wire      [7:0] n2825;
wire            n2826;
wire      [7:0] n2827;
wire            n2828;
wire      [7:0] n2829;
wire            n283;
wire            n2830;
wire      [7:0] n2831;
wire            n2832;
wire      [7:0] n2833;
wire            n2834;
wire      [7:0] n2835;
wire            n2836;
wire      [7:0] n2837;
wire            n2838;
wire      [7:0] n2839;
wire            n2840;
wire      [7:0] n2841;
wire            n2842;
wire      [7:0] n2843;
wire            n2844;
wire      [7:0] n2845;
wire            n2846;
wire      [7:0] n2847;
wire            n2848;
wire      [7:0] n2849;
wire      [7:0] n285;
wire            n2850;
wire      [7:0] n2851;
wire            n2852;
wire      [7:0] n2853;
wire            n2854;
wire      [7:0] n2855;
wire            n2856;
wire      [7:0] n2857;
wire            n2858;
wire      [7:0] n2859;
wire            n2860;
wire      [7:0] n2861;
wire            n2862;
wire      [7:0] n2863;
wire            n2864;
wire      [7:0] n2865;
wire            n2866;
wire      [7:0] n2867;
wire            n2868;
wire      [7:0] n2869;
wire            n287;
wire            n2870;
wire      [7:0] n2871;
wire            n2872;
wire      [7:0] n2873;
wire            n2874;
wire      [7:0] n2875;
wire            n2876;
wire      [7:0] n2877;
wire            n2878;
wire      [7:0] n2879;
wire            n2880;
wire      [7:0] n2881;
wire            n2882;
wire      [7:0] n2883;
wire            n2884;
wire      [7:0] n2885;
wire            n2886;
wire      [7:0] n2887;
wire            n2888;
wire      [7:0] n2889;
wire      [7:0] n289;
wire            n2890;
wire      [7:0] n2891;
wire            n2892;
wire      [7:0] n2893;
wire            n2894;
wire      [7:0] n2895;
wire            n2896;
wire      [7:0] n2897;
wire            n2898;
wire      [7:0] n2899;
wire            n29;
wire            n2900;
wire      [7:0] n2901;
wire            n2902;
wire      [7:0] n2903;
wire            n2904;
wire      [7:0] n2905;
wire            n2906;
wire      [7:0] n2907;
wire            n2908;
wire      [7:0] n2909;
wire            n291;
wire            n2910;
wire      [7:0] n2911;
wire            n2912;
wire      [7:0] n2913;
wire            n2914;
wire      [7:0] n2915;
wire            n2916;
wire      [7:0] n2917;
wire            n2918;
wire      [7:0] n2919;
wire            n2920;
wire      [7:0] n2921;
wire            n2922;
wire      [7:0] n2923;
wire            n2924;
wire      [7:0] n2925;
wire            n2926;
wire      [7:0] n2927;
wire            n2928;
wire      [7:0] n2929;
wire      [7:0] n293;
wire            n2930;
wire      [7:0] n2931;
wire            n2932;
wire      [7:0] n2933;
wire            n2934;
wire      [7:0] n2935;
wire            n2936;
wire      [7:0] n2937;
wire            n2938;
wire      [7:0] n2939;
wire            n2940;
wire      [7:0] n2941;
wire            n2942;
wire      [7:0] n2943;
wire            n2944;
wire      [7:0] n2945;
wire            n2946;
wire      [7:0] n2947;
wire            n2948;
wire      [7:0] n2949;
wire            n295;
wire            n2950;
wire      [7:0] n2951;
wire            n2952;
wire      [7:0] n2953;
wire            n2954;
wire      [7:0] n2955;
wire            n2956;
wire      [7:0] n2957;
wire            n2958;
wire      [7:0] n2959;
wire      [7:0] n296;
wire            n2960;
wire      [7:0] n2961;
wire            n2962;
wire      [7:0] n2963;
wire            n2964;
wire      [7:0] n2965;
wire            n2966;
wire      [7:0] n2967;
wire            n2968;
wire      [7:0] n2969;
wire            n297;
wire            n2970;
wire      [7:0] n2971;
wire            n2972;
wire      [7:0] n2973;
wire            n2974;
wire      [7:0] n2975;
wire            n2976;
wire      [7:0] n2977;
wire            n2978;
wire      [7:0] n2979;
wire      [7:0] n298;
wire            n2980;
wire      [7:0] n2981;
wire            n2982;
wire      [7:0] n2983;
wire            n2984;
wire      [7:0] n2985;
wire            n2986;
wire      [7:0] n2987;
wire            n2988;
wire      [7:0] n2989;
wire            n2990;
wire      [7:0] n2991;
wire            n2992;
wire      [7:0] n2993;
wire            n2994;
wire      [7:0] n2995;
wire            n2996;
wire      [7:0] n2997;
wire            n2998;
wire      [7:0] n2999;
wire      [7:0] n3;
wire            n300;
wire            n3000;
wire      [7:0] n3001;
wire            n3002;
wire      [7:0] n3003;
wire            n3004;
wire      [7:0] n3005;
wire            n3006;
wire      [7:0] n3007;
wire            n3008;
wire      [7:0] n3009;
wire            n3010;
wire      [7:0] n3011;
wire            n3012;
wire      [7:0] n3013;
wire            n3014;
wire      [7:0] n3015;
wire            n3016;
wire      [7:0] n3017;
wire            n3018;
wire      [7:0] n3019;
wire      [7:0] n302;
wire            n3020;
wire      [7:0] n3021;
wire            n3022;
wire      [7:0] n3023;
wire            n3024;
wire      [7:0] n3025;
wire            n3026;
wire      [7:0] n3027;
wire            n3028;
wire      [7:0] n3029;
wire            n303;
wire            n3030;
wire      [7:0] n3031;
wire            n3032;
wire      [7:0] n3033;
wire            n3034;
wire      [7:0] n3035;
wire            n3036;
wire      [7:0] n3037;
wire            n3038;
wire      [7:0] n3039;
wire      [7:0] n304;
wire            n3040;
wire      [7:0] n3041;
wire            n3042;
wire      [7:0] n3043;
wire            n3044;
wire      [7:0] n3045;
wire            n3046;
wire      [7:0] n3047;
wire            n3048;
wire      [7:0] n3049;
wire            n3050;
wire      [7:0] n3051;
wire            n3052;
wire      [7:0] n3053;
wire            n3054;
wire      [7:0] n3055;
wire            n3056;
wire      [7:0] n3057;
wire            n3058;
wire      [7:0] n3059;
wire            n306;
wire            n3060;
wire      [7:0] n3061;
wire            n3062;
wire      [7:0] n3063;
wire            n3064;
wire      [7:0] n3065;
wire            n3066;
wire      [7:0] n3067;
wire            n3068;
wire      [7:0] n3069;
wire            n3070;
wire      [7:0] n3071;
wire            n3072;
wire      [7:0] n3073;
wire            n3074;
wire      [7:0] n3075;
wire            n3076;
wire      [7:0] n3077;
wire            n3078;
wire      [7:0] n3079;
wire      [7:0] n308;
wire            n3080;
wire      [7:0] n3081;
wire            n3082;
wire      [7:0] n3083;
wire      [7:0] n3084;
wire      [7:0] n3085;
wire      [7:0] n3086;
wire      [7:0] n3087;
wire      [7:0] n3088;
wire      [7:0] n3089;
wire      [7:0] n3090;
wire      [7:0] n3091;
wire      [7:0] n3092;
wire      [7:0] n3093;
wire      [7:0] n3094;
wire      [7:0] n3095;
wire      [7:0] n3096;
wire      [7:0] n3097;
wire      [7:0] n3098;
wire      [7:0] n3099;
wire      [7:0] n31;
wire            n310;
wire      [7:0] n3100;
wire      [7:0] n3101;
wire      [7:0] n3102;
wire      [7:0] n3103;
wire      [7:0] n3104;
wire      [7:0] n3105;
wire      [7:0] n3106;
wire      [7:0] n3107;
wire      [7:0] n3108;
wire      [7:0] n3109;
wire      [7:0] n3110;
wire      [7:0] n3111;
wire      [7:0] n3112;
wire      [7:0] n3113;
wire      [7:0] n3114;
wire      [7:0] n3115;
wire      [7:0] n3116;
wire      [7:0] n3117;
wire      [7:0] n3118;
wire      [7:0] n3119;
wire      [7:0] n312;
wire      [7:0] n3120;
wire      [7:0] n3121;
wire      [7:0] n3122;
wire      [7:0] n3123;
wire      [7:0] n3124;
wire      [7:0] n3125;
wire      [7:0] n3126;
wire      [7:0] n3127;
wire      [7:0] n3128;
wire      [7:0] n3129;
wire      [7:0] n3130;
wire      [7:0] n3131;
wire      [7:0] n3132;
wire      [7:0] n3133;
wire      [7:0] n3134;
wire      [7:0] n3135;
wire      [7:0] n3136;
wire      [7:0] n3137;
wire      [7:0] n3138;
wire      [7:0] n3139;
wire            n314;
wire      [7:0] n3140;
wire      [7:0] n3141;
wire      [7:0] n3142;
wire      [7:0] n3143;
wire      [7:0] n3144;
wire      [7:0] n3145;
wire      [7:0] n3146;
wire      [7:0] n3147;
wire      [7:0] n3148;
wire      [7:0] n3149;
wire      [7:0] n3150;
wire      [7:0] n3151;
wire      [7:0] n3152;
wire      [7:0] n3153;
wire      [7:0] n3154;
wire      [7:0] n3155;
wire      [7:0] n3156;
wire      [7:0] n3157;
wire      [7:0] n3158;
wire      [7:0] n3159;
wire      [7:0] n316;
wire      [7:0] n3160;
wire      [7:0] n3161;
wire      [7:0] n3162;
wire      [7:0] n3163;
wire      [7:0] n3164;
wire      [7:0] n3165;
wire      [7:0] n3166;
wire      [7:0] n3167;
wire      [7:0] n3168;
wire      [7:0] n3169;
wire      [7:0] n3170;
wire      [7:0] n3171;
wire      [7:0] n3172;
wire      [7:0] n3173;
wire      [7:0] n3174;
wire      [7:0] n3175;
wire      [7:0] n3176;
wire      [7:0] n3177;
wire      [7:0] n3178;
wire      [7:0] n3179;
wire            n318;
wire      [7:0] n3180;
wire      [7:0] n3181;
wire      [7:0] n3182;
wire      [7:0] n3183;
wire      [7:0] n3184;
wire      [7:0] n3185;
wire      [7:0] n3186;
wire      [7:0] n3187;
wire      [7:0] n3188;
wire      [7:0] n3189;
wire      [7:0] n319;
wire      [7:0] n3190;
wire      [7:0] n3191;
wire      [7:0] n3192;
wire      [7:0] n3193;
wire      [7:0] n3194;
wire      [7:0] n3195;
wire      [7:0] n3196;
wire      [7:0] n3197;
wire      [7:0] n3198;
wire      [7:0] n3199;
wire            n320;
wire      [7:0] n3200;
wire      [7:0] n3201;
wire      [7:0] n3202;
wire      [7:0] n3203;
wire      [7:0] n3204;
wire      [7:0] n3205;
wire      [7:0] n3206;
wire      [7:0] n3207;
wire      [7:0] n3208;
wire      [7:0] n3209;
wire      [7:0] n321;
wire      [7:0] n3210;
wire      [7:0] n3211;
wire      [7:0] n3212;
wire      [7:0] n3213;
wire      [7:0] n3214;
wire      [7:0] n3215;
wire      [7:0] n3216;
wire      [7:0] n3217;
wire      [7:0] n3218;
wire      [7:0] n3219;
wire      [7:0] n3220;
wire      [7:0] n3221;
wire      [7:0] n3222;
wire      [7:0] n3223;
wire      [7:0] n3224;
wire      [7:0] n3225;
wire      [7:0] n3226;
wire      [7:0] n3227;
wire      [7:0] n3228;
wire      [7:0] n3229;
wire            n323;
wire      [7:0] n3230;
wire      [7:0] n3231;
wire      [7:0] n3232;
wire      [7:0] n3233;
wire      [7:0] n3234;
wire      [7:0] n3235;
wire      [7:0] n3236;
wire      [7:0] n3237;
wire      [7:0] n3238;
wire      [7:0] n3239;
wire      [7:0] n324;
wire      [7:0] n3240;
wire      [7:0] n3241;
wire      [7:0] n3242;
wire      [7:0] n3243;
wire      [7:0] n3244;
wire      [7:0] n3245;
wire      [7:0] n3246;
wire      [7:0] n3247;
wire      [7:0] n3248;
wire      [7:0] n3249;
wire      [7:0] n3250;
wire      [7:0] n3251;
wire      [7:0] n3252;
wire      [7:0] n3253;
wire      [7:0] n3254;
wire      [7:0] n3255;
wire      [7:0] n3256;
wire      [7:0] n3257;
wire      [7:0] n3258;
wire      [7:0] n3259;
wire            n326;
wire      [7:0] n3260;
wire      [7:0] n3261;
wire      [7:0] n3262;
wire      [7:0] n3263;
wire      [7:0] n3264;
wire      [7:0] n3265;
wire      [7:0] n3266;
wire      [7:0] n3267;
wire      [7:0] n3268;
wire      [7:0] n3269;
wire      [7:0] n3270;
wire      [7:0] n3271;
wire      [7:0] n3272;
wire      [7:0] n3273;
wire      [7:0] n3274;
wire      [7:0] n3275;
wire      [7:0] n3276;
wire      [7:0] n3277;
wire      [7:0] n3278;
wire      [7:0] n3279;
wire      [7:0] n328;
wire      [7:0] n3280;
wire      [7:0] n3281;
wire      [7:0] n3282;
wire      [7:0] n3283;
wire      [7:0] n3284;
wire      [7:0] n3285;
wire      [7:0] n3286;
wire      [7:0] n3287;
wire      [7:0] n3288;
wire      [7:0] n3289;
wire            n329;
wire      [7:0] n3290;
wire      [7:0] n3291;
wire      [7:0] n3292;
wire      [7:0] n3293;
wire      [7:0] n3294;
wire      [7:0] n3295;
wire      [7:0] n3296;
wire      [7:0] n3297;
wire      [7:0] n3298;
wire      [7:0] n3299;
wire            n33;
wire      [7:0] n3300;
wire      [7:0] n3301;
wire      [7:0] n3302;
wire      [7:0] n3303;
wire      [7:0] n3304;
wire      [7:0] n3305;
wire      [7:0] n3306;
wire      [7:0] n3307;
wire      [7:0] n3308;
wire      [7:0] n3309;
wire      [7:0] n331;
wire      [7:0] n3310;
wire      [7:0] n3311;
wire      [7:0] n3312;
wire      [7:0] n3313;
wire      [7:0] n3314;
wire      [7:0] n3315;
wire      [7:0] n3316;
wire      [7:0] n3317;
wire      [7:0] n3318;
wire      [7:0] n3319;
wire      [7:0] n3320;
wire      [7:0] n3321;
wire      [7:0] n3322;
wire      [7:0] n3323;
wire      [7:0] n3324;
wire      [7:0] n3325;
wire      [7:0] n3326;
wire      [7:0] n3327;
wire      [7:0] n3328;
wire      [7:0] n3329;
wire            n333;
wire      [7:0] n3330;
wire      [7:0] n3331;
wire      [7:0] n3332;
wire      [7:0] n3333;
wire      [7:0] n3334;
wire      [7:0] n3335;
wire      [7:0] n3336;
wire      [7:0] n3337;
wire      [7:0] n3338;
wire      [7:0] n3339;
wire     [31:0] n3340;
wire      [7:0] n3341;
wire      [7:0] n3342;
wire      [7:0] n3343;
wire      [7:0] n3344;
wire      [7:0] n3345;
wire     [39:0] n3346;
wire      [7:0] n3347;
wire      [7:0] n3348;
wire      [7:0] n3349;
wire      [7:0] n335;
wire      [7:0] n3350;
wire     [47:0] n3351;
wire      [7:0] n3352;
wire      [7:0] n3353;
wire      [7:0] n3354;
wire      [7:0] n3355;
wire     [55:0] n3356;
wire      [7:0] n3357;
wire      [7:0] n3358;
wire      [7:0] n3359;
wire      [7:0] n3360;
wire     [63:0] n3361;
wire      [7:0] n3362;
wire      [7:0] n3363;
wire      [7:0] n3364;
wire      [7:0] n3365;
wire      [7:0] n3366;
wire      [7:0] n3367;
wire      [7:0] n3368;
wire     [71:0] n3369;
wire            n337;
wire      [7:0] n3370;
wire      [7:0] n3371;
wire      [7:0] n3372;
wire      [7:0] n3373;
wire      [7:0] n3374;
wire      [7:0] n3375;
wire     [79:0] n3376;
wire      [7:0] n3377;
wire      [7:0] n3378;
wire      [7:0] n3379;
wire      [7:0] n3380;
wire      [7:0] n3381;
wire      [7:0] n3382;
wire     [87:0] n3383;
wire      [7:0] n3384;
wire      [7:0] n3385;
wire      [7:0] n3386;
wire      [7:0] n3387;
wire      [7:0] n3388;
wire      [7:0] n3389;
wire      [7:0] n339;
wire     [95:0] n3390;
wire      [7:0] n3391;
wire      [7:0] n3392;
wire      [7:0] n3393;
wire      [7:0] n3394;
wire      [7:0] n3395;
wire      [7:0] n3396;
wire      [7:0] n3397;
wire      [7:0] n3398;
wire      [7:0] n3399;
wire    [103:0] n3400;
wire      [7:0] n3401;
wire      [7:0] n3402;
wire      [7:0] n3403;
wire      [7:0] n3404;
wire      [7:0] n3405;
wire      [7:0] n3406;
wire      [7:0] n3407;
wire      [7:0] n3408;
wire    [111:0] n3409;
wire            n341;
wire      [7:0] n3410;
wire      [7:0] n3411;
wire      [7:0] n3412;
wire      [7:0] n3413;
wire      [7:0] n3414;
wire      [7:0] n3415;
wire      [7:0] n3416;
wire      [7:0] n3417;
wire    [119:0] n3418;
wire      [7:0] n3419;
wire      [7:0] n3420;
wire      [7:0] n3421;
wire      [7:0] n3422;
wire      [7:0] n3423;
wire      [7:0] n3424;
wire      [7:0] n3425;
wire      [7:0] n3426;
wire    [127:0] n3427;
wire      [7:0] n343;
wire            n345;
wire      [7:0] n347;
wire            n348;
wire      [7:0] n35;
wire      [7:0] n350;
wire            n352;
wire      [7:0] n353;
wire            n355;
wire      [7:0] n356;
wire            n357;
wire      [7:0] n359;
wire            n361;
wire      [7:0] n363;
wire            n365;
wire      [7:0] n366;
wire            n367;
wire      [7:0] n369;
wire            n37;
wire            n371;
wire      [7:0] n372;
wire            n373;
wire      [7:0] n374;
wire            n375;
wire      [7:0] n377;
wire            n379;
wire      [7:0] n381;
wire            n383;
wire      [7:0] n385;
wire            n386;
wire      [7:0] n388;
wire            n389;
wire      [7:0] n39;
wire      [7:0] n391;
wire            n393;
wire      [7:0] n394;
wire            n396;
wire      [7:0] n398;
wire            n399;
wire      [7:0] n401;
wire            n402;
wire      [7:0] n404;
wire            n406;
wire      [7:0] n408;
wire            n409;
wire            n41;
wire      [7:0] n411;
wire            n412;
wire      [7:0] n414;
wire            n415;
wire      [7:0] n417;
wire            n418;
wire      [7:0] n420;
wire            n421;
wire      [7:0] n423;
wire            n424;
wire      [7:0] n425;
wire            n426;
wire      [7:0] n427;
wire            n428;
wire      [7:0] n43;
wire      [7:0] n430;
wire            n431;
wire      [7:0] n433;
wire            n435;
wire      [7:0] n436;
wire            n438;
wire      [7:0] n440;
wire            n442;
wire      [7:0] n443;
wire            n445;
wire      [7:0] n447;
wire            n448;
wire            n45;
wire      [7:0] n450;
wire            n452;
wire      [7:0] n453;
wire            n455;
wire      [7:0] n456;
wire            n457;
wire      [7:0] n458;
wire            n460;
wire      [7:0] n461;
wire            n463;
wire      [7:0] n465;
wire            n467;
wire      [7:0] n469;
wire      [7:0] n47;
wire            n470;
wire      [7:0] n471;
wire            n472;
wire      [7:0] n473;
wire            n474;
wire      [7:0] n475;
wire            n477;
wire      [7:0] n478;
wire            n480;
wire      [7:0] n482;
wire            n484;
wire      [7:0] n485;
wire            n486;
wire      [7:0] n487;
wire            n488;
wire      [7:0] n489;
wire            n49;
wire            n491;
wire      [7:0] n493;
wire            n495;
wire      [7:0] n496;
wire            n497;
wire      [7:0] n499;
wire            n5;
wire            n501;
wire      [7:0] n502;
wire            n504;
wire      [7:0] n505;
wire            n506;
wire      [7:0] n508;
wire            n509;
wire      [7:0] n51;
wire      [7:0] n511;
wire            n513;
wire      [7:0] n514;
wire            n516;
wire      [7:0] n518;
wire            n519;
wire      [7:0] n520;
wire            n521;
wire      [7:0] n523;
wire            n525;
wire      [7:0] n526;
wire            n527;
wire      [7:0] n529;
wire            n53;
wire            n530;
wire      [7:0] n532;
wire            n533;
wire      [7:0] n535;
wire            n537;
wire      [7:0] n538;
wire            n539;
wire      [7:0] n540;
wire            n541;
wire      [7:0] n542;
wire            n543;
wire      [7:0] n544;
wire            n545;
wire      [7:0] n546;
wire            n547;
wire      [7:0] n549;
wire      [7:0] n55;
wire            n550;
wire      [7:0] n552;
wire            n553;
wire      [7:0] n555;
wire            n557;
wire      [7:0] n559;
wire            n561;
wire      [7:0] n562;
wire            n564;
wire      [7:0] n565;
wire            n566;
wire      [7:0] n567;
wire            n568;
wire      [7:0] n569;
wire            n57;
wire            n570;
wire      [7:0] n571;
wire            n572;
wire      [7:0] n573;
wire            n574;
wire      [7:0] n576;
wire            n578;
wire      [7:0] n579;
wire            n581;
wire      [7:0] n583;
wire            n584;
wire      [7:0] n585;
wire            n586;
wire      [7:0] n587;
wire            n588;
wire      [7:0] n589;
wire      [7:0] n59;
wire            n590;
wire      [7:0] n592;
wire            n593;
wire      [7:0] n594;
wire            n595;
wire      [7:0] n597;
wire            n598;
wire      [7:0] n599;
wire            n600;
wire      [7:0] n601;
wire            n602;
wire      [7:0] n604;
wire            n605;
wire      [7:0] n606;
wire            n608;
wire      [7:0] n609;
wire            n61;
wire            n610;
wire      [7:0] n611;
wire            n612;
wire      [7:0] n613;
wire            n614;
wire      [7:0] n616;
wire            n617;
wire      [7:0] n619;
wire            n620;
wire      [7:0] n622;
wire            n623;
wire      [7:0] n624;
wire            n625;
wire      [7:0] n627;
wire            n629;
wire      [7:0] n63;
wire      [7:0] n630;
wire            n631;
wire      [7:0] n632;
wire            n633;
wire      [7:0] n635;
wire            n636;
wire      [7:0] n637;
wire            n638;
wire      [7:0] n639;
wire            n640;
wire      [7:0] n641;
wire            n642;
wire      [7:0] n644;
wire            n645;
wire      [7:0] n647;
wire            n648;
wire      [7:0] n649;
wire            n65;
wire            n651;
wire      [7:0] n653;
wire            n654;
wire      [7:0] n655;
wire            n657;
wire      [7:0] n659;
wire            n660;
wire      [7:0] n661;
wire            n662;
wire      [7:0] n664;
wire            n666;
wire      [7:0] n667;
wire            n669;
wire      [7:0] n67;
wire      [7:0] n671;
wire            n672;
wire      [7:0] n674;
wire            n675;
wire      [7:0] n676;
wire            n677;
wire      [7:0] n678;
wire            n679;
wire      [7:0] n680;
wire            n682;
wire      [7:0] n683;
wire            n684;
wire      [7:0] n685;
wire            n686;
wire      [7:0] n687;
wire            n688;
wire      [7:0] n689;
wire            n69;
wire            n690;
wire      [7:0] n691;
wire            n693;
wire      [7:0] n694;
wire            n695;
wire      [7:0] n696;
wire            n697;
wire      [7:0] n698;
wire            n699;
wire      [7:0] n7;
wire      [7:0] n700;
wire            n701;
wire      [7:0] n702;
wire            n703;
wire      [7:0] n704;
wire            n705;
wire      [7:0] n706;
wire            n707;
wire      [7:0] n708;
wire            n709;
wire      [7:0] n71;
wire      [7:0] n710;
wire            n711;
wire      [7:0] n712;
wire            n713;
wire      [7:0] n714;
wire            n715;
wire      [7:0] n716;
wire            n717;
wire      [7:0] n718;
wire            n719;
wire      [7:0] n720;
wire            n721;
wire      [7:0] n722;
wire            n723;
wire      [7:0] n724;
wire            n725;
wire      [7:0] n726;
wire            n727;
wire      [7:0] n728;
wire            n729;
wire            n73;
wire      [7:0] n730;
wire            n731;
wire      [7:0] n732;
wire            n733;
wire      [7:0] n734;
wire            n735;
wire      [7:0] n736;
wire            n737;
wire      [7:0] n738;
wire            n739;
wire      [7:0] n740;
wire            n741;
wire      [7:0] n742;
wire            n743;
wire      [7:0] n744;
wire            n745;
wire      [7:0] n746;
wire            n747;
wire      [7:0] n748;
wire            n749;
wire      [7:0] n75;
wire      [7:0] n750;
wire            n751;
wire      [7:0] n753;
wire            n754;
wire      [7:0] n755;
wire            n756;
wire      [7:0] n757;
wire            n758;
wire      [7:0] n759;
wire            n760;
wire      [7:0] n761;
wire            n762;
wire      [7:0] n763;
wire            n764;
wire      [7:0] n765;
wire            n766;
wire      [7:0] n767;
wire            n768;
wire      [7:0] n769;
wire            n77;
wire            n770;
wire      [7:0] n771;
wire      [7:0] n772;
wire      [7:0] n773;
wire      [7:0] n774;
wire      [7:0] n775;
wire      [7:0] n776;
wire      [7:0] n777;
wire      [7:0] n778;
wire      [7:0] n779;
wire      [7:0] n780;
wire      [7:0] n781;
wire      [7:0] n782;
wire      [7:0] n783;
wire      [7:0] n784;
wire      [7:0] n785;
wire      [7:0] n786;
wire      [7:0] n787;
wire      [7:0] n788;
wire      [7:0] n789;
wire      [7:0] n79;
wire      [7:0] n790;
wire      [7:0] n791;
wire      [7:0] n792;
wire      [7:0] n793;
wire      [7:0] n794;
wire      [7:0] n795;
wire      [7:0] n796;
wire      [7:0] n797;
wire      [7:0] n798;
wire      [7:0] n799;
wire      [7:0] n800;
wire      [7:0] n801;
wire      [7:0] n802;
wire      [7:0] n803;
wire      [7:0] n804;
wire      [7:0] n805;
wire      [7:0] n806;
wire      [7:0] n807;
wire      [7:0] n808;
wire      [7:0] n809;
wire            n81;
wire      [7:0] n810;
wire      [7:0] n811;
wire      [7:0] n812;
wire      [7:0] n813;
wire      [7:0] n814;
wire      [7:0] n815;
wire      [7:0] n816;
wire      [7:0] n817;
wire      [7:0] n818;
wire      [7:0] n819;
wire      [7:0] n820;
wire      [7:0] n821;
wire      [7:0] n822;
wire      [7:0] n823;
wire      [7:0] n824;
wire      [7:0] n825;
wire      [7:0] n826;
wire      [7:0] n827;
wire      [7:0] n828;
wire      [7:0] n829;
wire      [7:0] n83;
wire      [7:0] n830;
wire      [7:0] n831;
wire      [7:0] n832;
wire      [7:0] n833;
wire      [7:0] n834;
wire      [7:0] n835;
wire      [7:0] n836;
wire      [7:0] n837;
wire      [7:0] n838;
wire      [7:0] n839;
wire      [7:0] n840;
wire      [7:0] n841;
wire      [7:0] n842;
wire      [7:0] n843;
wire      [7:0] n844;
wire      [7:0] n845;
wire      [7:0] n846;
wire      [7:0] n847;
wire      [7:0] n848;
wire      [7:0] n849;
wire            n85;
wire      [7:0] n850;
wire      [7:0] n851;
wire      [7:0] n852;
wire      [7:0] n853;
wire      [7:0] n854;
wire      [7:0] n855;
wire      [7:0] n856;
wire      [7:0] n857;
wire      [7:0] n858;
wire      [7:0] n859;
wire      [7:0] n860;
wire      [7:0] n861;
wire      [7:0] n862;
wire      [7:0] n863;
wire      [7:0] n864;
wire      [7:0] n865;
wire      [7:0] n866;
wire      [7:0] n867;
wire      [7:0] n868;
wire      [7:0] n869;
wire      [7:0] n87;
wire      [7:0] n870;
wire      [7:0] n871;
wire      [7:0] n872;
wire      [7:0] n873;
wire      [7:0] n874;
wire      [7:0] n875;
wire      [7:0] n876;
wire      [7:0] n877;
wire      [7:0] n878;
wire      [7:0] n879;
wire      [7:0] n880;
wire      [7:0] n881;
wire      [7:0] n882;
wire      [7:0] n883;
wire      [7:0] n884;
wire      [7:0] n885;
wire      [7:0] n886;
wire      [7:0] n887;
wire      [7:0] n888;
wire      [7:0] n889;
wire            n89;
wire      [7:0] n890;
wire      [7:0] n891;
wire      [7:0] n892;
wire      [7:0] n893;
wire      [7:0] n894;
wire      [7:0] n895;
wire      [7:0] n896;
wire      [7:0] n897;
wire      [7:0] n898;
wire      [7:0] n899;
wire            n9;
wire      [7:0] n900;
wire      [7:0] n901;
wire      [7:0] n902;
wire      [7:0] n903;
wire      [7:0] n904;
wire      [7:0] n905;
wire      [7:0] n906;
wire      [7:0] n907;
wire      [7:0] n908;
wire      [7:0] n909;
wire      [7:0] n91;
wire      [7:0] n910;
wire      [7:0] n911;
wire      [7:0] n912;
wire      [7:0] n913;
wire      [7:0] n914;
wire      [7:0] n915;
wire      [7:0] n916;
wire      [7:0] n917;
wire      [7:0] n918;
wire      [7:0] n919;
wire            n92;
wire      [7:0] n920;
wire      [7:0] n921;
wire      [7:0] n922;
wire      [7:0] n923;
wire      [7:0] n924;
wire      [7:0] n925;
wire      [7:0] n926;
wire      [7:0] n927;
wire      [7:0] n928;
wire      [7:0] n929;
wire      [7:0] n930;
wire      [7:0] n931;
wire      [7:0] n932;
wire      [7:0] n933;
wire      [7:0] n934;
wire      [7:0] n935;
wire      [7:0] n936;
wire      [7:0] n937;
wire      [7:0] n938;
wire      [7:0] n939;
wire      [7:0] n94;
wire      [7:0] n940;
wire      [7:0] n941;
wire      [7:0] n942;
wire      [7:0] n943;
wire      [7:0] n944;
wire      [7:0] n945;
wire      [7:0] n946;
wire      [7:0] n947;
wire      [7:0] n948;
wire      [7:0] n949;
wire      [7:0] n950;
wire      [7:0] n951;
wire      [7:0] n952;
wire      [7:0] n953;
wire      [7:0] n954;
wire      [7:0] n955;
wire      [7:0] n956;
wire      [7:0] n957;
wire      [7:0] n958;
wire      [7:0] n959;
wire            n96;
wire      [7:0] n960;
wire      [7:0] n961;
wire      [7:0] n962;
wire      [7:0] n963;
wire      [7:0] n964;
wire      [7:0] n965;
wire      [7:0] n966;
wire      [7:0] n967;
wire      [7:0] n968;
wire      [7:0] n969;
wire      [7:0] n970;
wire      [7:0] n971;
wire      [7:0] n972;
wire      [7:0] n973;
wire      [7:0] n974;
wire      [7:0] n975;
wire      [7:0] n976;
wire      [7:0] n977;
wire      [7:0] n978;
wire      [7:0] n979;
wire      [7:0] n98;
wire      [7:0] n980;
wire      [7:0] n981;
wire      [7:0] n982;
wire      [7:0] n983;
wire      [7:0] n984;
wire      [7:0] n985;
wire      [7:0] n986;
wire      [7:0] n987;
wire      [7:0] n988;
wire      [7:0] n989;
wire      [7:0] n990;
wire      [7:0] n991;
wire      [7:0] n992;
wire      [7:0] n993;
wire      [7:0] n994;
wire      [7:0] n995;
wire      [7:0] n996;
wire      [7:0] n997;
wire      [7:0] n998;
wire      [7:0] n999;
(* keep *) wire    [127:0] out_1_randinit;
(* keep *) wire      [7:0] rcon_randinit;
wire            rst;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign n1 = in[127:120] ;
assign n2 =  ( n1 ) ^ ( rcon )  ;
assign n3 = in[23:16] ;
assign bv_8_255_n4 = 8'hff ;
assign n5 =  ( n3 ) == ( bv_8_255_n4 )  ;
assign bv_8_22_n6 = 8'h16 ;
assign n7 = in[23:16] ;
assign bv_8_254_n8 = 8'hfe ;
assign n9 =  ( n7 ) == ( bv_8_254_n8 )  ;
assign bv_8_187_n10 = 8'hbb ;
assign n11 = in[23:16] ;
assign bv_8_253_n12 = 8'hfd ;
assign n13 =  ( n11 ) == ( bv_8_253_n12 )  ;
assign bv_8_84_n14 = 8'h54 ;
assign n15 = in[23:16] ;
assign bv_8_252_n16 = 8'hfc ;
assign n17 =  ( n15 ) == ( bv_8_252_n16 )  ;
assign bv_8_176_n18 = 8'hb0 ;
assign n19 = in[23:16] ;
assign bv_8_251_n20 = 8'hfb ;
assign n21 =  ( n19 ) == ( bv_8_251_n20 )  ;
assign bv_8_15_n22 = 8'hf ;
assign n23 = in[23:16] ;
assign bv_8_250_n24 = 8'hfa ;
assign n25 =  ( n23 ) == ( bv_8_250_n24 )  ;
assign bv_8_45_n26 = 8'h2d ;
assign n27 = in[23:16] ;
assign bv_8_249_n28 = 8'hf9 ;
assign n29 =  ( n27 ) == ( bv_8_249_n28 )  ;
assign bv_8_153_n30 = 8'h99 ;
assign n31 = in[23:16] ;
assign bv_8_248_n32 = 8'hf8 ;
assign n33 =  ( n31 ) == ( bv_8_248_n32 )  ;
assign bv_8_65_n34 = 8'h41 ;
assign n35 = in[23:16] ;
assign bv_8_247_n36 = 8'hf7 ;
assign n37 =  ( n35 ) == ( bv_8_247_n36 )  ;
assign bv_8_104_n38 = 8'h68 ;
assign n39 = in[23:16] ;
assign bv_8_246_n40 = 8'hf6 ;
assign n41 =  ( n39 ) == ( bv_8_246_n40 )  ;
assign bv_8_66_n42 = 8'h42 ;
assign n43 = in[23:16] ;
assign bv_8_245_n44 = 8'hf5 ;
assign n45 =  ( n43 ) == ( bv_8_245_n44 )  ;
assign bv_8_230_n46 = 8'he6 ;
assign n47 = in[23:16] ;
assign bv_8_244_n48 = 8'hf4 ;
assign n49 =  ( n47 ) == ( bv_8_244_n48 )  ;
assign bv_8_191_n50 = 8'hbf ;
assign n51 = in[23:16] ;
assign bv_8_243_n52 = 8'hf3 ;
assign n53 =  ( n51 ) == ( bv_8_243_n52 )  ;
assign bv_8_13_n54 = 8'hd ;
assign n55 = in[23:16] ;
assign bv_8_242_n56 = 8'hf2 ;
assign n57 =  ( n55 ) == ( bv_8_242_n56 )  ;
assign bv_8_137_n58 = 8'h89 ;
assign n59 = in[23:16] ;
assign bv_8_241_n60 = 8'hf1 ;
assign n61 =  ( n59 ) == ( bv_8_241_n60 )  ;
assign bv_8_161_n62 = 8'ha1 ;
assign n63 = in[23:16] ;
assign bv_8_240_n64 = 8'hf0 ;
assign n65 =  ( n63 ) == ( bv_8_240_n64 )  ;
assign bv_8_140_n66 = 8'h8c ;
assign n67 = in[23:16] ;
assign bv_8_239_n68 = 8'hef ;
assign n69 =  ( n67 ) == ( bv_8_239_n68 )  ;
assign bv_8_223_n70 = 8'hdf ;
assign n71 = in[23:16] ;
assign bv_8_238_n72 = 8'hee ;
assign n73 =  ( n71 ) == ( bv_8_238_n72 )  ;
assign bv_8_40_n74 = 8'h28 ;
assign n75 = in[23:16] ;
assign bv_8_237_n76 = 8'hed ;
assign n77 =  ( n75 ) == ( bv_8_237_n76 )  ;
assign bv_8_85_n78 = 8'h55 ;
assign n79 = in[23:16] ;
assign bv_8_236_n80 = 8'hec ;
assign n81 =  ( n79 ) == ( bv_8_236_n80 )  ;
assign bv_8_206_n82 = 8'hce ;
assign n83 = in[23:16] ;
assign bv_8_235_n84 = 8'heb ;
assign n85 =  ( n83 ) == ( bv_8_235_n84 )  ;
assign bv_8_233_n86 = 8'he9 ;
assign n87 = in[23:16] ;
assign bv_8_234_n88 = 8'hea ;
assign n89 =  ( n87 ) == ( bv_8_234_n88 )  ;
assign bv_8_135_n90 = 8'h87 ;
assign n91 = in[23:16] ;
assign n92 =  ( n91 ) == ( bv_8_233_n86 )  ;
assign bv_8_30_n93 = 8'h1e ;
assign n94 = in[23:16] ;
assign bv_8_232_n95 = 8'he8 ;
assign n96 =  ( n94 ) == ( bv_8_232_n95 )  ;
assign bv_8_155_n97 = 8'h9b ;
assign n98 = in[23:16] ;
assign bv_8_231_n99 = 8'he7 ;
assign n100 =  ( n98 ) == ( bv_8_231_n99 )  ;
assign bv_8_148_n101 = 8'h94 ;
assign n102 = in[23:16] ;
assign n103 =  ( n102 ) == ( bv_8_230_n46 )  ;
assign bv_8_142_n104 = 8'h8e ;
assign n105 = in[23:16] ;
assign bv_8_229_n106 = 8'he5 ;
assign n107 =  ( n105 ) == ( bv_8_229_n106 )  ;
assign bv_8_217_n108 = 8'hd9 ;
assign n109 = in[23:16] ;
assign bv_8_228_n110 = 8'he4 ;
assign n111 =  ( n109 ) == ( bv_8_228_n110 )  ;
assign bv_8_105_n112 = 8'h69 ;
assign n113 = in[23:16] ;
assign bv_8_227_n114 = 8'he3 ;
assign n115 =  ( n113 ) == ( bv_8_227_n114 )  ;
assign bv_8_17_n116 = 8'h11 ;
assign n117 = in[23:16] ;
assign bv_8_226_n118 = 8'he2 ;
assign n119 =  ( n117 ) == ( bv_8_226_n118 )  ;
assign bv_8_152_n120 = 8'h98 ;
assign n121 = in[23:16] ;
assign bv_8_225_n122 = 8'he1 ;
assign n123 =  ( n121 ) == ( bv_8_225_n122 )  ;
assign n124 = in[23:16] ;
assign bv_8_224_n125 = 8'he0 ;
assign n126 =  ( n124 ) == ( bv_8_224_n125 )  ;
assign n127 = in[23:16] ;
assign n128 =  ( n127 ) == ( bv_8_223_n70 )  ;
assign bv_8_158_n129 = 8'h9e ;
assign n130 = in[23:16] ;
assign bv_8_222_n131 = 8'hde ;
assign n132 =  ( n130 ) == ( bv_8_222_n131 )  ;
assign bv_8_29_n133 = 8'h1d ;
assign n134 = in[23:16] ;
assign bv_8_221_n135 = 8'hdd ;
assign n136 =  ( n134 ) == ( bv_8_221_n135 )  ;
assign bv_8_193_n137 = 8'hc1 ;
assign n138 = in[23:16] ;
assign bv_8_220_n139 = 8'hdc ;
assign n140 =  ( n138 ) == ( bv_8_220_n139 )  ;
assign bv_8_134_n141 = 8'h86 ;
assign n142 = in[23:16] ;
assign bv_8_219_n143 = 8'hdb ;
assign n144 =  ( n142 ) == ( bv_8_219_n143 )  ;
assign bv_8_185_n145 = 8'hb9 ;
assign n146 = in[23:16] ;
assign bv_8_218_n147 = 8'hda ;
assign n148 =  ( n146 ) == ( bv_8_218_n147 )  ;
assign bv_8_87_n149 = 8'h57 ;
assign n150 = in[23:16] ;
assign n151 =  ( n150 ) == ( bv_8_217_n108 )  ;
assign bv_8_53_n152 = 8'h35 ;
assign n153 = in[23:16] ;
assign bv_8_216_n154 = 8'hd8 ;
assign n155 =  ( n153 ) == ( bv_8_216_n154 )  ;
assign bv_8_97_n156 = 8'h61 ;
assign n157 = in[23:16] ;
assign bv_8_215_n158 = 8'hd7 ;
assign n159 =  ( n157 ) == ( bv_8_215_n158 )  ;
assign bv_8_14_n160 = 8'he ;
assign n161 = in[23:16] ;
assign bv_8_214_n162 = 8'hd6 ;
assign n163 =  ( n161 ) == ( bv_8_214_n162 )  ;
assign n164 = in[23:16] ;
assign bv_8_213_n165 = 8'hd5 ;
assign n166 =  ( n164 ) == ( bv_8_213_n165 )  ;
assign bv_8_3_n167 = 8'h3 ;
assign n168 = in[23:16] ;
assign bv_8_212_n169 = 8'hd4 ;
assign n170 =  ( n168 ) == ( bv_8_212_n169 )  ;
assign bv_8_72_n171 = 8'h48 ;
assign n172 = in[23:16] ;
assign bv_8_211_n173 = 8'hd3 ;
assign n174 =  ( n172 ) == ( bv_8_211_n173 )  ;
assign bv_8_102_n175 = 8'h66 ;
assign n176 = in[23:16] ;
assign bv_8_210_n177 = 8'hd2 ;
assign n178 =  ( n176 ) == ( bv_8_210_n177 )  ;
assign bv_8_181_n179 = 8'hb5 ;
assign n180 = in[23:16] ;
assign bv_8_209_n181 = 8'hd1 ;
assign n182 =  ( n180 ) == ( bv_8_209_n181 )  ;
assign bv_8_62_n183 = 8'h3e ;
assign n184 = in[23:16] ;
assign bv_8_208_n185 = 8'hd0 ;
assign n186 =  ( n184 ) == ( bv_8_208_n185 )  ;
assign bv_8_112_n187 = 8'h70 ;
assign n188 = in[23:16] ;
assign bv_8_207_n189 = 8'hcf ;
assign n190 =  ( n188 ) == ( bv_8_207_n189 )  ;
assign bv_8_138_n191 = 8'h8a ;
assign n192 = in[23:16] ;
assign n193 =  ( n192 ) == ( bv_8_206_n82 )  ;
assign bv_8_139_n194 = 8'h8b ;
assign n195 = in[23:16] ;
assign bv_8_205_n196 = 8'hcd ;
assign n197 =  ( n195 ) == ( bv_8_205_n196 )  ;
assign bv_8_189_n198 = 8'hbd ;
assign n199 = in[23:16] ;
assign bv_8_204_n200 = 8'hcc ;
assign n201 =  ( n199 ) == ( bv_8_204_n200 )  ;
assign bv_8_75_n202 = 8'h4b ;
assign n203 = in[23:16] ;
assign bv_8_203_n204 = 8'hcb ;
assign n205 =  ( n203 ) == ( bv_8_203_n204 )  ;
assign bv_8_31_n206 = 8'h1f ;
assign n207 = in[23:16] ;
assign bv_8_202_n208 = 8'hca ;
assign n209 =  ( n207 ) == ( bv_8_202_n208 )  ;
assign bv_8_116_n210 = 8'h74 ;
assign n211 = in[23:16] ;
assign bv_8_201_n212 = 8'hc9 ;
assign n213 =  ( n211 ) == ( bv_8_201_n212 )  ;
assign n214 = in[23:16] ;
assign bv_8_200_n215 = 8'hc8 ;
assign n216 =  ( n214 ) == ( bv_8_200_n215 )  ;
assign n217 = in[23:16] ;
assign bv_8_199_n218 = 8'hc7 ;
assign n219 =  ( n217 ) == ( bv_8_199_n218 )  ;
assign bv_8_198_n220 = 8'hc6 ;
assign n221 = in[23:16] ;
assign n222 =  ( n221 ) == ( bv_8_198_n220 )  ;
assign bv_8_180_n223 = 8'hb4 ;
assign n224 = in[23:16] ;
assign bv_8_197_n225 = 8'hc5 ;
assign n226 =  ( n224 ) == ( bv_8_197_n225 )  ;
assign bv_8_166_n227 = 8'ha6 ;
assign n228 = in[23:16] ;
assign bv_8_196_n229 = 8'hc4 ;
assign n230 =  ( n228 ) == ( bv_8_196_n229 )  ;
assign bv_8_28_n231 = 8'h1c ;
assign n232 = in[23:16] ;
assign bv_8_195_n233 = 8'hc3 ;
assign n234 =  ( n232 ) == ( bv_8_195_n233 )  ;
assign bv_8_46_n235 = 8'h2e ;
assign n236 = in[23:16] ;
assign bv_8_194_n237 = 8'hc2 ;
assign n238 =  ( n236 ) == ( bv_8_194_n237 )  ;
assign bv_8_37_n239 = 8'h25 ;
assign n240 = in[23:16] ;
assign n241 =  ( n240 ) == ( bv_8_193_n137 )  ;
assign bv_8_120_n242 = 8'h78 ;
assign n243 = in[23:16] ;
assign bv_8_192_n244 = 8'hc0 ;
assign n245 =  ( n243 ) == ( bv_8_192_n244 )  ;
assign bv_8_186_n246 = 8'hba ;
assign n247 = in[23:16] ;
assign n248 =  ( n247 ) == ( bv_8_191_n50 )  ;
assign bv_8_8_n249 = 8'h8 ;
assign n250 = in[23:16] ;
assign bv_8_190_n251 = 8'hbe ;
assign n252 =  ( n250 ) == ( bv_8_190_n251 )  ;
assign bv_8_174_n253 = 8'hae ;
assign n254 = in[23:16] ;
assign n255 =  ( n254 ) == ( bv_8_189_n198 )  ;
assign bv_8_122_n256 = 8'h7a ;
assign n257 = in[23:16] ;
assign bv_8_188_n258 = 8'hbc ;
assign n259 =  ( n257 ) == ( bv_8_188_n258 )  ;
assign bv_8_101_n260 = 8'h65 ;
assign n261 = in[23:16] ;
assign n262 =  ( n261 ) == ( bv_8_187_n10 )  ;
assign n263 = in[23:16] ;
assign n264 =  ( n263 ) == ( bv_8_186_n246 )  ;
assign n265 = in[23:16] ;
assign n266 =  ( n265 ) == ( bv_8_185_n145 )  ;
assign bv_8_86_n267 = 8'h56 ;
assign n268 = in[23:16] ;
assign bv_8_184_n269 = 8'hb8 ;
assign n270 =  ( n268 ) == ( bv_8_184_n269 )  ;
assign bv_8_108_n271 = 8'h6c ;
assign n272 = in[23:16] ;
assign bv_8_183_n273 = 8'hb7 ;
assign n274 =  ( n272 ) == ( bv_8_183_n273 )  ;
assign bv_8_169_n275 = 8'ha9 ;
assign n276 = in[23:16] ;
assign bv_8_182_n277 = 8'hb6 ;
assign n278 =  ( n276 ) == ( bv_8_182_n277 )  ;
assign bv_8_78_n279 = 8'h4e ;
assign n280 = in[23:16] ;
assign n281 =  ( n280 ) == ( bv_8_181_n179 )  ;
assign n282 = in[23:16] ;
assign n283 =  ( n282 ) == ( bv_8_180_n223 )  ;
assign bv_8_141_n284 = 8'h8d ;
assign n285 = in[23:16] ;
assign bv_8_179_n286 = 8'hb3 ;
assign n287 =  ( n285 ) == ( bv_8_179_n286 )  ;
assign bv_8_109_n288 = 8'h6d ;
assign n289 = in[23:16] ;
assign bv_8_178_n290 = 8'hb2 ;
assign n291 =  ( n289 ) == ( bv_8_178_n290 )  ;
assign bv_8_55_n292 = 8'h37 ;
assign n293 = in[23:16] ;
assign bv_8_177_n294 = 8'hb1 ;
assign n295 =  ( n293 ) == ( bv_8_177_n294 )  ;
assign n296 = in[23:16] ;
assign n297 =  ( n296 ) == ( bv_8_176_n18 )  ;
assign n298 = in[23:16] ;
assign bv_8_175_n299 = 8'haf ;
assign n300 =  ( n298 ) == ( bv_8_175_n299 )  ;
assign bv_8_121_n301 = 8'h79 ;
assign n302 = in[23:16] ;
assign n303 =  ( n302 ) == ( bv_8_174_n253 )  ;
assign n304 = in[23:16] ;
assign bv_8_173_n305 = 8'had ;
assign n306 =  ( n304 ) == ( bv_8_173_n305 )  ;
assign bv_8_149_n307 = 8'h95 ;
assign n308 = in[23:16] ;
assign bv_8_172_n309 = 8'hac ;
assign n310 =  ( n308 ) == ( bv_8_172_n309 )  ;
assign bv_8_145_n311 = 8'h91 ;
assign n312 = in[23:16] ;
assign bv_8_171_n313 = 8'hab ;
assign n314 =  ( n312 ) == ( bv_8_171_n313 )  ;
assign bv_8_98_n315 = 8'h62 ;
assign n316 = in[23:16] ;
assign bv_8_170_n317 = 8'haa ;
assign n318 =  ( n316 ) == ( bv_8_170_n317 )  ;
assign n319 = in[23:16] ;
assign n320 =  ( n319 ) == ( bv_8_169_n275 )  ;
assign n321 = in[23:16] ;
assign bv_8_168_n322 = 8'ha8 ;
assign n323 =  ( n321 ) == ( bv_8_168_n322 )  ;
assign n324 = in[23:16] ;
assign bv_8_167_n325 = 8'ha7 ;
assign n326 =  ( n324 ) == ( bv_8_167_n325 )  ;
assign bv_8_92_n327 = 8'h5c ;
assign n328 = in[23:16] ;
assign n329 =  ( n328 ) == ( bv_8_166_n227 )  ;
assign bv_8_36_n330 = 8'h24 ;
assign n331 = in[23:16] ;
assign bv_8_165_n332 = 8'ha5 ;
assign n333 =  ( n331 ) == ( bv_8_165_n332 )  ;
assign bv_8_6_n334 = 8'h6 ;
assign n335 = in[23:16] ;
assign bv_8_164_n336 = 8'ha4 ;
assign n337 =  ( n335 ) == ( bv_8_164_n336 )  ;
assign bv_8_73_n338 = 8'h49 ;
assign n339 = in[23:16] ;
assign bv_8_163_n340 = 8'ha3 ;
assign n341 =  ( n339 ) == ( bv_8_163_n340 )  ;
assign bv_8_10_n342 = 8'ha ;
assign n343 = in[23:16] ;
assign bv_8_162_n344 = 8'ha2 ;
assign n345 =  ( n343 ) == ( bv_8_162_n344 )  ;
assign bv_8_58_n346 = 8'h3a ;
assign n347 = in[23:16] ;
assign n348 =  ( n347 ) == ( bv_8_161_n62 )  ;
assign bv_8_50_n349 = 8'h32 ;
assign n350 = in[23:16] ;
assign bv_8_160_n351 = 8'ha0 ;
assign n352 =  ( n350 ) == ( bv_8_160_n351 )  ;
assign n353 = in[23:16] ;
assign bv_8_159_n354 = 8'h9f ;
assign n355 =  ( n353 ) == ( bv_8_159_n354 )  ;
assign n356 = in[23:16] ;
assign n357 =  ( n356 ) == ( bv_8_158_n129 )  ;
assign bv_8_11_n358 = 8'hb ;
assign n359 = in[23:16] ;
assign bv_8_157_n360 = 8'h9d ;
assign n361 =  ( n359 ) == ( bv_8_157_n360 )  ;
assign bv_8_94_n362 = 8'h5e ;
assign n363 = in[23:16] ;
assign bv_8_156_n364 = 8'h9c ;
assign n365 =  ( n363 ) == ( bv_8_156_n364 )  ;
assign n366 = in[23:16] ;
assign n367 =  ( n366 ) == ( bv_8_155_n97 )  ;
assign bv_8_20_n368 = 8'h14 ;
assign n369 = in[23:16] ;
assign bv_8_154_n370 = 8'h9a ;
assign n371 =  ( n369 ) == ( bv_8_154_n370 )  ;
assign n372 = in[23:16] ;
assign n373 =  ( n372 ) == ( bv_8_153_n30 )  ;
assign n374 = in[23:16] ;
assign n375 =  ( n374 ) == ( bv_8_152_n120 )  ;
assign bv_8_70_n376 = 8'h46 ;
assign n377 = in[23:16] ;
assign bv_8_151_n378 = 8'h97 ;
assign n379 =  ( n377 ) == ( bv_8_151_n378 )  ;
assign bv_8_136_n380 = 8'h88 ;
assign n381 = in[23:16] ;
assign bv_8_150_n382 = 8'h96 ;
assign n383 =  ( n381 ) == ( bv_8_150_n382 )  ;
assign bv_8_144_n384 = 8'h90 ;
assign n385 = in[23:16] ;
assign n386 =  ( n385 ) == ( bv_8_149_n307 )  ;
assign bv_8_42_n387 = 8'h2a ;
assign n388 = in[23:16] ;
assign n389 =  ( n388 ) == ( bv_8_148_n101 )  ;
assign bv_8_34_n390 = 8'h22 ;
assign n391 = in[23:16] ;
assign bv_8_147_n392 = 8'h93 ;
assign n393 =  ( n391 ) == ( bv_8_147_n392 )  ;
assign n394 = in[23:16] ;
assign bv_8_146_n395 = 8'h92 ;
assign n396 =  ( n394 ) == ( bv_8_146_n395 )  ;
assign bv_8_79_n397 = 8'h4f ;
assign n398 = in[23:16] ;
assign n399 =  ( n398 ) == ( bv_8_145_n311 )  ;
assign bv_8_129_n400 = 8'h81 ;
assign n401 = in[23:16] ;
assign n402 =  ( n401 ) == ( bv_8_144_n384 )  ;
assign bv_8_96_n403 = 8'h60 ;
assign n404 = in[23:16] ;
assign bv_8_143_n405 = 8'h8f ;
assign n406 =  ( n404 ) == ( bv_8_143_n405 )  ;
assign bv_8_115_n407 = 8'h73 ;
assign n408 = in[23:16] ;
assign n409 =  ( n408 ) == ( bv_8_142_n104 )  ;
assign bv_8_25_n410 = 8'h19 ;
assign n411 = in[23:16] ;
assign n412 =  ( n411 ) == ( bv_8_141_n284 )  ;
assign bv_8_93_n413 = 8'h5d ;
assign n414 = in[23:16] ;
assign n415 =  ( n414 ) == ( bv_8_140_n66 )  ;
assign bv_8_100_n416 = 8'h64 ;
assign n417 = in[23:16] ;
assign n418 =  ( n417 ) == ( bv_8_139_n194 )  ;
assign bv_8_61_n419 = 8'h3d ;
assign n420 = in[23:16] ;
assign n421 =  ( n420 ) == ( bv_8_138_n191 )  ;
assign bv_8_126_n422 = 8'h7e ;
assign n423 = in[23:16] ;
assign n424 =  ( n423 ) == ( bv_8_137_n58 )  ;
assign n425 = in[23:16] ;
assign n426 =  ( n425 ) == ( bv_8_136_n380 )  ;
assign n427 = in[23:16] ;
assign n428 =  ( n427 ) == ( bv_8_135_n90 )  ;
assign bv_8_23_n429 = 8'h17 ;
assign n430 = in[23:16] ;
assign n431 =  ( n430 ) == ( bv_8_134_n141 )  ;
assign bv_8_68_n432 = 8'h44 ;
assign n433 = in[23:16] ;
assign bv_8_133_n434 = 8'h85 ;
assign n435 =  ( n433 ) == ( bv_8_133_n434 )  ;
assign n436 = in[23:16] ;
assign bv_8_132_n437 = 8'h84 ;
assign n438 =  ( n436 ) == ( bv_8_132_n437 )  ;
assign bv_8_95_n439 = 8'h5f ;
assign n440 = in[23:16] ;
assign bv_8_131_n441 = 8'h83 ;
assign n442 =  ( n440 ) == ( bv_8_131_n441 )  ;
assign n443 = in[23:16] ;
assign bv_8_130_n444 = 8'h82 ;
assign n445 =  ( n443 ) == ( bv_8_130_n444 )  ;
assign bv_8_19_n446 = 8'h13 ;
assign n447 = in[23:16] ;
assign n448 =  ( n447 ) == ( bv_8_129_n400 )  ;
assign bv_8_12_n449 = 8'hc ;
assign n450 = in[23:16] ;
assign bv_8_128_n451 = 8'h80 ;
assign n452 =  ( n450 ) == ( bv_8_128_n451 )  ;
assign n453 = in[23:16] ;
assign bv_8_127_n454 = 8'h7f ;
assign n455 =  ( n453 ) == ( bv_8_127_n454 )  ;
assign n456 = in[23:16] ;
assign n457 =  ( n456 ) == ( bv_8_126_n422 )  ;
assign n458 = in[23:16] ;
assign bv_8_125_n459 = 8'h7d ;
assign n460 =  ( n458 ) == ( bv_8_125_n459 )  ;
assign n461 = in[23:16] ;
assign bv_8_124_n462 = 8'h7c ;
assign n463 =  ( n461 ) == ( bv_8_124_n462 )  ;
assign bv_8_16_n464 = 8'h10 ;
assign n465 = in[23:16] ;
assign bv_8_123_n466 = 8'h7b ;
assign n467 =  ( n465 ) == ( bv_8_123_n466 )  ;
assign bv_8_33_n468 = 8'h21 ;
assign n469 = in[23:16] ;
assign n470 =  ( n469 ) == ( bv_8_122_n256 )  ;
assign n471 = in[23:16] ;
assign n472 =  ( n471 ) == ( bv_8_121_n301 )  ;
assign n473 = in[23:16] ;
assign n474 =  ( n473 ) == ( bv_8_120_n242 )  ;
assign n475 = in[23:16] ;
assign bv_8_119_n476 = 8'h77 ;
assign n477 =  ( n475 ) == ( bv_8_119_n476 )  ;
assign n478 = in[23:16] ;
assign bv_8_118_n479 = 8'h76 ;
assign n480 =  ( n478 ) == ( bv_8_118_n479 )  ;
assign bv_8_56_n481 = 8'h38 ;
assign n482 = in[23:16] ;
assign bv_8_117_n483 = 8'h75 ;
assign n484 =  ( n482 ) == ( bv_8_117_n483 )  ;
assign n485 = in[23:16] ;
assign n486 =  ( n485 ) == ( bv_8_116_n210 )  ;
assign n487 = in[23:16] ;
assign n488 =  ( n487 ) == ( bv_8_115_n407 )  ;
assign n489 = in[23:16] ;
assign bv_8_114_n490 = 8'h72 ;
assign n491 =  ( n489 ) == ( bv_8_114_n490 )  ;
assign bv_8_64_n492 = 8'h40 ;
assign n493 = in[23:16] ;
assign bv_8_113_n494 = 8'h71 ;
assign n495 =  ( n493 ) == ( bv_8_113_n494 )  ;
assign n496 = in[23:16] ;
assign n497 =  ( n496 ) == ( bv_8_112_n187 )  ;
assign bv_8_81_n498 = 8'h51 ;
assign n499 = in[23:16] ;
assign bv_8_111_n500 = 8'h6f ;
assign n501 =  ( n499 ) == ( bv_8_111_n500 )  ;
assign n502 = in[23:16] ;
assign bv_8_110_n503 = 8'h6e ;
assign n504 =  ( n502 ) == ( bv_8_110_n503 )  ;
assign n505 = in[23:16] ;
assign n506 =  ( n505 ) == ( bv_8_109_n288 )  ;
assign bv_8_60_n507 = 8'h3c ;
assign n508 = in[23:16] ;
assign n509 =  ( n508 ) == ( bv_8_108_n271 )  ;
assign bv_8_80_n510 = 8'h50 ;
assign n511 = in[23:16] ;
assign bv_8_107_n512 = 8'h6b ;
assign n513 =  ( n511 ) == ( bv_8_107_n512 )  ;
assign n514 = in[23:16] ;
assign bv_8_106_n515 = 8'h6a ;
assign n516 =  ( n514 ) == ( bv_8_106_n515 )  ;
assign bv_8_2_n517 = 8'h2 ;
assign n518 = in[23:16] ;
assign n519 =  ( n518 ) == ( bv_8_105_n112 )  ;
assign n520 = in[23:16] ;
assign n521 =  ( n520 ) == ( bv_8_104_n38 )  ;
assign bv_8_69_n522 = 8'h45 ;
assign n523 = in[23:16] ;
assign bv_8_103_n524 = 8'h67 ;
assign n525 =  ( n523 ) == ( bv_8_103_n524 )  ;
assign n526 = in[23:16] ;
assign n527 =  ( n526 ) == ( bv_8_102_n175 )  ;
assign bv_8_51_n528 = 8'h33 ;
assign n529 = in[23:16] ;
assign n530 =  ( n529 ) == ( bv_8_101_n260 )  ;
assign bv_8_77_n531 = 8'h4d ;
assign n532 = in[23:16] ;
assign n533 =  ( n532 ) == ( bv_8_100_n416 )  ;
assign bv_8_67_n534 = 8'h43 ;
assign n535 = in[23:16] ;
assign bv_8_99_n536 = 8'h63 ;
assign n537 =  ( n535 ) == ( bv_8_99_n536 )  ;
assign n538 = in[23:16] ;
assign n539 =  ( n538 ) == ( bv_8_98_n315 )  ;
assign n540 = in[23:16] ;
assign n541 =  ( n540 ) == ( bv_8_97_n156 )  ;
assign n542 = in[23:16] ;
assign n543 =  ( n542 ) == ( bv_8_96_n403 )  ;
assign n544 = in[23:16] ;
assign n545 =  ( n544 ) == ( bv_8_95_n439 )  ;
assign n546 = in[23:16] ;
assign n547 =  ( n546 ) == ( bv_8_94_n362 )  ;
assign bv_8_88_n548 = 8'h58 ;
assign n549 = in[23:16] ;
assign n550 =  ( n549 ) == ( bv_8_93_n413 )  ;
assign bv_8_76_n551 = 8'h4c ;
assign n552 = in[23:16] ;
assign n553 =  ( n552 ) == ( bv_8_92_n327 )  ;
assign bv_8_74_n554 = 8'h4a ;
assign n555 = in[23:16] ;
assign bv_8_91_n556 = 8'h5b ;
assign n557 =  ( n555 ) == ( bv_8_91_n556 )  ;
assign bv_8_57_n558 = 8'h39 ;
assign n559 = in[23:16] ;
assign bv_8_90_n560 = 8'h5a ;
assign n561 =  ( n559 ) == ( bv_8_90_n560 )  ;
assign n562 = in[23:16] ;
assign bv_8_89_n563 = 8'h59 ;
assign n564 =  ( n562 ) == ( bv_8_89_n563 )  ;
assign n565 = in[23:16] ;
assign n566 =  ( n565 ) == ( bv_8_88_n548 )  ;
assign n567 = in[23:16] ;
assign n568 =  ( n567 ) == ( bv_8_87_n149 )  ;
assign n569 = in[23:16] ;
assign n570 =  ( n569 ) == ( bv_8_86_n267 )  ;
assign n571 = in[23:16] ;
assign n572 =  ( n571 ) == ( bv_8_85_n78 )  ;
assign n573 = in[23:16] ;
assign n574 =  ( n573 ) == ( bv_8_84_n14 )  ;
assign bv_8_32_n575 = 8'h20 ;
assign n576 = in[23:16] ;
assign bv_8_83_n577 = 8'h53 ;
assign n578 =  ( n576 ) == ( bv_8_83_n577 )  ;
assign n579 = in[23:16] ;
assign bv_8_82_n580 = 8'h52 ;
assign n581 =  ( n579 ) == ( bv_8_82_n580 )  ;
assign bv_8_0_n582 = 8'h0 ;
assign n583 = in[23:16] ;
assign n584 =  ( n583 ) == ( bv_8_81_n498 )  ;
assign n585 = in[23:16] ;
assign n586 =  ( n585 ) == ( bv_8_80_n510 )  ;
assign n587 = in[23:16] ;
assign n588 =  ( n587 ) == ( bv_8_79_n397 )  ;
assign n589 = in[23:16] ;
assign n590 =  ( n589 ) == ( bv_8_78_n279 )  ;
assign bv_8_47_n591 = 8'h2f ;
assign n592 = in[23:16] ;
assign n593 =  ( n592 ) == ( bv_8_77_n531 )  ;
assign n594 = in[23:16] ;
assign n595 =  ( n594 ) == ( bv_8_76_n551 )  ;
assign bv_8_41_n596 = 8'h29 ;
assign n597 = in[23:16] ;
assign n598 =  ( n597 ) == ( bv_8_75_n202 )  ;
assign n599 = in[23:16] ;
assign n600 =  ( n599 ) == ( bv_8_74_n554 )  ;
assign n601 = in[23:16] ;
assign n602 =  ( n601 ) == ( bv_8_73_n338 )  ;
assign bv_8_59_n603 = 8'h3b ;
assign n604 = in[23:16] ;
assign n605 =  ( n604 ) == ( bv_8_72_n171 )  ;
assign n606 = in[23:16] ;
assign bv_8_71_n607 = 8'h47 ;
assign n608 =  ( n606 ) == ( bv_8_71_n607 )  ;
assign n609 = in[23:16] ;
assign n610 =  ( n609 ) == ( bv_8_70_n376 )  ;
assign n611 = in[23:16] ;
assign n612 =  ( n611 ) == ( bv_8_69_n522 )  ;
assign n613 = in[23:16] ;
assign n614 =  ( n613 ) == ( bv_8_68_n432 )  ;
assign bv_8_27_n615 = 8'h1b ;
assign n616 = in[23:16] ;
assign n617 =  ( n616 ) == ( bv_8_67_n534 )  ;
assign bv_8_26_n618 = 8'h1a ;
assign n619 = in[23:16] ;
assign n620 =  ( n619 ) == ( bv_8_66_n42 )  ;
assign bv_8_44_n621 = 8'h2c ;
assign n622 = in[23:16] ;
assign n623 =  ( n622 ) == ( bv_8_65_n34 )  ;
assign n624 = in[23:16] ;
assign n625 =  ( n624 ) == ( bv_8_64_n492 )  ;
assign bv_8_9_n626 = 8'h9 ;
assign n627 = in[23:16] ;
assign bv_8_63_n628 = 8'h3f ;
assign n629 =  ( n627 ) == ( bv_8_63_n628 )  ;
assign n630 = in[23:16] ;
assign n631 =  ( n630 ) == ( bv_8_62_n183 )  ;
assign n632 = in[23:16] ;
assign n633 =  ( n632 ) == ( bv_8_61_n419 )  ;
assign bv_8_39_n634 = 8'h27 ;
assign n635 = in[23:16] ;
assign n636 =  ( n635 ) == ( bv_8_60_n507 )  ;
assign n637 = in[23:16] ;
assign n638 =  ( n637 ) == ( bv_8_59_n603 )  ;
assign n639 = in[23:16] ;
assign n640 =  ( n639 ) == ( bv_8_58_n346 )  ;
assign n641 = in[23:16] ;
assign n642 =  ( n641 ) == ( bv_8_57_n558 )  ;
assign bv_8_18_n643 = 8'h12 ;
assign n644 = in[23:16] ;
assign n645 =  ( n644 ) == ( bv_8_56_n481 )  ;
assign bv_8_7_n646 = 8'h7 ;
assign n647 = in[23:16] ;
assign n648 =  ( n647 ) == ( bv_8_55_n292 )  ;
assign n649 = in[23:16] ;
assign bv_8_54_n650 = 8'h36 ;
assign n651 =  ( n649 ) == ( bv_8_54_n650 )  ;
assign bv_8_5_n652 = 8'h5 ;
assign n653 = in[23:16] ;
assign n654 =  ( n653 ) == ( bv_8_53_n152 )  ;
assign n655 = in[23:16] ;
assign bv_8_52_n656 = 8'h34 ;
assign n657 =  ( n655 ) == ( bv_8_52_n656 )  ;
assign bv_8_24_n658 = 8'h18 ;
assign n659 = in[23:16] ;
assign n660 =  ( n659 ) == ( bv_8_51_n528 )  ;
assign n661 = in[23:16] ;
assign n662 =  ( n661 ) == ( bv_8_50_n349 )  ;
assign bv_8_35_n663 = 8'h23 ;
assign n664 = in[23:16] ;
assign bv_8_49_n665 = 8'h31 ;
assign n666 =  ( n664 ) == ( bv_8_49_n665 )  ;
assign n667 = in[23:16] ;
assign bv_8_48_n668 = 8'h30 ;
assign n669 =  ( n667 ) == ( bv_8_48_n668 )  ;
assign bv_8_4_n670 = 8'h4 ;
assign n671 = in[23:16] ;
assign n672 =  ( n671 ) == ( bv_8_47_n591 )  ;
assign bv_8_21_n673 = 8'h15 ;
assign n674 = in[23:16] ;
assign n675 =  ( n674 ) == ( bv_8_46_n235 )  ;
assign n676 = in[23:16] ;
assign n677 =  ( n676 ) == ( bv_8_45_n26 )  ;
assign n678 = in[23:16] ;
assign n679 =  ( n678 ) == ( bv_8_44_n621 )  ;
assign n680 = in[23:16] ;
assign bv_8_43_n681 = 8'h2b ;
assign n682 =  ( n680 ) == ( bv_8_43_n681 )  ;
assign n683 = in[23:16] ;
assign n684 =  ( n683 ) == ( bv_8_42_n387 )  ;
assign n685 = in[23:16] ;
assign n686 =  ( n685 ) == ( bv_8_41_n596 )  ;
assign n687 = in[23:16] ;
assign n688 =  ( n687 ) == ( bv_8_40_n74 )  ;
assign n689 = in[23:16] ;
assign n690 =  ( n689 ) == ( bv_8_39_n634 )  ;
assign n691 = in[23:16] ;
assign bv_8_38_n692 = 8'h26 ;
assign n693 =  ( n691 ) == ( bv_8_38_n692 )  ;
assign n694 = in[23:16] ;
assign n695 =  ( n694 ) == ( bv_8_37_n239 )  ;
assign n696 = in[23:16] ;
assign n697 =  ( n696 ) == ( bv_8_36_n330 )  ;
assign n698 = in[23:16] ;
assign n699 =  ( n698 ) == ( bv_8_35_n663 )  ;
assign n700 = in[23:16] ;
assign n701 =  ( n700 ) == ( bv_8_34_n390 )  ;
assign n702 = in[23:16] ;
assign n703 =  ( n702 ) == ( bv_8_33_n468 )  ;
assign n704 = in[23:16] ;
assign n705 =  ( n704 ) == ( bv_8_32_n575 )  ;
assign n706 = in[23:16] ;
assign n707 =  ( n706 ) == ( bv_8_31_n206 )  ;
assign n708 = in[23:16] ;
assign n709 =  ( n708 ) == ( bv_8_30_n93 )  ;
assign n710 = in[23:16] ;
assign n711 =  ( n710 ) == ( bv_8_29_n133 )  ;
assign n712 = in[23:16] ;
assign n713 =  ( n712 ) == ( bv_8_28_n231 )  ;
assign n714 = in[23:16] ;
assign n715 =  ( n714 ) == ( bv_8_27_n615 )  ;
assign n716 = in[23:16] ;
assign n717 =  ( n716 ) == ( bv_8_26_n618 )  ;
assign n718 = in[23:16] ;
assign n719 =  ( n718 ) == ( bv_8_25_n410 )  ;
assign n720 = in[23:16] ;
assign n721 =  ( n720 ) == ( bv_8_24_n658 )  ;
assign n722 = in[23:16] ;
assign n723 =  ( n722 ) == ( bv_8_23_n429 )  ;
assign n724 = in[23:16] ;
assign n725 =  ( n724 ) == ( bv_8_22_n6 )  ;
assign n726 = in[23:16] ;
assign n727 =  ( n726 ) == ( bv_8_21_n673 )  ;
assign n728 = in[23:16] ;
assign n729 =  ( n728 ) == ( bv_8_20_n368 )  ;
assign n730 = in[23:16] ;
assign n731 =  ( n730 ) == ( bv_8_19_n446 )  ;
assign n732 = in[23:16] ;
assign n733 =  ( n732 ) == ( bv_8_18_n643 )  ;
assign n734 = in[23:16] ;
assign n735 =  ( n734 ) == ( bv_8_17_n116 )  ;
assign n736 = in[23:16] ;
assign n737 =  ( n736 ) == ( bv_8_16_n464 )  ;
assign n738 = in[23:16] ;
assign n739 =  ( n738 ) == ( bv_8_15_n22 )  ;
assign n740 = in[23:16] ;
assign n741 =  ( n740 ) == ( bv_8_14_n160 )  ;
assign n742 = in[23:16] ;
assign n743 =  ( n742 ) == ( bv_8_13_n54 )  ;
assign n744 = in[23:16] ;
assign n745 =  ( n744 ) == ( bv_8_12_n449 )  ;
assign n746 = in[23:16] ;
assign n747 =  ( n746 ) == ( bv_8_11_n358 )  ;
assign n748 = in[23:16] ;
assign n749 =  ( n748 ) == ( bv_8_10_n342 )  ;
assign n750 = in[23:16] ;
assign n751 =  ( n750 ) == ( bv_8_9_n626 )  ;
assign bv_8_1_n752 = 8'h1 ;
assign n753 = in[23:16] ;
assign n754 =  ( n753 ) == ( bv_8_8_n249 )  ;
assign n755 = in[23:16] ;
assign n756 =  ( n755 ) == ( bv_8_7_n646 )  ;
assign n757 = in[23:16] ;
assign n758 =  ( n757 ) == ( bv_8_6_n334 )  ;
assign n759 = in[23:16] ;
assign n760 =  ( n759 ) == ( bv_8_5_n652 )  ;
assign n761 = in[23:16] ;
assign n762 =  ( n761 ) == ( bv_8_4_n670 )  ;
assign n763 = in[23:16] ;
assign n764 =  ( n763 ) == ( bv_8_3_n167 )  ;
assign n765 = in[23:16] ;
assign n766 =  ( n765 ) == ( bv_8_2_n517 )  ;
assign n767 = in[23:16] ;
assign n768 =  ( n767 ) == ( bv_8_1_n752 )  ;
assign n769 = in[23:16] ;
assign n770 =  ( n769 ) == ( bv_8_0_n582 )  ;
assign n771 =  ( n770 ) ? ( bv_8_99_n536 ) : ( bv_8_0_n582 ) ;
assign n772 =  ( n768 ) ? ( bv_8_124_n462 ) : ( n771 ) ;
assign n773 =  ( n766 ) ? ( bv_8_119_n476 ) : ( n772 ) ;
assign n774 =  ( n764 ) ? ( bv_8_123_n466 ) : ( n773 ) ;
assign n775 =  ( n762 ) ? ( bv_8_242_n56 ) : ( n774 ) ;
assign n776 =  ( n760 ) ? ( bv_8_107_n512 ) : ( n775 ) ;
assign n777 =  ( n758 ) ? ( bv_8_111_n500 ) : ( n776 ) ;
assign n778 =  ( n756 ) ? ( bv_8_197_n225 ) : ( n777 ) ;
assign n779 =  ( n754 ) ? ( bv_8_48_n668 ) : ( n778 ) ;
assign n780 =  ( n751 ) ? ( bv_8_1_n752 ) : ( n779 ) ;
assign n781 =  ( n749 ) ? ( bv_8_103_n524 ) : ( n780 ) ;
assign n782 =  ( n747 ) ? ( bv_8_43_n681 ) : ( n781 ) ;
assign n783 =  ( n745 ) ? ( bv_8_254_n8 ) : ( n782 ) ;
assign n784 =  ( n743 ) ? ( bv_8_215_n158 ) : ( n783 ) ;
assign n785 =  ( n741 ) ? ( bv_8_171_n313 ) : ( n784 ) ;
assign n786 =  ( n739 ) ? ( bv_8_118_n479 ) : ( n785 ) ;
assign n787 =  ( n737 ) ? ( bv_8_202_n208 ) : ( n786 ) ;
assign n788 =  ( n735 ) ? ( bv_8_130_n444 ) : ( n787 ) ;
assign n789 =  ( n733 ) ? ( bv_8_201_n212 ) : ( n788 ) ;
assign n790 =  ( n731 ) ? ( bv_8_125_n459 ) : ( n789 ) ;
assign n791 =  ( n729 ) ? ( bv_8_250_n24 ) : ( n790 ) ;
assign n792 =  ( n727 ) ? ( bv_8_89_n563 ) : ( n791 ) ;
assign n793 =  ( n725 ) ? ( bv_8_71_n607 ) : ( n792 ) ;
assign n794 =  ( n723 ) ? ( bv_8_240_n64 ) : ( n793 ) ;
assign n795 =  ( n721 ) ? ( bv_8_173_n305 ) : ( n794 ) ;
assign n796 =  ( n719 ) ? ( bv_8_212_n169 ) : ( n795 ) ;
assign n797 =  ( n717 ) ? ( bv_8_162_n344 ) : ( n796 ) ;
assign n798 =  ( n715 ) ? ( bv_8_175_n299 ) : ( n797 ) ;
assign n799 =  ( n713 ) ? ( bv_8_156_n364 ) : ( n798 ) ;
assign n800 =  ( n711 ) ? ( bv_8_164_n336 ) : ( n799 ) ;
assign n801 =  ( n709 ) ? ( bv_8_114_n490 ) : ( n800 ) ;
assign n802 =  ( n707 ) ? ( bv_8_192_n244 ) : ( n801 ) ;
assign n803 =  ( n705 ) ? ( bv_8_183_n273 ) : ( n802 ) ;
assign n804 =  ( n703 ) ? ( bv_8_253_n12 ) : ( n803 ) ;
assign n805 =  ( n701 ) ? ( bv_8_147_n392 ) : ( n804 ) ;
assign n806 =  ( n699 ) ? ( bv_8_38_n692 ) : ( n805 ) ;
assign n807 =  ( n697 ) ? ( bv_8_54_n650 ) : ( n806 ) ;
assign n808 =  ( n695 ) ? ( bv_8_63_n628 ) : ( n807 ) ;
assign n809 =  ( n693 ) ? ( bv_8_247_n36 ) : ( n808 ) ;
assign n810 =  ( n690 ) ? ( bv_8_204_n200 ) : ( n809 ) ;
assign n811 =  ( n688 ) ? ( bv_8_52_n656 ) : ( n810 ) ;
assign n812 =  ( n686 ) ? ( bv_8_165_n332 ) : ( n811 ) ;
assign n813 =  ( n684 ) ? ( bv_8_229_n106 ) : ( n812 ) ;
assign n814 =  ( n682 ) ? ( bv_8_241_n60 ) : ( n813 ) ;
assign n815 =  ( n679 ) ? ( bv_8_113_n494 ) : ( n814 ) ;
assign n816 =  ( n677 ) ? ( bv_8_216_n154 ) : ( n815 ) ;
assign n817 =  ( n675 ) ? ( bv_8_49_n665 ) : ( n816 ) ;
assign n818 =  ( n672 ) ? ( bv_8_21_n673 ) : ( n817 ) ;
assign n819 =  ( n669 ) ? ( bv_8_4_n670 ) : ( n818 ) ;
assign n820 =  ( n666 ) ? ( bv_8_199_n218 ) : ( n819 ) ;
assign n821 =  ( n662 ) ? ( bv_8_35_n663 ) : ( n820 ) ;
assign n822 =  ( n660 ) ? ( bv_8_195_n233 ) : ( n821 ) ;
assign n823 =  ( n657 ) ? ( bv_8_24_n658 ) : ( n822 ) ;
assign n824 =  ( n654 ) ? ( bv_8_150_n382 ) : ( n823 ) ;
assign n825 =  ( n651 ) ? ( bv_8_5_n652 ) : ( n824 ) ;
assign n826 =  ( n648 ) ? ( bv_8_154_n370 ) : ( n825 ) ;
assign n827 =  ( n645 ) ? ( bv_8_7_n646 ) : ( n826 ) ;
assign n828 =  ( n642 ) ? ( bv_8_18_n643 ) : ( n827 ) ;
assign n829 =  ( n640 ) ? ( bv_8_128_n451 ) : ( n828 ) ;
assign n830 =  ( n638 ) ? ( bv_8_226_n118 ) : ( n829 ) ;
assign n831 =  ( n636 ) ? ( bv_8_235_n84 ) : ( n830 ) ;
assign n832 =  ( n633 ) ? ( bv_8_39_n634 ) : ( n831 ) ;
assign n833 =  ( n631 ) ? ( bv_8_178_n290 ) : ( n832 ) ;
assign n834 =  ( n629 ) ? ( bv_8_117_n483 ) : ( n833 ) ;
assign n835 =  ( n625 ) ? ( bv_8_9_n626 ) : ( n834 ) ;
assign n836 =  ( n623 ) ? ( bv_8_131_n441 ) : ( n835 ) ;
assign n837 =  ( n620 ) ? ( bv_8_44_n621 ) : ( n836 ) ;
assign n838 =  ( n617 ) ? ( bv_8_26_n618 ) : ( n837 ) ;
assign n839 =  ( n614 ) ? ( bv_8_27_n615 ) : ( n838 ) ;
assign n840 =  ( n612 ) ? ( bv_8_110_n503 ) : ( n839 ) ;
assign n841 =  ( n610 ) ? ( bv_8_90_n560 ) : ( n840 ) ;
assign n842 =  ( n608 ) ? ( bv_8_160_n351 ) : ( n841 ) ;
assign n843 =  ( n605 ) ? ( bv_8_82_n580 ) : ( n842 ) ;
assign n844 =  ( n602 ) ? ( bv_8_59_n603 ) : ( n843 ) ;
assign n845 =  ( n600 ) ? ( bv_8_214_n162 ) : ( n844 ) ;
assign n846 =  ( n598 ) ? ( bv_8_179_n286 ) : ( n845 ) ;
assign n847 =  ( n595 ) ? ( bv_8_41_n596 ) : ( n846 ) ;
assign n848 =  ( n593 ) ? ( bv_8_227_n114 ) : ( n847 ) ;
assign n849 =  ( n590 ) ? ( bv_8_47_n591 ) : ( n848 ) ;
assign n850 =  ( n588 ) ? ( bv_8_132_n437 ) : ( n849 ) ;
assign n851 =  ( n586 ) ? ( bv_8_83_n577 ) : ( n850 ) ;
assign n852 =  ( n584 ) ? ( bv_8_209_n181 ) : ( n851 ) ;
assign n853 =  ( n581 ) ? ( bv_8_0_n582 ) : ( n852 ) ;
assign n854 =  ( n578 ) ? ( bv_8_237_n76 ) : ( n853 ) ;
assign n855 =  ( n574 ) ? ( bv_8_32_n575 ) : ( n854 ) ;
assign n856 =  ( n572 ) ? ( bv_8_252_n16 ) : ( n855 ) ;
assign n857 =  ( n570 ) ? ( bv_8_177_n294 ) : ( n856 ) ;
assign n858 =  ( n568 ) ? ( bv_8_91_n556 ) : ( n857 ) ;
assign n859 =  ( n566 ) ? ( bv_8_106_n515 ) : ( n858 ) ;
assign n860 =  ( n564 ) ? ( bv_8_203_n204 ) : ( n859 ) ;
assign n861 =  ( n561 ) ? ( bv_8_190_n251 ) : ( n860 ) ;
assign n862 =  ( n557 ) ? ( bv_8_57_n558 ) : ( n861 ) ;
assign n863 =  ( n553 ) ? ( bv_8_74_n554 ) : ( n862 ) ;
assign n864 =  ( n550 ) ? ( bv_8_76_n551 ) : ( n863 ) ;
assign n865 =  ( n547 ) ? ( bv_8_88_n548 ) : ( n864 ) ;
assign n866 =  ( n545 ) ? ( bv_8_207_n189 ) : ( n865 ) ;
assign n867 =  ( n543 ) ? ( bv_8_208_n185 ) : ( n866 ) ;
assign n868 =  ( n541 ) ? ( bv_8_239_n68 ) : ( n867 ) ;
assign n869 =  ( n539 ) ? ( bv_8_170_n317 ) : ( n868 ) ;
assign n870 =  ( n537 ) ? ( bv_8_251_n20 ) : ( n869 ) ;
assign n871 =  ( n533 ) ? ( bv_8_67_n534 ) : ( n870 ) ;
assign n872 =  ( n530 ) ? ( bv_8_77_n531 ) : ( n871 ) ;
assign n873 =  ( n527 ) ? ( bv_8_51_n528 ) : ( n872 ) ;
assign n874 =  ( n525 ) ? ( bv_8_133_n434 ) : ( n873 ) ;
assign n875 =  ( n521 ) ? ( bv_8_69_n522 ) : ( n874 ) ;
assign n876 =  ( n519 ) ? ( bv_8_249_n28 ) : ( n875 ) ;
assign n877 =  ( n516 ) ? ( bv_8_2_n517 ) : ( n876 ) ;
assign n878 =  ( n513 ) ? ( bv_8_127_n454 ) : ( n877 ) ;
assign n879 =  ( n509 ) ? ( bv_8_80_n510 ) : ( n878 ) ;
assign n880 =  ( n506 ) ? ( bv_8_60_n507 ) : ( n879 ) ;
assign n881 =  ( n504 ) ? ( bv_8_159_n354 ) : ( n880 ) ;
assign n882 =  ( n501 ) ? ( bv_8_168_n322 ) : ( n881 ) ;
assign n883 =  ( n497 ) ? ( bv_8_81_n498 ) : ( n882 ) ;
assign n884 =  ( n495 ) ? ( bv_8_163_n340 ) : ( n883 ) ;
assign n885 =  ( n491 ) ? ( bv_8_64_n492 ) : ( n884 ) ;
assign n886 =  ( n488 ) ? ( bv_8_143_n405 ) : ( n885 ) ;
assign n887 =  ( n486 ) ? ( bv_8_146_n395 ) : ( n886 ) ;
assign n888 =  ( n484 ) ? ( bv_8_157_n360 ) : ( n887 ) ;
assign n889 =  ( n480 ) ? ( bv_8_56_n481 ) : ( n888 ) ;
assign n890 =  ( n477 ) ? ( bv_8_245_n44 ) : ( n889 ) ;
assign n891 =  ( n474 ) ? ( bv_8_188_n258 ) : ( n890 ) ;
assign n892 =  ( n472 ) ? ( bv_8_182_n277 ) : ( n891 ) ;
assign n893 =  ( n470 ) ? ( bv_8_218_n147 ) : ( n892 ) ;
assign n894 =  ( n467 ) ? ( bv_8_33_n468 ) : ( n893 ) ;
assign n895 =  ( n463 ) ? ( bv_8_16_n464 ) : ( n894 ) ;
assign n896 =  ( n460 ) ? ( bv_8_255_n4 ) : ( n895 ) ;
assign n897 =  ( n457 ) ? ( bv_8_243_n52 ) : ( n896 ) ;
assign n898 =  ( n455 ) ? ( bv_8_210_n177 ) : ( n897 ) ;
assign n899 =  ( n452 ) ? ( bv_8_205_n196 ) : ( n898 ) ;
assign n900 =  ( n448 ) ? ( bv_8_12_n449 ) : ( n899 ) ;
assign n901 =  ( n445 ) ? ( bv_8_19_n446 ) : ( n900 ) ;
assign n902 =  ( n442 ) ? ( bv_8_236_n80 ) : ( n901 ) ;
assign n903 =  ( n438 ) ? ( bv_8_95_n439 ) : ( n902 ) ;
assign n904 =  ( n435 ) ? ( bv_8_151_n378 ) : ( n903 ) ;
assign n905 =  ( n431 ) ? ( bv_8_68_n432 ) : ( n904 ) ;
assign n906 =  ( n428 ) ? ( bv_8_23_n429 ) : ( n905 ) ;
assign n907 =  ( n426 ) ? ( bv_8_196_n229 ) : ( n906 ) ;
assign n908 =  ( n424 ) ? ( bv_8_167_n325 ) : ( n907 ) ;
assign n909 =  ( n421 ) ? ( bv_8_126_n422 ) : ( n908 ) ;
assign n910 =  ( n418 ) ? ( bv_8_61_n419 ) : ( n909 ) ;
assign n911 =  ( n415 ) ? ( bv_8_100_n416 ) : ( n910 ) ;
assign n912 =  ( n412 ) ? ( bv_8_93_n413 ) : ( n911 ) ;
assign n913 =  ( n409 ) ? ( bv_8_25_n410 ) : ( n912 ) ;
assign n914 =  ( n406 ) ? ( bv_8_115_n407 ) : ( n913 ) ;
assign n915 =  ( n402 ) ? ( bv_8_96_n403 ) : ( n914 ) ;
assign n916 =  ( n399 ) ? ( bv_8_129_n400 ) : ( n915 ) ;
assign n917 =  ( n396 ) ? ( bv_8_79_n397 ) : ( n916 ) ;
assign n918 =  ( n393 ) ? ( bv_8_220_n139 ) : ( n917 ) ;
assign n919 =  ( n389 ) ? ( bv_8_34_n390 ) : ( n918 ) ;
assign n920 =  ( n386 ) ? ( bv_8_42_n387 ) : ( n919 ) ;
assign n921 =  ( n383 ) ? ( bv_8_144_n384 ) : ( n920 ) ;
assign n922 =  ( n379 ) ? ( bv_8_136_n380 ) : ( n921 ) ;
assign n923 =  ( n375 ) ? ( bv_8_70_n376 ) : ( n922 ) ;
assign n924 =  ( n373 ) ? ( bv_8_238_n72 ) : ( n923 ) ;
assign n925 =  ( n371 ) ? ( bv_8_184_n269 ) : ( n924 ) ;
assign n926 =  ( n367 ) ? ( bv_8_20_n368 ) : ( n925 ) ;
assign n927 =  ( n365 ) ? ( bv_8_222_n131 ) : ( n926 ) ;
assign n928 =  ( n361 ) ? ( bv_8_94_n362 ) : ( n927 ) ;
assign n929 =  ( n357 ) ? ( bv_8_11_n358 ) : ( n928 ) ;
assign n930 =  ( n355 ) ? ( bv_8_219_n143 ) : ( n929 ) ;
assign n931 =  ( n352 ) ? ( bv_8_224_n125 ) : ( n930 ) ;
assign n932 =  ( n348 ) ? ( bv_8_50_n349 ) : ( n931 ) ;
assign n933 =  ( n345 ) ? ( bv_8_58_n346 ) : ( n932 ) ;
assign n934 =  ( n341 ) ? ( bv_8_10_n342 ) : ( n933 ) ;
assign n935 =  ( n337 ) ? ( bv_8_73_n338 ) : ( n934 ) ;
assign n936 =  ( n333 ) ? ( bv_8_6_n334 ) : ( n935 ) ;
assign n937 =  ( n329 ) ? ( bv_8_36_n330 ) : ( n936 ) ;
assign n938 =  ( n326 ) ? ( bv_8_92_n327 ) : ( n937 ) ;
assign n939 =  ( n323 ) ? ( bv_8_194_n237 ) : ( n938 ) ;
assign n940 =  ( n320 ) ? ( bv_8_211_n173 ) : ( n939 ) ;
assign n941 =  ( n318 ) ? ( bv_8_172_n309 ) : ( n940 ) ;
assign n942 =  ( n314 ) ? ( bv_8_98_n315 ) : ( n941 ) ;
assign n943 =  ( n310 ) ? ( bv_8_145_n311 ) : ( n942 ) ;
assign n944 =  ( n306 ) ? ( bv_8_149_n307 ) : ( n943 ) ;
assign n945 =  ( n303 ) ? ( bv_8_228_n110 ) : ( n944 ) ;
assign n946 =  ( n300 ) ? ( bv_8_121_n301 ) : ( n945 ) ;
assign n947 =  ( n297 ) ? ( bv_8_231_n99 ) : ( n946 ) ;
assign n948 =  ( n295 ) ? ( bv_8_200_n215 ) : ( n947 ) ;
assign n949 =  ( n291 ) ? ( bv_8_55_n292 ) : ( n948 ) ;
assign n950 =  ( n287 ) ? ( bv_8_109_n288 ) : ( n949 ) ;
assign n951 =  ( n283 ) ? ( bv_8_141_n284 ) : ( n950 ) ;
assign n952 =  ( n281 ) ? ( bv_8_213_n165 ) : ( n951 ) ;
assign n953 =  ( n278 ) ? ( bv_8_78_n279 ) : ( n952 ) ;
assign n954 =  ( n274 ) ? ( bv_8_169_n275 ) : ( n953 ) ;
assign n955 =  ( n270 ) ? ( bv_8_108_n271 ) : ( n954 ) ;
assign n956 =  ( n266 ) ? ( bv_8_86_n267 ) : ( n955 ) ;
assign n957 =  ( n264 ) ? ( bv_8_244_n48 ) : ( n956 ) ;
assign n958 =  ( n262 ) ? ( bv_8_234_n88 ) : ( n957 ) ;
assign n959 =  ( n259 ) ? ( bv_8_101_n260 ) : ( n958 ) ;
assign n960 =  ( n255 ) ? ( bv_8_122_n256 ) : ( n959 ) ;
assign n961 =  ( n252 ) ? ( bv_8_174_n253 ) : ( n960 ) ;
assign n962 =  ( n248 ) ? ( bv_8_8_n249 ) : ( n961 ) ;
assign n963 =  ( n245 ) ? ( bv_8_186_n246 ) : ( n962 ) ;
assign n964 =  ( n241 ) ? ( bv_8_120_n242 ) : ( n963 ) ;
assign n965 =  ( n238 ) ? ( bv_8_37_n239 ) : ( n964 ) ;
assign n966 =  ( n234 ) ? ( bv_8_46_n235 ) : ( n965 ) ;
assign n967 =  ( n230 ) ? ( bv_8_28_n231 ) : ( n966 ) ;
assign n968 =  ( n226 ) ? ( bv_8_166_n227 ) : ( n967 ) ;
assign n969 =  ( n222 ) ? ( bv_8_180_n223 ) : ( n968 ) ;
assign n970 =  ( n219 ) ? ( bv_8_198_n220 ) : ( n969 ) ;
assign n971 =  ( n216 ) ? ( bv_8_232_n95 ) : ( n970 ) ;
assign n972 =  ( n213 ) ? ( bv_8_221_n135 ) : ( n971 ) ;
assign n973 =  ( n209 ) ? ( bv_8_116_n210 ) : ( n972 ) ;
assign n974 =  ( n205 ) ? ( bv_8_31_n206 ) : ( n973 ) ;
assign n975 =  ( n201 ) ? ( bv_8_75_n202 ) : ( n974 ) ;
assign n976 =  ( n197 ) ? ( bv_8_189_n198 ) : ( n975 ) ;
assign n977 =  ( n193 ) ? ( bv_8_139_n194 ) : ( n976 ) ;
assign n978 =  ( n190 ) ? ( bv_8_138_n191 ) : ( n977 ) ;
assign n979 =  ( n186 ) ? ( bv_8_112_n187 ) : ( n978 ) ;
assign n980 =  ( n182 ) ? ( bv_8_62_n183 ) : ( n979 ) ;
assign n981 =  ( n178 ) ? ( bv_8_181_n179 ) : ( n980 ) ;
assign n982 =  ( n174 ) ? ( bv_8_102_n175 ) : ( n981 ) ;
assign n983 =  ( n170 ) ? ( bv_8_72_n171 ) : ( n982 ) ;
assign n984 =  ( n166 ) ? ( bv_8_3_n167 ) : ( n983 ) ;
assign n985 =  ( n163 ) ? ( bv_8_246_n40 ) : ( n984 ) ;
assign n986 =  ( n159 ) ? ( bv_8_14_n160 ) : ( n985 ) ;
assign n987 =  ( n155 ) ? ( bv_8_97_n156 ) : ( n986 ) ;
assign n988 =  ( n151 ) ? ( bv_8_53_n152 ) : ( n987 ) ;
assign n989 =  ( n148 ) ? ( bv_8_87_n149 ) : ( n988 ) ;
assign n990 =  ( n144 ) ? ( bv_8_185_n145 ) : ( n989 ) ;
assign n991 =  ( n140 ) ? ( bv_8_134_n141 ) : ( n990 ) ;
assign n992 =  ( n136 ) ? ( bv_8_193_n137 ) : ( n991 ) ;
assign n993 =  ( n132 ) ? ( bv_8_29_n133 ) : ( n992 ) ;
assign n994 =  ( n128 ) ? ( bv_8_158_n129 ) : ( n993 ) ;
assign n995 =  ( n126 ) ? ( bv_8_225_n122 ) : ( n994 ) ;
assign n996 =  ( n123 ) ? ( bv_8_248_n32 ) : ( n995 ) ;
assign n997 =  ( n119 ) ? ( bv_8_152_n120 ) : ( n996 ) ;
assign n998 =  ( n115 ) ? ( bv_8_17_n116 ) : ( n997 ) ;
assign n999 =  ( n111 ) ? ( bv_8_105_n112 ) : ( n998 ) ;
assign n1000 =  ( n107 ) ? ( bv_8_217_n108 ) : ( n999 ) ;
assign n1001 =  ( n103 ) ? ( bv_8_142_n104 ) : ( n1000 ) ;
assign n1002 =  ( n100 ) ? ( bv_8_148_n101 ) : ( n1001 ) ;
assign n1003 =  ( n96 ) ? ( bv_8_155_n97 ) : ( n1002 ) ;
assign n1004 =  ( n92 ) ? ( bv_8_30_n93 ) : ( n1003 ) ;
assign n1005 =  ( n89 ) ? ( bv_8_135_n90 ) : ( n1004 ) ;
assign n1006 =  ( n85 ) ? ( bv_8_233_n86 ) : ( n1005 ) ;
assign n1007 =  ( n81 ) ? ( bv_8_206_n82 ) : ( n1006 ) ;
assign n1008 =  ( n77 ) ? ( bv_8_85_n78 ) : ( n1007 ) ;
assign n1009 =  ( n73 ) ? ( bv_8_40_n74 ) : ( n1008 ) ;
assign n1010 =  ( n69 ) ? ( bv_8_223_n70 ) : ( n1009 ) ;
assign n1011 =  ( n65 ) ? ( bv_8_140_n66 ) : ( n1010 ) ;
assign n1012 =  ( n61 ) ? ( bv_8_161_n62 ) : ( n1011 ) ;
assign n1013 =  ( n57 ) ? ( bv_8_137_n58 ) : ( n1012 ) ;
assign n1014 =  ( n53 ) ? ( bv_8_13_n54 ) : ( n1013 ) ;
assign n1015 =  ( n49 ) ? ( bv_8_191_n50 ) : ( n1014 ) ;
assign n1016 =  ( n45 ) ? ( bv_8_230_n46 ) : ( n1015 ) ;
assign n1017 =  ( n41 ) ? ( bv_8_66_n42 ) : ( n1016 ) ;
assign n1018 =  ( n37 ) ? ( bv_8_104_n38 ) : ( n1017 ) ;
assign n1019 =  ( n33 ) ? ( bv_8_65_n34 ) : ( n1018 ) ;
assign n1020 =  ( n29 ) ? ( bv_8_153_n30 ) : ( n1019 ) ;
assign n1021 =  ( n25 ) ? ( bv_8_45_n26 ) : ( n1020 ) ;
assign n1022 =  ( n21 ) ? ( bv_8_15_n22 ) : ( n1021 ) ;
assign n1023 =  ( n17 ) ? ( bv_8_176_n18 ) : ( n1022 ) ;
assign n1024 =  ( n13 ) ? ( bv_8_84_n14 ) : ( n1023 ) ;
assign n1025 =  ( n9 ) ? ( bv_8_187_n10 ) : ( n1024 ) ;
assign n1026 =  ( n5 ) ? ( bv_8_22_n6 ) : ( n1025 ) ;
assign n1027 =  ( n2 ) ^ ( n1026 )  ;
assign n1028 = in[119:112] ;
assign n1029 = in[15:8] ;
assign n1030 =  ( n1029 ) == ( bv_8_255_n4 )  ;
assign n1031 = in[15:8] ;
assign n1032 =  ( n1031 ) == ( bv_8_254_n8 )  ;
assign n1033 = in[15:8] ;
assign n1034 =  ( n1033 ) == ( bv_8_253_n12 )  ;
assign n1035 = in[15:8] ;
assign n1036 =  ( n1035 ) == ( bv_8_252_n16 )  ;
assign n1037 = in[15:8] ;
assign n1038 =  ( n1037 ) == ( bv_8_251_n20 )  ;
assign n1039 = in[15:8] ;
assign n1040 =  ( n1039 ) == ( bv_8_250_n24 )  ;
assign n1041 = in[15:8] ;
assign n1042 =  ( n1041 ) == ( bv_8_249_n28 )  ;
assign n1043 = in[15:8] ;
assign n1044 =  ( n1043 ) == ( bv_8_248_n32 )  ;
assign n1045 = in[15:8] ;
assign n1046 =  ( n1045 ) == ( bv_8_247_n36 )  ;
assign n1047 = in[15:8] ;
assign n1048 =  ( n1047 ) == ( bv_8_246_n40 )  ;
assign n1049 = in[15:8] ;
assign n1050 =  ( n1049 ) == ( bv_8_245_n44 )  ;
assign n1051 = in[15:8] ;
assign n1052 =  ( n1051 ) == ( bv_8_244_n48 )  ;
assign n1053 = in[15:8] ;
assign n1054 =  ( n1053 ) == ( bv_8_243_n52 )  ;
assign n1055 = in[15:8] ;
assign n1056 =  ( n1055 ) == ( bv_8_242_n56 )  ;
assign n1057 = in[15:8] ;
assign n1058 =  ( n1057 ) == ( bv_8_241_n60 )  ;
assign n1059 = in[15:8] ;
assign n1060 =  ( n1059 ) == ( bv_8_240_n64 )  ;
assign n1061 = in[15:8] ;
assign n1062 =  ( n1061 ) == ( bv_8_239_n68 )  ;
assign n1063 = in[15:8] ;
assign n1064 =  ( n1063 ) == ( bv_8_238_n72 )  ;
assign n1065 = in[15:8] ;
assign n1066 =  ( n1065 ) == ( bv_8_237_n76 )  ;
assign n1067 = in[15:8] ;
assign n1068 =  ( n1067 ) == ( bv_8_236_n80 )  ;
assign n1069 = in[15:8] ;
assign n1070 =  ( n1069 ) == ( bv_8_235_n84 )  ;
assign n1071 = in[15:8] ;
assign n1072 =  ( n1071 ) == ( bv_8_234_n88 )  ;
assign n1073 = in[15:8] ;
assign n1074 =  ( n1073 ) == ( bv_8_233_n86 )  ;
assign n1075 = in[15:8] ;
assign n1076 =  ( n1075 ) == ( bv_8_232_n95 )  ;
assign n1077 = in[15:8] ;
assign n1078 =  ( n1077 ) == ( bv_8_231_n99 )  ;
assign n1079 = in[15:8] ;
assign n1080 =  ( n1079 ) == ( bv_8_230_n46 )  ;
assign n1081 = in[15:8] ;
assign n1082 =  ( n1081 ) == ( bv_8_229_n106 )  ;
assign n1083 = in[15:8] ;
assign n1084 =  ( n1083 ) == ( bv_8_228_n110 )  ;
assign n1085 = in[15:8] ;
assign n1086 =  ( n1085 ) == ( bv_8_227_n114 )  ;
assign n1087 = in[15:8] ;
assign n1088 =  ( n1087 ) == ( bv_8_226_n118 )  ;
assign n1089 = in[15:8] ;
assign n1090 =  ( n1089 ) == ( bv_8_225_n122 )  ;
assign n1091 = in[15:8] ;
assign n1092 =  ( n1091 ) == ( bv_8_224_n125 )  ;
assign n1093 = in[15:8] ;
assign n1094 =  ( n1093 ) == ( bv_8_223_n70 )  ;
assign n1095 = in[15:8] ;
assign n1096 =  ( n1095 ) == ( bv_8_222_n131 )  ;
assign n1097 = in[15:8] ;
assign n1098 =  ( n1097 ) == ( bv_8_221_n135 )  ;
assign n1099 = in[15:8] ;
assign n1100 =  ( n1099 ) == ( bv_8_220_n139 )  ;
assign n1101 = in[15:8] ;
assign n1102 =  ( n1101 ) == ( bv_8_219_n143 )  ;
assign n1103 = in[15:8] ;
assign n1104 =  ( n1103 ) == ( bv_8_218_n147 )  ;
assign n1105 = in[15:8] ;
assign n1106 =  ( n1105 ) == ( bv_8_217_n108 )  ;
assign n1107 = in[15:8] ;
assign n1108 =  ( n1107 ) == ( bv_8_216_n154 )  ;
assign n1109 = in[15:8] ;
assign n1110 =  ( n1109 ) == ( bv_8_215_n158 )  ;
assign n1111 = in[15:8] ;
assign n1112 =  ( n1111 ) == ( bv_8_214_n162 )  ;
assign n1113 = in[15:8] ;
assign n1114 =  ( n1113 ) == ( bv_8_213_n165 )  ;
assign n1115 = in[15:8] ;
assign n1116 =  ( n1115 ) == ( bv_8_212_n169 )  ;
assign n1117 = in[15:8] ;
assign n1118 =  ( n1117 ) == ( bv_8_211_n173 )  ;
assign n1119 = in[15:8] ;
assign n1120 =  ( n1119 ) == ( bv_8_210_n177 )  ;
assign n1121 = in[15:8] ;
assign n1122 =  ( n1121 ) == ( bv_8_209_n181 )  ;
assign n1123 = in[15:8] ;
assign n1124 =  ( n1123 ) == ( bv_8_208_n185 )  ;
assign n1125 = in[15:8] ;
assign n1126 =  ( n1125 ) == ( bv_8_207_n189 )  ;
assign n1127 = in[15:8] ;
assign n1128 =  ( n1127 ) == ( bv_8_206_n82 )  ;
assign n1129 = in[15:8] ;
assign n1130 =  ( n1129 ) == ( bv_8_205_n196 )  ;
assign n1131 = in[15:8] ;
assign n1132 =  ( n1131 ) == ( bv_8_204_n200 )  ;
assign n1133 = in[15:8] ;
assign n1134 =  ( n1133 ) == ( bv_8_203_n204 )  ;
assign n1135 = in[15:8] ;
assign n1136 =  ( n1135 ) == ( bv_8_202_n208 )  ;
assign n1137 = in[15:8] ;
assign n1138 =  ( n1137 ) == ( bv_8_201_n212 )  ;
assign n1139 = in[15:8] ;
assign n1140 =  ( n1139 ) == ( bv_8_200_n215 )  ;
assign n1141 = in[15:8] ;
assign n1142 =  ( n1141 ) == ( bv_8_199_n218 )  ;
assign n1143 = in[15:8] ;
assign n1144 =  ( n1143 ) == ( bv_8_198_n220 )  ;
assign n1145 = in[15:8] ;
assign n1146 =  ( n1145 ) == ( bv_8_197_n225 )  ;
assign n1147 = in[15:8] ;
assign n1148 =  ( n1147 ) == ( bv_8_196_n229 )  ;
assign n1149 = in[15:8] ;
assign n1150 =  ( n1149 ) == ( bv_8_195_n233 )  ;
assign n1151 = in[15:8] ;
assign n1152 =  ( n1151 ) == ( bv_8_194_n237 )  ;
assign n1153 = in[15:8] ;
assign n1154 =  ( n1153 ) == ( bv_8_193_n137 )  ;
assign n1155 = in[15:8] ;
assign n1156 =  ( n1155 ) == ( bv_8_192_n244 )  ;
assign n1157 = in[15:8] ;
assign n1158 =  ( n1157 ) == ( bv_8_191_n50 )  ;
assign n1159 = in[15:8] ;
assign n1160 =  ( n1159 ) == ( bv_8_190_n251 )  ;
assign n1161 = in[15:8] ;
assign n1162 =  ( n1161 ) == ( bv_8_189_n198 )  ;
assign n1163 = in[15:8] ;
assign n1164 =  ( n1163 ) == ( bv_8_188_n258 )  ;
assign n1165 = in[15:8] ;
assign n1166 =  ( n1165 ) == ( bv_8_187_n10 )  ;
assign n1167 = in[15:8] ;
assign n1168 =  ( n1167 ) == ( bv_8_186_n246 )  ;
assign n1169 = in[15:8] ;
assign n1170 =  ( n1169 ) == ( bv_8_185_n145 )  ;
assign n1171 = in[15:8] ;
assign n1172 =  ( n1171 ) == ( bv_8_184_n269 )  ;
assign n1173 = in[15:8] ;
assign n1174 =  ( n1173 ) == ( bv_8_183_n273 )  ;
assign n1175 = in[15:8] ;
assign n1176 =  ( n1175 ) == ( bv_8_182_n277 )  ;
assign n1177 = in[15:8] ;
assign n1178 =  ( n1177 ) == ( bv_8_181_n179 )  ;
assign n1179 = in[15:8] ;
assign n1180 =  ( n1179 ) == ( bv_8_180_n223 )  ;
assign n1181 = in[15:8] ;
assign n1182 =  ( n1181 ) == ( bv_8_179_n286 )  ;
assign n1183 = in[15:8] ;
assign n1184 =  ( n1183 ) == ( bv_8_178_n290 )  ;
assign n1185 = in[15:8] ;
assign n1186 =  ( n1185 ) == ( bv_8_177_n294 )  ;
assign n1187 = in[15:8] ;
assign n1188 =  ( n1187 ) == ( bv_8_176_n18 )  ;
assign n1189 = in[15:8] ;
assign n1190 =  ( n1189 ) == ( bv_8_175_n299 )  ;
assign n1191 = in[15:8] ;
assign n1192 =  ( n1191 ) == ( bv_8_174_n253 )  ;
assign n1193 = in[15:8] ;
assign n1194 =  ( n1193 ) == ( bv_8_173_n305 )  ;
assign n1195 = in[15:8] ;
assign n1196 =  ( n1195 ) == ( bv_8_172_n309 )  ;
assign n1197 = in[15:8] ;
assign n1198 =  ( n1197 ) == ( bv_8_171_n313 )  ;
assign n1199 = in[15:8] ;
assign n1200 =  ( n1199 ) == ( bv_8_170_n317 )  ;
assign n1201 = in[15:8] ;
assign n1202 =  ( n1201 ) == ( bv_8_169_n275 )  ;
assign n1203 = in[15:8] ;
assign n1204 =  ( n1203 ) == ( bv_8_168_n322 )  ;
assign n1205 = in[15:8] ;
assign n1206 =  ( n1205 ) == ( bv_8_167_n325 )  ;
assign n1207 = in[15:8] ;
assign n1208 =  ( n1207 ) == ( bv_8_166_n227 )  ;
assign n1209 = in[15:8] ;
assign n1210 =  ( n1209 ) == ( bv_8_165_n332 )  ;
assign n1211 = in[15:8] ;
assign n1212 =  ( n1211 ) == ( bv_8_164_n336 )  ;
assign n1213 = in[15:8] ;
assign n1214 =  ( n1213 ) == ( bv_8_163_n340 )  ;
assign n1215 = in[15:8] ;
assign n1216 =  ( n1215 ) == ( bv_8_162_n344 )  ;
assign n1217 = in[15:8] ;
assign n1218 =  ( n1217 ) == ( bv_8_161_n62 )  ;
assign n1219 = in[15:8] ;
assign n1220 =  ( n1219 ) == ( bv_8_160_n351 )  ;
assign n1221 = in[15:8] ;
assign n1222 =  ( n1221 ) == ( bv_8_159_n354 )  ;
assign n1223 = in[15:8] ;
assign n1224 =  ( n1223 ) == ( bv_8_158_n129 )  ;
assign n1225 = in[15:8] ;
assign n1226 =  ( n1225 ) == ( bv_8_157_n360 )  ;
assign n1227 = in[15:8] ;
assign n1228 =  ( n1227 ) == ( bv_8_156_n364 )  ;
assign n1229 = in[15:8] ;
assign n1230 =  ( n1229 ) == ( bv_8_155_n97 )  ;
assign n1231 = in[15:8] ;
assign n1232 =  ( n1231 ) == ( bv_8_154_n370 )  ;
assign n1233 = in[15:8] ;
assign n1234 =  ( n1233 ) == ( bv_8_153_n30 )  ;
assign n1235 = in[15:8] ;
assign n1236 =  ( n1235 ) == ( bv_8_152_n120 )  ;
assign n1237 = in[15:8] ;
assign n1238 =  ( n1237 ) == ( bv_8_151_n378 )  ;
assign n1239 = in[15:8] ;
assign n1240 =  ( n1239 ) == ( bv_8_150_n382 )  ;
assign n1241 = in[15:8] ;
assign n1242 =  ( n1241 ) == ( bv_8_149_n307 )  ;
assign n1243 = in[15:8] ;
assign n1244 =  ( n1243 ) == ( bv_8_148_n101 )  ;
assign n1245 = in[15:8] ;
assign n1246 =  ( n1245 ) == ( bv_8_147_n392 )  ;
assign n1247 = in[15:8] ;
assign n1248 =  ( n1247 ) == ( bv_8_146_n395 )  ;
assign n1249 = in[15:8] ;
assign n1250 =  ( n1249 ) == ( bv_8_145_n311 )  ;
assign n1251 = in[15:8] ;
assign n1252 =  ( n1251 ) == ( bv_8_144_n384 )  ;
assign n1253 = in[15:8] ;
assign n1254 =  ( n1253 ) == ( bv_8_143_n405 )  ;
assign n1255 = in[15:8] ;
assign n1256 =  ( n1255 ) == ( bv_8_142_n104 )  ;
assign n1257 = in[15:8] ;
assign n1258 =  ( n1257 ) == ( bv_8_141_n284 )  ;
assign n1259 = in[15:8] ;
assign n1260 =  ( n1259 ) == ( bv_8_140_n66 )  ;
assign n1261 = in[15:8] ;
assign n1262 =  ( n1261 ) == ( bv_8_139_n194 )  ;
assign n1263 = in[15:8] ;
assign n1264 =  ( n1263 ) == ( bv_8_138_n191 )  ;
assign n1265 = in[15:8] ;
assign n1266 =  ( n1265 ) == ( bv_8_137_n58 )  ;
assign n1267 = in[15:8] ;
assign n1268 =  ( n1267 ) == ( bv_8_136_n380 )  ;
assign n1269 = in[15:8] ;
assign n1270 =  ( n1269 ) == ( bv_8_135_n90 )  ;
assign n1271 = in[15:8] ;
assign n1272 =  ( n1271 ) == ( bv_8_134_n141 )  ;
assign n1273 = in[15:8] ;
assign n1274 =  ( n1273 ) == ( bv_8_133_n434 )  ;
assign n1275 = in[15:8] ;
assign n1276 =  ( n1275 ) == ( bv_8_132_n437 )  ;
assign n1277 = in[15:8] ;
assign n1278 =  ( n1277 ) == ( bv_8_131_n441 )  ;
assign n1279 = in[15:8] ;
assign n1280 =  ( n1279 ) == ( bv_8_130_n444 )  ;
assign n1281 = in[15:8] ;
assign n1282 =  ( n1281 ) == ( bv_8_129_n400 )  ;
assign n1283 = in[15:8] ;
assign n1284 =  ( n1283 ) == ( bv_8_128_n451 )  ;
assign n1285 = in[15:8] ;
assign n1286 =  ( n1285 ) == ( bv_8_127_n454 )  ;
assign n1287 = in[15:8] ;
assign n1288 =  ( n1287 ) == ( bv_8_126_n422 )  ;
assign n1289 = in[15:8] ;
assign n1290 =  ( n1289 ) == ( bv_8_125_n459 )  ;
assign n1291 = in[15:8] ;
assign n1292 =  ( n1291 ) == ( bv_8_124_n462 )  ;
assign n1293 = in[15:8] ;
assign n1294 =  ( n1293 ) == ( bv_8_123_n466 )  ;
assign n1295 = in[15:8] ;
assign n1296 =  ( n1295 ) == ( bv_8_122_n256 )  ;
assign n1297 = in[15:8] ;
assign n1298 =  ( n1297 ) == ( bv_8_121_n301 )  ;
assign n1299 = in[15:8] ;
assign n1300 =  ( n1299 ) == ( bv_8_120_n242 )  ;
assign n1301 = in[15:8] ;
assign n1302 =  ( n1301 ) == ( bv_8_119_n476 )  ;
assign n1303 = in[15:8] ;
assign n1304 =  ( n1303 ) == ( bv_8_118_n479 )  ;
assign n1305 = in[15:8] ;
assign n1306 =  ( n1305 ) == ( bv_8_117_n483 )  ;
assign n1307 = in[15:8] ;
assign n1308 =  ( n1307 ) == ( bv_8_116_n210 )  ;
assign n1309 = in[15:8] ;
assign n1310 =  ( n1309 ) == ( bv_8_115_n407 )  ;
assign n1311 = in[15:8] ;
assign n1312 =  ( n1311 ) == ( bv_8_114_n490 )  ;
assign n1313 = in[15:8] ;
assign n1314 =  ( n1313 ) == ( bv_8_113_n494 )  ;
assign n1315 = in[15:8] ;
assign n1316 =  ( n1315 ) == ( bv_8_112_n187 )  ;
assign n1317 = in[15:8] ;
assign n1318 =  ( n1317 ) == ( bv_8_111_n500 )  ;
assign n1319 = in[15:8] ;
assign n1320 =  ( n1319 ) == ( bv_8_110_n503 )  ;
assign n1321 = in[15:8] ;
assign n1322 =  ( n1321 ) == ( bv_8_109_n288 )  ;
assign n1323 = in[15:8] ;
assign n1324 =  ( n1323 ) == ( bv_8_108_n271 )  ;
assign n1325 = in[15:8] ;
assign n1326 =  ( n1325 ) == ( bv_8_107_n512 )  ;
assign n1327 = in[15:8] ;
assign n1328 =  ( n1327 ) == ( bv_8_106_n515 )  ;
assign n1329 = in[15:8] ;
assign n1330 =  ( n1329 ) == ( bv_8_105_n112 )  ;
assign n1331 = in[15:8] ;
assign n1332 =  ( n1331 ) == ( bv_8_104_n38 )  ;
assign n1333 = in[15:8] ;
assign n1334 =  ( n1333 ) == ( bv_8_103_n524 )  ;
assign n1335 = in[15:8] ;
assign n1336 =  ( n1335 ) == ( bv_8_102_n175 )  ;
assign n1337 = in[15:8] ;
assign n1338 =  ( n1337 ) == ( bv_8_101_n260 )  ;
assign n1339 = in[15:8] ;
assign n1340 =  ( n1339 ) == ( bv_8_100_n416 )  ;
assign n1341 = in[15:8] ;
assign n1342 =  ( n1341 ) == ( bv_8_99_n536 )  ;
assign n1343 = in[15:8] ;
assign n1344 =  ( n1343 ) == ( bv_8_98_n315 )  ;
assign n1345 = in[15:8] ;
assign n1346 =  ( n1345 ) == ( bv_8_97_n156 )  ;
assign n1347 = in[15:8] ;
assign n1348 =  ( n1347 ) == ( bv_8_96_n403 )  ;
assign n1349 = in[15:8] ;
assign n1350 =  ( n1349 ) == ( bv_8_95_n439 )  ;
assign n1351 = in[15:8] ;
assign n1352 =  ( n1351 ) == ( bv_8_94_n362 )  ;
assign n1353 = in[15:8] ;
assign n1354 =  ( n1353 ) == ( bv_8_93_n413 )  ;
assign n1355 = in[15:8] ;
assign n1356 =  ( n1355 ) == ( bv_8_92_n327 )  ;
assign n1357 = in[15:8] ;
assign n1358 =  ( n1357 ) == ( bv_8_91_n556 )  ;
assign n1359 = in[15:8] ;
assign n1360 =  ( n1359 ) == ( bv_8_90_n560 )  ;
assign n1361 = in[15:8] ;
assign n1362 =  ( n1361 ) == ( bv_8_89_n563 )  ;
assign n1363 = in[15:8] ;
assign n1364 =  ( n1363 ) == ( bv_8_88_n548 )  ;
assign n1365 = in[15:8] ;
assign n1366 =  ( n1365 ) == ( bv_8_87_n149 )  ;
assign n1367 = in[15:8] ;
assign n1368 =  ( n1367 ) == ( bv_8_86_n267 )  ;
assign n1369 = in[15:8] ;
assign n1370 =  ( n1369 ) == ( bv_8_85_n78 )  ;
assign n1371 = in[15:8] ;
assign n1372 =  ( n1371 ) == ( bv_8_84_n14 )  ;
assign n1373 = in[15:8] ;
assign n1374 =  ( n1373 ) == ( bv_8_83_n577 )  ;
assign n1375 = in[15:8] ;
assign n1376 =  ( n1375 ) == ( bv_8_82_n580 )  ;
assign n1377 = in[15:8] ;
assign n1378 =  ( n1377 ) == ( bv_8_81_n498 )  ;
assign n1379 = in[15:8] ;
assign n1380 =  ( n1379 ) == ( bv_8_80_n510 )  ;
assign n1381 = in[15:8] ;
assign n1382 =  ( n1381 ) == ( bv_8_79_n397 )  ;
assign n1383 = in[15:8] ;
assign n1384 =  ( n1383 ) == ( bv_8_78_n279 )  ;
assign n1385 = in[15:8] ;
assign n1386 =  ( n1385 ) == ( bv_8_77_n531 )  ;
assign n1387 = in[15:8] ;
assign n1388 =  ( n1387 ) == ( bv_8_76_n551 )  ;
assign n1389 = in[15:8] ;
assign n1390 =  ( n1389 ) == ( bv_8_75_n202 )  ;
assign n1391 = in[15:8] ;
assign n1392 =  ( n1391 ) == ( bv_8_74_n554 )  ;
assign n1393 = in[15:8] ;
assign n1394 =  ( n1393 ) == ( bv_8_73_n338 )  ;
assign n1395 = in[15:8] ;
assign n1396 =  ( n1395 ) == ( bv_8_72_n171 )  ;
assign n1397 = in[15:8] ;
assign n1398 =  ( n1397 ) == ( bv_8_71_n607 )  ;
assign n1399 = in[15:8] ;
assign n1400 =  ( n1399 ) == ( bv_8_70_n376 )  ;
assign n1401 = in[15:8] ;
assign n1402 =  ( n1401 ) == ( bv_8_69_n522 )  ;
assign n1403 = in[15:8] ;
assign n1404 =  ( n1403 ) == ( bv_8_68_n432 )  ;
assign n1405 = in[15:8] ;
assign n1406 =  ( n1405 ) == ( bv_8_67_n534 )  ;
assign n1407 = in[15:8] ;
assign n1408 =  ( n1407 ) == ( bv_8_66_n42 )  ;
assign n1409 = in[15:8] ;
assign n1410 =  ( n1409 ) == ( bv_8_65_n34 )  ;
assign n1411 = in[15:8] ;
assign n1412 =  ( n1411 ) == ( bv_8_64_n492 )  ;
assign n1413 = in[15:8] ;
assign n1414 =  ( n1413 ) == ( bv_8_63_n628 )  ;
assign n1415 = in[15:8] ;
assign n1416 =  ( n1415 ) == ( bv_8_62_n183 )  ;
assign n1417 = in[15:8] ;
assign n1418 =  ( n1417 ) == ( bv_8_61_n419 )  ;
assign n1419 = in[15:8] ;
assign n1420 =  ( n1419 ) == ( bv_8_60_n507 )  ;
assign n1421 = in[15:8] ;
assign n1422 =  ( n1421 ) == ( bv_8_59_n603 )  ;
assign n1423 = in[15:8] ;
assign n1424 =  ( n1423 ) == ( bv_8_58_n346 )  ;
assign n1425 = in[15:8] ;
assign n1426 =  ( n1425 ) == ( bv_8_57_n558 )  ;
assign n1427 = in[15:8] ;
assign n1428 =  ( n1427 ) == ( bv_8_56_n481 )  ;
assign n1429 = in[15:8] ;
assign n1430 =  ( n1429 ) == ( bv_8_55_n292 )  ;
assign n1431 = in[15:8] ;
assign n1432 =  ( n1431 ) == ( bv_8_54_n650 )  ;
assign n1433 = in[15:8] ;
assign n1434 =  ( n1433 ) == ( bv_8_53_n152 )  ;
assign n1435 = in[15:8] ;
assign n1436 =  ( n1435 ) == ( bv_8_52_n656 )  ;
assign n1437 = in[15:8] ;
assign n1438 =  ( n1437 ) == ( bv_8_51_n528 )  ;
assign n1439 = in[15:8] ;
assign n1440 =  ( n1439 ) == ( bv_8_50_n349 )  ;
assign n1441 = in[15:8] ;
assign n1442 =  ( n1441 ) == ( bv_8_49_n665 )  ;
assign n1443 = in[15:8] ;
assign n1444 =  ( n1443 ) == ( bv_8_48_n668 )  ;
assign n1445 = in[15:8] ;
assign n1446 =  ( n1445 ) == ( bv_8_47_n591 )  ;
assign n1447 = in[15:8] ;
assign n1448 =  ( n1447 ) == ( bv_8_46_n235 )  ;
assign n1449 = in[15:8] ;
assign n1450 =  ( n1449 ) == ( bv_8_45_n26 )  ;
assign n1451 = in[15:8] ;
assign n1452 =  ( n1451 ) == ( bv_8_44_n621 )  ;
assign n1453 = in[15:8] ;
assign n1454 =  ( n1453 ) == ( bv_8_43_n681 )  ;
assign n1455 = in[15:8] ;
assign n1456 =  ( n1455 ) == ( bv_8_42_n387 )  ;
assign n1457 = in[15:8] ;
assign n1458 =  ( n1457 ) == ( bv_8_41_n596 )  ;
assign n1459 = in[15:8] ;
assign n1460 =  ( n1459 ) == ( bv_8_40_n74 )  ;
assign n1461 = in[15:8] ;
assign n1462 =  ( n1461 ) == ( bv_8_39_n634 )  ;
assign n1463 = in[15:8] ;
assign n1464 =  ( n1463 ) == ( bv_8_38_n692 )  ;
assign n1465 = in[15:8] ;
assign n1466 =  ( n1465 ) == ( bv_8_37_n239 )  ;
assign n1467 = in[15:8] ;
assign n1468 =  ( n1467 ) == ( bv_8_36_n330 )  ;
assign n1469 = in[15:8] ;
assign n1470 =  ( n1469 ) == ( bv_8_35_n663 )  ;
assign n1471 = in[15:8] ;
assign n1472 =  ( n1471 ) == ( bv_8_34_n390 )  ;
assign n1473 = in[15:8] ;
assign n1474 =  ( n1473 ) == ( bv_8_33_n468 )  ;
assign n1475 = in[15:8] ;
assign n1476 =  ( n1475 ) == ( bv_8_32_n575 )  ;
assign n1477 = in[15:8] ;
assign n1478 =  ( n1477 ) == ( bv_8_31_n206 )  ;
assign n1479 = in[15:8] ;
assign n1480 =  ( n1479 ) == ( bv_8_30_n93 )  ;
assign n1481 = in[15:8] ;
assign n1482 =  ( n1481 ) == ( bv_8_29_n133 )  ;
assign n1483 = in[15:8] ;
assign n1484 =  ( n1483 ) == ( bv_8_28_n231 )  ;
assign n1485 = in[15:8] ;
assign n1486 =  ( n1485 ) == ( bv_8_27_n615 )  ;
assign n1487 = in[15:8] ;
assign n1488 =  ( n1487 ) == ( bv_8_26_n618 )  ;
assign n1489 = in[15:8] ;
assign n1490 =  ( n1489 ) == ( bv_8_25_n410 )  ;
assign n1491 = in[15:8] ;
assign n1492 =  ( n1491 ) == ( bv_8_24_n658 )  ;
assign n1493 = in[15:8] ;
assign n1494 =  ( n1493 ) == ( bv_8_23_n429 )  ;
assign n1495 = in[15:8] ;
assign n1496 =  ( n1495 ) == ( bv_8_22_n6 )  ;
assign n1497 = in[15:8] ;
assign n1498 =  ( n1497 ) == ( bv_8_21_n673 )  ;
assign n1499 = in[15:8] ;
assign n1500 =  ( n1499 ) == ( bv_8_20_n368 )  ;
assign n1501 = in[15:8] ;
assign n1502 =  ( n1501 ) == ( bv_8_19_n446 )  ;
assign n1503 = in[15:8] ;
assign n1504 =  ( n1503 ) == ( bv_8_18_n643 )  ;
assign n1505 = in[15:8] ;
assign n1506 =  ( n1505 ) == ( bv_8_17_n116 )  ;
assign n1507 = in[15:8] ;
assign n1508 =  ( n1507 ) == ( bv_8_16_n464 )  ;
assign n1509 = in[15:8] ;
assign n1510 =  ( n1509 ) == ( bv_8_15_n22 )  ;
assign n1511 = in[15:8] ;
assign n1512 =  ( n1511 ) == ( bv_8_14_n160 )  ;
assign n1513 = in[15:8] ;
assign n1514 =  ( n1513 ) == ( bv_8_13_n54 )  ;
assign n1515 = in[15:8] ;
assign n1516 =  ( n1515 ) == ( bv_8_12_n449 )  ;
assign n1517 = in[15:8] ;
assign n1518 =  ( n1517 ) == ( bv_8_11_n358 )  ;
assign n1519 = in[15:8] ;
assign n1520 =  ( n1519 ) == ( bv_8_10_n342 )  ;
assign n1521 = in[15:8] ;
assign n1522 =  ( n1521 ) == ( bv_8_9_n626 )  ;
assign n1523 = in[15:8] ;
assign n1524 =  ( n1523 ) == ( bv_8_8_n249 )  ;
assign n1525 = in[15:8] ;
assign n1526 =  ( n1525 ) == ( bv_8_7_n646 )  ;
assign n1527 = in[15:8] ;
assign n1528 =  ( n1527 ) == ( bv_8_6_n334 )  ;
assign n1529 = in[15:8] ;
assign n1530 =  ( n1529 ) == ( bv_8_5_n652 )  ;
assign n1531 = in[15:8] ;
assign n1532 =  ( n1531 ) == ( bv_8_4_n670 )  ;
assign n1533 = in[15:8] ;
assign n1534 =  ( n1533 ) == ( bv_8_3_n167 )  ;
assign n1535 = in[15:8] ;
assign n1536 =  ( n1535 ) == ( bv_8_2_n517 )  ;
assign n1537 = in[15:8] ;
assign n1538 =  ( n1537 ) == ( bv_8_1_n752 )  ;
assign n1539 = in[15:8] ;
assign n1540 =  ( n1539 ) == ( bv_8_0_n582 )  ;
assign n1541 =  ( n1540 ) ? ( bv_8_99_n536 ) : ( bv_8_0_n582 ) ;
assign n1542 =  ( n1538 ) ? ( bv_8_124_n462 ) : ( n1541 ) ;
assign n1543 =  ( n1536 ) ? ( bv_8_119_n476 ) : ( n1542 ) ;
assign n1544 =  ( n1534 ) ? ( bv_8_123_n466 ) : ( n1543 ) ;
assign n1545 =  ( n1532 ) ? ( bv_8_242_n56 ) : ( n1544 ) ;
assign n1546 =  ( n1530 ) ? ( bv_8_107_n512 ) : ( n1545 ) ;
assign n1547 =  ( n1528 ) ? ( bv_8_111_n500 ) : ( n1546 ) ;
assign n1548 =  ( n1526 ) ? ( bv_8_197_n225 ) : ( n1547 ) ;
assign n1549 =  ( n1524 ) ? ( bv_8_48_n668 ) : ( n1548 ) ;
assign n1550 =  ( n1522 ) ? ( bv_8_1_n752 ) : ( n1549 ) ;
assign n1551 =  ( n1520 ) ? ( bv_8_103_n524 ) : ( n1550 ) ;
assign n1552 =  ( n1518 ) ? ( bv_8_43_n681 ) : ( n1551 ) ;
assign n1553 =  ( n1516 ) ? ( bv_8_254_n8 ) : ( n1552 ) ;
assign n1554 =  ( n1514 ) ? ( bv_8_215_n158 ) : ( n1553 ) ;
assign n1555 =  ( n1512 ) ? ( bv_8_171_n313 ) : ( n1554 ) ;
assign n1556 =  ( n1510 ) ? ( bv_8_118_n479 ) : ( n1555 ) ;
assign n1557 =  ( n1508 ) ? ( bv_8_202_n208 ) : ( n1556 ) ;
assign n1558 =  ( n1506 ) ? ( bv_8_130_n444 ) : ( n1557 ) ;
assign n1559 =  ( n1504 ) ? ( bv_8_201_n212 ) : ( n1558 ) ;
assign n1560 =  ( n1502 ) ? ( bv_8_125_n459 ) : ( n1559 ) ;
assign n1561 =  ( n1500 ) ? ( bv_8_250_n24 ) : ( n1560 ) ;
assign n1562 =  ( n1498 ) ? ( bv_8_89_n563 ) : ( n1561 ) ;
assign n1563 =  ( n1496 ) ? ( bv_8_71_n607 ) : ( n1562 ) ;
assign n1564 =  ( n1494 ) ? ( bv_8_240_n64 ) : ( n1563 ) ;
assign n1565 =  ( n1492 ) ? ( bv_8_173_n305 ) : ( n1564 ) ;
assign n1566 =  ( n1490 ) ? ( bv_8_212_n169 ) : ( n1565 ) ;
assign n1567 =  ( n1488 ) ? ( bv_8_162_n344 ) : ( n1566 ) ;
assign n1568 =  ( n1486 ) ? ( bv_8_175_n299 ) : ( n1567 ) ;
assign n1569 =  ( n1484 ) ? ( bv_8_156_n364 ) : ( n1568 ) ;
assign n1570 =  ( n1482 ) ? ( bv_8_164_n336 ) : ( n1569 ) ;
assign n1571 =  ( n1480 ) ? ( bv_8_114_n490 ) : ( n1570 ) ;
assign n1572 =  ( n1478 ) ? ( bv_8_192_n244 ) : ( n1571 ) ;
assign n1573 =  ( n1476 ) ? ( bv_8_183_n273 ) : ( n1572 ) ;
assign n1574 =  ( n1474 ) ? ( bv_8_253_n12 ) : ( n1573 ) ;
assign n1575 =  ( n1472 ) ? ( bv_8_147_n392 ) : ( n1574 ) ;
assign n1576 =  ( n1470 ) ? ( bv_8_38_n692 ) : ( n1575 ) ;
assign n1577 =  ( n1468 ) ? ( bv_8_54_n650 ) : ( n1576 ) ;
assign n1578 =  ( n1466 ) ? ( bv_8_63_n628 ) : ( n1577 ) ;
assign n1579 =  ( n1464 ) ? ( bv_8_247_n36 ) : ( n1578 ) ;
assign n1580 =  ( n1462 ) ? ( bv_8_204_n200 ) : ( n1579 ) ;
assign n1581 =  ( n1460 ) ? ( bv_8_52_n656 ) : ( n1580 ) ;
assign n1582 =  ( n1458 ) ? ( bv_8_165_n332 ) : ( n1581 ) ;
assign n1583 =  ( n1456 ) ? ( bv_8_229_n106 ) : ( n1582 ) ;
assign n1584 =  ( n1454 ) ? ( bv_8_241_n60 ) : ( n1583 ) ;
assign n1585 =  ( n1452 ) ? ( bv_8_113_n494 ) : ( n1584 ) ;
assign n1586 =  ( n1450 ) ? ( bv_8_216_n154 ) : ( n1585 ) ;
assign n1587 =  ( n1448 ) ? ( bv_8_49_n665 ) : ( n1586 ) ;
assign n1588 =  ( n1446 ) ? ( bv_8_21_n673 ) : ( n1587 ) ;
assign n1589 =  ( n1444 ) ? ( bv_8_4_n670 ) : ( n1588 ) ;
assign n1590 =  ( n1442 ) ? ( bv_8_199_n218 ) : ( n1589 ) ;
assign n1591 =  ( n1440 ) ? ( bv_8_35_n663 ) : ( n1590 ) ;
assign n1592 =  ( n1438 ) ? ( bv_8_195_n233 ) : ( n1591 ) ;
assign n1593 =  ( n1436 ) ? ( bv_8_24_n658 ) : ( n1592 ) ;
assign n1594 =  ( n1434 ) ? ( bv_8_150_n382 ) : ( n1593 ) ;
assign n1595 =  ( n1432 ) ? ( bv_8_5_n652 ) : ( n1594 ) ;
assign n1596 =  ( n1430 ) ? ( bv_8_154_n370 ) : ( n1595 ) ;
assign n1597 =  ( n1428 ) ? ( bv_8_7_n646 ) : ( n1596 ) ;
assign n1598 =  ( n1426 ) ? ( bv_8_18_n643 ) : ( n1597 ) ;
assign n1599 =  ( n1424 ) ? ( bv_8_128_n451 ) : ( n1598 ) ;
assign n1600 =  ( n1422 ) ? ( bv_8_226_n118 ) : ( n1599 ) ;
assign n1601 =  ( n1420 ) ? ( bv_8_235_n84 ) : ( n1600 ) ;
assign n1602 =  ( n1418 ) ? ( bv_8_39_n634 ) : ( n1601 ) ;
assign n1603 =  ( n1416 ) ? ( bv_8_178_n290 ) : ( n1602 ) ;
assign n1604 =  ( n1414 ) ? ( bv_8_117_n483 ) : ( n1603 ) ;
assign n1605 =  ( n1412 ) ? ( bv_8_9_n626 ) : ( n1604 ) ;
assign n1606 =  ( n1410 ) ? ( bv_8_131_n441 ) : ( n1605 ) ;
assign n1607 =  ( n1408 ) ? ( bv_8_44_n621 ) : ( n1606 ) ;
assign n1608 =  ( n1406 ) ? ( bv_8_26_n618 ) : ( n1607 ) ;
assign n1609 =  ( n1404 ) ? ( bv_8_27_n615 ) : ( n1608 ) ;
assign n1610 =  ( n1402 ) ? ( bv_8_110_n503 ) : ( n1609 ) ;
assign n1611 =  ( n1400 ) ? ( bv_8_90_n560 ) : ( n1610 ) ;
assign n1612 =  ( n1398 ) ? ( bv_8_160_n351 ) : ( n1611 ) ;
assign n1613 =  ( n1396 ) ? ( bv_8_82_n580 ) : ( n1612 ) ;
assign n1614 =  ( n1394 ) ? ( bv_8_59_n603 ) : ( n1613 ) ;
assign n1615 =  ( n1392 ) ? ( bv_8_214_n162 ) : ( n1614 ) ;
assign n1616 =  ( n1390 ) ? ( bv_8_179_n286 ) : ( n1615 ) ;
assign n1617 =  ( n1388 ) ? ( bv_8_41_n596 ) : ( n1616 ) ;
assign n1618 =  ( n1386 ) ? ( bv_8_227_n114 ) : ( n1617 ) ;
assign n1619 =  ( n1384 ) ? ( bv_8_47_n591 ) : ( n1618 ) ;
assign n1620 =  ( n1382 ) ? ( bv_8_132_n437 ) : ( n1619 ) ;
assign n1621 =  ( n1380 ) ? ( bv_8_83_n577 ) : ( n1620 ) ;
assign n1622 =  ( n1378 ) ? ( bv_8_209_n181 ) : ( n1621 ) ;
assign n1623 =  ( n1376 ) ? ( bv_8_0_n582 ) : ( n1622 ) ;
assign n1624 =  ( n1374 ) ? ( bv_8_237_n76 ) : ( n1623 ) ;
assign n1625 =  ( n1372 ) ? ( bv_8_32_n575 ) : ( n1624 ) ;
assign n1626 =  ( n1370 ) ? ( bv_8_252_n16 ) : ( n1625 ) ;
assign n1627 =  ( n1368 ) ? ( bv_8_177_n294 ) : ( n1626 ) ;
assign n1628 =  ( n1366 ) ? ( bv_8_91_n556 ) : ( n1627 ) ;
assign n1629 =  ( n1364 ) ? ( bv_8_106_n515 ) : ( n1628 ) ;
assign n1630 =  ( n1362 ) ? ( bv_8_203_n204 ) : ( n1629 ) ;
assign n1631 =  ( n1360 ) ? ( bv_8_190_n251 ) : ( n1630 ) ;
assign n1632 =  ( n1358 ) ? ( bv_8_57_n558 ) : ( n1631 ) ;
assign n1633 =  ( n1356 ) ? ( bv_8_74_n554 ) : ( n1632 ) ;
assign n1634 =  ( n1354 ) ? ( bv_8_76_n551 ) : ( n1633 ) ;
assign n1635 =  ( n1352 ) ? ( bv_8_88_n548 ) : ( n1634 ) ;
assign n1636 =  ( n1350 ) ? ( bv_8_207_n189 ) : ( n1635 ) ;
assign n1637 =  ( n1348 ) ? ( bv_8_208_n185 ) : ( n1636 ) ;
assign n1638 =  ( n1346 ) ? ( bv_8_239_n68 ) : ( n1637 ) ;
assign n1639 =  ( n1344 ) ? ( bv_8_170_n317 ) : ( n1638 ) ;
assign n1640 =  ( n1342 ) ? ( bv_8_251_n20 ) : ( n1639 ) ;
assign n1641 =  ( n1340 ) ? ( bv_8_67_n534 ) : ( n1640 ) ;
assign n1642 =  ( n1338 ) ? ( bv_8_77_n531 ) : ( n1641 ) ;
assign n1643 =  ( n1336 ) ? ( bv_8_51_n528 ) : ( n1642 ) ;
assign n1644 =  ( n1334 ) ? ( bv_8_133_n434 ) : ( n1643 ) ;
assign n1645 =  ( n1332 ) ? ( bv_8_69_n522 ) : ( n1644 ) ;
assign n1646 =  ( n1330 ) ? ( bv_8_249_n28 ) : ( n1645 ) ;
assign n1647 =  ( n1328 ) ? ( bv_8_2_n517 ) : ( n1646 ) ;
assign n1648 =  ( n1326 ) ? ( bv_8_127_n454 ) : ( n1647 ) ;
assign n1649 =  ( n1324 ) ? ( bv_8_80_n510 ) : ( n1648 ) ;
assign n1650 =  ( n1322 ) ? ( bv_8_60_n507 ) : ( n1649 ) ;
assign n1651 =  ( n1320 ) ? ( bv_8_159_n354 ) : ( n1650 ) ;
assign n1652 =  ( n1318 ) ? ( bv_8_168_n322 ) : ( n1651 ) ;
assign n1653 =  ( n1316 ) ? ( bv_8_81_n498 ) : ( n1652 ) ;
assign n1654 =  ( n1314 ) ? ( bv_8_163_n340 ) : ( n1653 ) ;
assign n1655 =  ( n1312 ) ? ( bv_8_64_n492 ) : ( n1654 ) ;
assign n1656 =  ( n1310 ) ? ( bv_8_143_n405 ) : ( n1655 ) ;
assign n1657 =  ( n1308 ) ? ( bv_8_146_n395 ) : ( n1656 ) ;
assign n1658 =  ( n1306 ) ? ( bv_8_157_n360 ) : ( n1657 ) ;
assign n1659 =  ( n1304 ) ? ( bv_8_56_n481 ) : ( n1658 ) ;
assign n1660 =  ( n1302 ) ? ( bv_8_245_n44 ) : ( n1659 ) ;
assign n1661 =  ( n1300 ) ? ( bv_8_188_n258 ) : ( n1660 ) ;
assign n1662 =  ( n1298 ) ? ( bv_8_182_n277 ) : ( n1661 ) ;
assign n1663 =  ( n1296 ) ? ( bv_8_218_n147 ) : ( n1662 ) ;
assign n1664 =  ( n1294 ) ? ( bv_8_33_n468 ) : ( n1663 ) ;
assign n1665 =  ( n1292 ) ? ( bv_8_16_n464 ) : ( n1664 ) ;
assign n1666 =  ( n1290 ) ? ( bv_8_255_n4 ) : ( n1665 ) ;
assign n1667 =  ( n1288 ) ? ( bv_8_243_n52 ) : ( n1666 ) ;
assign n1668 =  ( n1286 ) ? ( bv_8_210_n177 ) : ( n1667 ) ;
assign n1669 =  ( n1284 ) ? ( bv_8_205_n196 ) : ( n1668 ) ;
assign n1670 =  ( n1282 ) ? ( bv_8_12_n449 ) : ( n1669 ) ;
assign n1671 =  ( n1280 ) ? ( bv_8_19_n446 ) : ( n1670 ) ;
assign n1672 =  ( n1278 ) ? ( bv_8_236_n80 ) : ( n1671 ) ;
assign n1673 =  ( n1276 ) ? ( bv_8_95_n439 ) : ( n1672 ) ;
assign n1674 =  ( n1274 ) ? ( bv_8_151_n378 ) : ( n1673 ) ;
assign n1675 =  ( n1272 ) ? ( bv_8_68_n432 ) : ( n1674 ) ;
assign n1676 =  ( n1270 ) ? ( bv_8_23_n429 ) : ( n1675 ) ;
assign n1677 =  ( n1268 ) ? ( bv_8_196_n229 ) : ( n1676 ) ;
assign n1678 =  ( n1266 ) ? ( bv_8_167_n325 ) : ( n1677 ) ;
assign n1679 =  ( n1264 ) ? ( bv_8_126_n422 ) : ( n1678 ) ;
assign n1680 =  ( n1262 ) ? ( bv_8_61_n419 ) : ( n1679 ) ;
assign n1681 =  ( n1260 ) ? ( bv_8_100_n416 ) : ( n1680 ) ;
assign n1682 =  ( n1258 ) ? ( bv_8_93_n413 ) : ( n1681 ) ;
assign n1683 =  ( n1256 ) ? ( bv_8_25_n410 ) : ( n1682 ) ;
assign n1684 =  ( n1254 ) ? ( bv_8_115_n407 ) : ( n1683 ) ;
assign n1685 =  ( n1252 ) ? ( bv_8_96_n403 ) : ( n1684 ) ;
assign n1686 =  ( n1250 ) ? ( bv_8_129_n400 ) : ( n1685 ) ;
assign n1687 =  ( n1248 ) ? ( bv_8_79_n397 ) : ( n1686 ) ;
assign n1688 =  ( n1246 ) ? ( bv_8_220_n139 ) : ( n1687 ) ;
assign n1689 =  ( n1244 ) ? ( bv_8_34_n390 ) : ( n1688 ) ;
assign n1690 =  ( n1242 ) ? ( bv_8_42_n387 ) : ( n1689 ) ;
assign n1691 =  ( n1240 ) ? ( bv_8_144_n384 ) : ( n1690 ) ;
assign n1692 =  ( n1238 ) ? ( bv_8_136_n380 ) : ( n1691 ) ;
assign n1693 =  ( n1236 ) ? ( bv_8_70_n376 ) : ( n1692 ) ;
assign n1694 =  ( n1234 ) ? ( bv_8_238_n72 ) : ( n1693 ) ;
assign n1695 =  ( n1232 ) ? ( bv_8_184_n269 ) : ( n1694 ) ;
assign n1696 =  ( n1230 ) ? ( bv_8_20_n368 ) : ( n1695 ) ;
assign n1697 =  ( n1228 ) ? ( bv_8_222_n131 ) : ( n1696 ) ;
assign n1698 =  ( n1226 ) ? ( bv_8_94_n362 ) : ( n1697 ) ;
assign n1699 =  ( n1224 ) ? ( bv_8_11_n358 ) : ( n1698 ) ;
assign n1700 =  ( n1222 ) ? ( bv_8_219_n143 ) : ( n1699 ) ;
assign n1701 =  ( n1220 ) ? ( bv_8_224_n125 ) : ( n1700 ) ;
assign n1702 =  ( n1218 ) ? ( bv_8_50_n349 ) : ( n1701 ) ;
assign n1703 =  ( n1216 ) ? ( bv_8_58_n346 ) : ( n1702 ) ;
assign n1704 =  ( n1214 ) ? ( bv_8_10_n342 ) : ( n1703 ) ;
assign n1705 =  ( n1212 ) ? ( bv_8_73_n338 ) : ( n1704 ) ;
assign n1706 =  ( n1210 ) ? ( bv_8_6_n334 ) : ( n1705 ) ;
assign n1707 =  ( n1208 ) ? ( bv_8_36_n330 ) : ( n1706 ) ;
assign n1708 =  ( n1206 ) ? ( bv_8_92_n327 ) : ( n1707 ) ;
assign n1709 =  ( n1204 ) ? ( bv_8_194_n237 ) : ( n1708 ) ;
assign n1710 =  ( n1202 ) ? ( bv_8_211_n173 ) : ( n1709 ) ;
assign n1711 =  ( n1200 ) ? ( bv_8_172_n309 ) : ( n1710 ) ;
assign n1712 =  ( n1198 ) ? ( bv_8_98_n315 ) : ( n1711 ) ;
assign n1713 =  ( n1196 ) ? ( bv_8_145_n311 ) : ( n1712 ) ;
assign n1714 =  ( n1194 ) ? ( bv_8_149_n307 ) : ( n1713 ) ;
assign n1715 =  ( n1192 ) ? ( bv_8_228_n110 ) : ( n1714 ) ;
assign n1716 =  ( n1190 ) ? ( bv_8_121_n301 ) : ( n1715 ) ;
assign n1717 =  ( n1188 ) ? ( bv_8_231_n99 ) : ( n1716 ) ;
assign n1718 =  ( n1186 ) ? ( bv_8_200_n215 ) : ( n1717 ) ;
assign n1719 =  ( n1184 ) ? ( bv_8_55_n292 ) : ( n1718 ) ;
assign n1720 =  ( n1182 ) ? ( bv_8_109_n288 ) : ( n1719 ) ;
assign n1721 =  ( n1180 ) ? ( bv_8_141_n284 ) : ( n1720 ) ;
assign n1722 =  ( n1178 ) ? ( bv_8_213_n165 ) : ( n1721 ) ;
assign n1723 =  ( n1176 ) ? ( bv_8_78_n279 ) : ( n1722 ) ;
assign n1724 =  ( n1174 ) ? ( bv_8_169_n275 ) : ( n1723 ) ;
assign n1725 =  ( n1172 ) ? ( bv_8_108_n271 ) : ( n1724 ) ;
assign n1726 =  ( n1170 ) ? ( bv_8_86_n267 ) : ( n1725 ) ;
assign n1727 =  ( n1168 ) ? ( bv_8_244_n48 ) : ( n1726 ) ;
assign n1728 =  ( n1166 ) ? ( bv_8_234_n88 ) : ( n1727 ) ;
assign n1729 =  ( n1164 ) ? ( bv_8_101_n260 ) : ( n1728 ) ;
assign n1730 =  ( n1162 ) ? ( bv_8_122_n256 ) : ( n1729 ) ;
assign n1731 =  ( n1160 ) ? ( bv_8_174_n253 ) : ( n1730 ) ;
assign n1732 =  ( n1158 ) ? ( bv_8_8_n249 ) : ( n1731 ) ;
assign n1733 =  ( n1156 ) ? ( bv_8_186_n246 ) : ( n1732 ) ;
assign n1734 =  ( n1154 ) ? ( bv_8_120_n242 ) : ( n1733 ) ;
assign n1735 =  ( n1152 ) ? ( bv_8_37_n239 ) : ( n1734 ) ;
assign n1736 =  ( n1150 ) ? ( bv_8_46_n235 ) : ( n1735 ) ;
assign n1737 =  ( n1148 ) ? ( bv_8_28_n231 ) : ( n1736 ) ;
assign n1738 =  ( n1146 ) ? ( bv_8_166_n227 ) : ( n1737 ) ;
assign n1739 =  ( n1144 ) ? ( bv_8_180_n223 ) : ( n1738 ) ;
assign n1740 =  ( n1142 ) ? ( bv_8_198_n220 ) : ( n1739 ) ;
assign n1741 =  ( n1140 ) ? ( bv_8_232_n95 ) : ( n1740 ) ;
assign n1742 =  ( n1138 ) ? ( bv_8_221_n135 ) : ( n1741 ) ;
assign n1743 =  ( n1136 ) ? ( bv_8_116_n210 ) : ( n1742 ) ;
assign n1744 =  ( n1134 ) ? ( bv_8_31_n206 ) : ( n1743 ) ;
assign n1745 =  ( n1132 ) ? ( bv_8_75_n202 ) : ( n1744 ) ;
assign n1746 =  ( n1130 ) ? ( bv_8_189_n198 ) : ( n1745 ) ;
assign n1747 =  ( n1128 ) ? ( bv_8_139_n194 ) : ( n1746 ) ;
assign n1748 =  ( n1126 ) ? ( bv_8_138_n191 ) : ( n1747 ) ;
assign n1749 =  ( n1124 ) ? ( bv_8_112_n187 ) : ( n1748 ) ;
assign n1750 =  ( n1122 ) ? ( bv_8_62_n183 ) : ( n1749 ) ;
assign n1751 =  ( n1120 ) ? ( bv_8_181_n179 ) : ( n1750 ) ;
assign n1752 =  ( n1118 ) ? ( bv_8_102_n175 ) : ( n1751 ) ;
assign n1753 =  ( n1116 ) ? ( bv_8_72_n171 ) : ( n1752 ) ;
assign n1754 =  ( n1114 ) ? ( bv_8_3_n167 ) : ( n1753 ) ;
assign n1755 =  ( n1112 ) ? ( bv_8_246_n40 ) : ( n1754 ) ;
assign n1756 =  ( n1110 ) ? ( bv_8_14_n160 ) : ( n1755 ) ;
assign n1757 =  ( n1108 ) ? ( bv_8_97_n156 ) : ( n1756 ) ;
assign n1758 =  ( n1106 ) ? ( bv_8_53_n152 ) : ( n1757 ) ;
assign n1759 =  ( n1104 ) ? ( bv_8_87_n149 ) : ( n1758 ) ;
assign n1760 =  ( n1102 ) ? ( bv_8_185_n145 ) : ( n1759 ) ;
assign n1761 =  ( n1100 ) ? ( bv_8_134_n141 ) : ( n1760 ) ;
assign n1762 =  ( n1098 ) ? ( bv_8_193_n137 ) : ( n1761 ) ;
assign n1763 =  ( n1096 ) ? ( bv_8_29_n133 ) : ( n1762 ) ;
assign n1764 =  ( n1094 ) ? ( bv_8_158_n129 ) : ( n1763 ) ;
assign n1765 =  ( n1092 ) ? ( bv_8_225_n122 ) : ( n1764 ) ;
assign n1766 =  ( n1090 ) ? ( bv_8_248_n32 ) : ( n1765 ) ;
assign n1767 =  ( n1088 ) ? ( bv_8_152_n120 ) : ( n1766 ) ;
assign n1768 =  ( n1086 ) ? ( bv_8_17_n116 ) : ( n1767 ) ;
assign n1769 =  ( n1084 ) ? ( bv_8_105_n112 ) : ( n1768 ) ;
assign n1770 =  ( n1082 ) ? ( bv_8_217_n108 ) : ( n1769 ) ;
assign n1771 =  ( n1080 ) ? ( bv_8_142_n104 ) : ( n1770 ) ;
assign n1772 =  ( n1078 ) ? ( bv_8_148_n101 ) : ( n1771 ) ;
assign n1773 =  ( n1076 ) ? ( bv_8_155_n97 ) : ( n1772 ) ;
assign n1774 =  ( n1074 ) ? ( bv_8_30_n93 ) : ( n1773 ) ;
assign n1775 =  ( n1072 ) ? ( bv_8_135_n90 ) : ( n1774 ) ;
assign n1776 =  ( n1070 ) ? ( bv_8_233_n86 ) : ( n1775 ) ;
assign n1777 =  ( n1068 ) ? ( bv_8_206_n82 ) : ( n1776 ) ;
assign n1778 =  ( n1066 ) ? ( bv_8_85_n78 ) : ( n1777 ) ;
assign n1779 =  ( n1064 ) ? ( bv_8_40_n74 ) : ( n1778 ) ;
assign n1780 =  ( n1062 ) ? ( bv_8_223_n70 ) : ( n1779 ) ;
assign n1781 =  ( n1060 ) ? ( bv_8_140_n66 ) : ( n1780 ) ;
assign n1782 =  ( n1058 ) ? ( bv_8_161_n62 ) : ( n1781 ) ;
assign n1783 =  ( n1056 ) ? ( bv_8_137_n58 ) : ( n1782 ) ;
assign n1784 =  ( n1054 ) ? ( bv_8_13_n54 ) : ( n1783 ) ;
assign n1785 =  ( n1052 ) ? ( bv_8_191_n50 ) : ( n1784 ) ;
assign n1786 =  ( n1050 ) ? ( bv_8_230_n46 ) : ( n1785 ) ;
assign n1787 =  ( n1048 ) ? ( bv_8_66_n42 ) : ( n1786 ) ;
assign n1788 =  ( n1046 ) ? ( bv_8_104_n38 ) : ( n1787 ) ;
assign n1789 =  ( n1044 ) ? ( bv_8_65_n34 ) : ( n1788 ) ;
assign n1790 =  ( n1042 ) ? ( bv_8_153_n30 ) : ( n1789 ) ;
assign n1791 =  ( n1040 ) ? ( bv_8_45_n26 ) : ( n1790 ) ;
assign n1792 =  ( n1038 ) ? ( bv_8_15_n22 ) : ( n1791 ) ;
assign n1793 =  ( n1036 ) ? ( bv_8_176_n18 ) : ( n1792 ) ;
assign n1794 =  ( n1034 ) ? ( bv_8_84_n14 ) : ( n1793 ) ;
assign n1795 =  ( n1032 ) ? ( bv_8_187_n10 ) : ( n1794 ) ;
assign n1796 =  ( n1030 ) ? ( bv_8_22_n6 ) : ( n1795 ) ;
assign n1797 =  ( n1028 ) ^ ( n1796 )  ;
assign n1798 =  { ( n1027 ) , ( n1797 ) }  ;
assign n1799 = in[111:104] ;
assign n1800 = in[7:0] ;
assign n1801 =  ( n1800 ) == ( bv_8_255_n4 )  ;
assign n1802 = in[7:0] ;
assign n1803 =  ( n1802 ) == ( bv_8_254_n8 )  ;
assign n1804 = in[7:0] ;
assign n1805 =  ( n1804 ) == ( bv_8_253_n12 )  ;
assign n1806 = in[7:0] ;
assign n1807 =  ( n1806 ) == ( bv_8_252_n16 )  ;
assign n1808 = in[7:0] ;
assign n1809 =  ( n1808 ) == ( bv_8_251_n20 )  ;
assign n1810 = in[7:0] ;
assign n1811 =  ( n1810 ) == ( bv_8_250_n24 )  ;
assign n1812 = in[7:0] ;
assign n1813 =  ( n1812 ) == ( bv_8_249_n28 )  ;
assign n1814 = in[7:0] ;
assign n1815 =  ( n1814 ) == ( bv_8_248_n32 )  ;
assign n1816 = in[7:0] ;
assign n1817 =  ( n1816 ) == ( bv_8_247_n36 )  ;
assign n1818 = in[7:0] ;
assign n1819 =  ( n1818 ) == ( bv_8_246_n40 )  ;
assign n1820 = in[7:0] ;
assign n1821 =  ( n1820 ) == ( bv_8_245_n44 )  ;
assign n1822 = in[7:0] ;
assign n1823 =  ( n1822 ) == ( bv_8_244_n48 )  ;
assign n1824 = in[7:0] ;
assign n1825 =  ( n1824 ) == ( bv_8_243_n52 )  ;
assign n1826 = in[7:0] ;
assign n1827 =  ( n1826 ) == ( bv_8_242_n56 )  ;
assign n1828 = in[7:0] ;
assign n1829 =  ( n1828 ) == ( bv_8_241_n60 )  ;
assign n1830 = in[7:0] ;
assign n1831 =  ( n1830 ) == ( bv_8_240_n64 )  ;
assign n1832 = in[7:0] ;
assign n1833 =  ( n1832 ) == ( bv_8_239_n68 )  ;
assign n1834 = in[7:0] ;
assign n1835 =  ( n1834 ) == ( bv_8_238_n72 )  ;
assign n1836 = in[7:0] ;
assign n1837 =  ( n1836 ) == ( bv_8_237_n76 )  ;
assign n1838 = in[7:0] ;
assign n1839 =  ( n1838 ) == ( bv_8_236_n80 )  ;
assign n1840 = in[7:0] ;
assign n1841 =  ( n1840 ) == ( bv_8_235_n84 )  ;
assign n1842 = in[7:0] ;
assign n1843 =  ( n1842 ) == ( bv_8_234_n88 )  ;
assign n1844 = in[7:0] ;
assign n1845 =  ( n1844 ) == ( bv_8_233_n86 )  ;
assign n1846 = in[7:0] ;
assign n1847 =  ( n1846 ) == ( bv_8_232_n95 )  ;
assign n1848 = in[7:0] ;
assign n1849 =  ( n1848 ) == ( bv_8_231_n99 )  ;
assign n1850 = in[7:0] ;
assign n1851 =  ( n1850 ) == ( bv_8_230_n46 )  ;
assign n1852 = in[7:0] ;
assign n1853 =  ( n1852 ) == ( bv_8_229_n106 )  ;
assign n1854 = in[7:0] ;
assign n1855 =  ( n1854 ) == ( bv_8_228_n110 )  ;
assign n1856 = in[7:0] ;
assign n1857 =  ( n1856 ) == ( bv_8_227_n114 )  ;
assign n1858 = in[7:0] ;
assign n1859 =  ( n1858 ) == ( bv_8_226_n118 )  ;
assign n1860 = in[7:0] ;
assign n1861 =  ( n1860 ) == ( bv_8_225_n122 )  ;
assign n1862 = in[7:0] ;
assign n1863 =  ( n1862 ) == ( bv_8_224_n125 )  ;
assign n1864 = in[7:0] ;
assign n1865 =  ( n1864 ) == ( bv_8_223_n70 )  ;
assign n1866 = in[7:0] ;
assign n1867 =  ( n1866 ) == ( bv_8_222_n131 )  ;
assign n1868 = in[7:0] ;
assign n1869 =  ( n1868 ) == ( bv_8_221_n135 )  ;
assign n1870 = in[7:0] ;
assign n1871 =  ( n1870 ) == ( bv_8_220_n139 )  ;
assign n1872 = in[7:0] ;
assign n1873 =  ( n1872 ) == ( bv_8_219_n143 )  ;
assign n1874 = in[7:0] ;
assign n1875 =  ( n1874 ) == ( bv_8_218_n147 )  ;
assign n1876 = in[7:0] ;
assign n1877 =  ( n1876 ) == ( bv_8_217_n108 )  ;
assign n1878 = in[7:0] ;
assign n1879 =  ( n1878 ) == ( bv_8_216_n154 )  ;
assign n1880 = in[7:0] ;
assign n1881 =  ( n1880 ) == ( bv_8_215_n158 )  ;
assign n1882 = in[7:0] ;
assign n1883 =  ( n1882 ) == ( bv_8_214_n162 )  ;
assign n1884 = in[7:0] ;
assign n1885 =  ( n1884 ) == ( bv_8_213_n165 )  ;
assign n1886 = in[7:0] ;
assign n1887 =  ( n1886 ) == ( bv_8_212_n169 )  ;
assign n1888 = in[7:0] ;
assign n1889 =  ( n1888 ) == ( bv_8_211_n173 )  ;
assign n1890 = in[7:0] ;
assign n1891 =  ( n1890 ) == ( bv_8_210_n177 )  ;
assign n1892 = in[7:0] ;
assign n1893 =  ( n1892 ) == ( bv_8_209_n181 )  ;
assign n1894 = in[7:0] ;
assign n1895 =  ( n1894 ) == ( bv_8_208_n185 )  ;
assign n1896 = in[7:0] ;
assign n1897 =  ( n1896 ) == ( bv_8_207_n189 )  ;
assign n1898 = in[7:0] ;
assign n1899 =  ( n1898 ) == ( bv_8_206_n82 )  ;
assign n1900 = in[7:0] ;
assign n1901 =  ( n1900 ) == ( bv_8_205_n196 )  ;
assign n1902 = in[7:0] ;
assign n1903 =  ( n1902 ) == ( bv_8_204_n200 )  ;
assign n1904 = in[7:0] ;
assign n1905 =  ( n1904 ) == ( bv_8_203_n204 )  ;
assign n1906 = in[7:0] ;
assign n1907 =  ( n1906 ) == ( bv_8_202_n208 )  ;
assign n1908 = in[7:0] ;
assign n1909 =  ( n1908 ) == ( bv_8_201_n212 )  ;
assign n1910 = in[7:0] ;
assign n1911 =  ( n1910 ) == ( bv_8_200_n215 )  ;
assign n1912 = in[7:0] ;
assign n1913 =  ( n1912 ) == ( bv_8_199_n218 )  ;
assign n1914 = in[7:0] ;
assign n1915 =  ( n1914 ) == ( bv_8_198_n220 )  ;
assign n1916 = in[7:0] ;
assign n1917 =  ( n1916 ) == ( bv_8_197_n225 )  ;
assign n1918 = in[7:0] ;
assign n1919 =  ( n1918 ) == ( bv_8_196_n229 )  ;
assign n1920 = in[7:0] ;
assign n1921 =  ( n1920 ) == ( bv_8_195_n233 )  ;
assign n1922 = in[7:0] ;
assign n1923 =  ( n1922 ) == ( bv_8_194_n237 )  ;
assign n1924 = in[7:0] ;
assign n1925 =  ( n1924 ) == ( bv_8_193_n137 )  ;
assign n1926 = in[7:0] ;
assign n1927 =  ( n1926 ) == ( bv_8_192_n244 )  ;
assign n1928 = in[7:0] ;
assign n1929 =  ( n1928 ) == ( bv_8_191_n50 )  ;
assign n1930 = in[7:0] ;
assign n1931 =  ( n1930 ) == ( bv_8_190_n251 )  ;
assign n1932 = in[7:0] ;
assign n1933 =  ( n1932 ) == ( bv_8_189_n198 )  ;
assign n1934 = in[7:0] ;
assign n1935 =  ( n1934 ) == ( bv_8_188_n258 )  ;
assign n1936 = in[7:0] ;
assign n1937 =  ( n1936 ) == ( bv_8_187_n10 )  ;
assign n1938 = in[7:0] ;
assign n1939 =  ( n1938 ) == ( bv_8_186_n246 )  ;
assign n1940 = in[7:0] ;
assign n1941 =  ( n1940 ) == ( bv_8_185_n145 )  ;
assign n1942 = in[7:0] ;
assign n1943 =  ( n1942 ) == ( bv_8_184_n269 )  ;
assign n1944 = in[7:0] ;
assign n1945 =  ( n1944 ) == ( bv_8_183_n273 )  ;
assign n1946 = in[7:0] ;
assign n1947 =  ( n1946 ) == ( bv_8_182_n277 )  ;
assign n1948 = in[7:0] ;
assign n1949 =  ( n1948 ) == ( bv_8_181_n179 )  ;
assign n1950 = in[7:0] ;
assign n1951 =  ( n1950 ) == ( bv_8_180_n223 )  ;
assign n1952 = in[7:0] ;
assign n1953 =  ( n1952 ) == ( bv_8_179_n286 )  ;
assign n1954 = in[7:0] ;
assign n1955 =  ( n1954 ) == ( bv_8_178_n290 )  ;
assign n1956 = in[7:0] ;
assign n1957 =  ( n1956 ) == ( bv_8_177_n294 )  ;
assign n1958 = in[7:0] ;
assign n1959 =  ( n1958 ) == ( bv_8_176_n18 )  ;
assign n1960 = in[7:0] ;
assign n1961 =  ( n1960 ) == ( bv_8_175_n299 )  ;
assign n1962 = in[7:0] ;
assign n1963 =  ( n1962 ) == ( bv_8_174_n253 )  ;
assign n1964 = in[7:0] ;
assign n1965 =  ( n1964 ) == ( bv_8_173_n305 )  ;
assign n1966 = in[7:0] ;
assign n1967 =  ( n1966 ) == ( bv_8_172_n309 )  ;
assign n1968 = in[7:0] ;
assign n1969 =  ( n1968 ) == ( bv_8_171_n313 )  ;
assign n1970 = in[7:0] ;
assign n1971 =  ( n1970 ) == ( bv_8_170_n317 )  ;
assign n1972 = in[7:0] ;
assign n1973 =  ( n1972 ) == ( bv_8_169_n275 )  ;
assign n1974 = in[7:0] ;
assign n1975 =  ( n1974 ) == ( bv_8_168_n322 )  ;
assign n1976 = in[7:0] ;
assign n1977 =  ( n1976 ) == ( bv_8_167_n325 )  ;
assign n1978 = in[7:0] ;
assign n1979 =  ( n1978 ) == ( bv_8_166_n227 )  ;
assign n1980 = in[7:0] ;
assign n1981 =  ( n1980 ) == ( bv_8_165_n332 )  ;
assign n1982 = in[7:0] ;
assign n1983 =  ( n1982 ) == ( bv_8_164_n336 )  ;
assign n1984 = in[7:0] ;
assign n1985 =  ( n1984 ) == ( bv_8_163_n340 )  ;
assign n1986 = in[7:0] ;
assign n1987 =  ( n1986 ) == ( bv_8_162_n344 )  ;
assign n1988 = in[7:0] ;
assign n1989 =  ( n1988 ) == ( bv_8_161_n62 )  ;
assign n1990 = in[7:0] ;
assign n1991 =  ( n1990 ) == ( bv_8_160_n351 )  ;
assign n1992 = in[7:0] ;
assign n1993 =  ( n1992 ) == ( bv_8_159_n354 )  ;
assign n1994 = in[7:0] ;
assign n1995 =  ( n1994 ) == ( bv_8_158_n129 )  ;
assign n1996 = in[7:0] ;
assign n1997 =  ( n1996 ) == ( bv_8_157_n360 )  ;
assign n1998 = in[7:0] ;
assign n1999 =  ( n1998 ) == ( bv_8_156_n364 )  ;
assign n2000 = in[7:0] ;
assign n2001 =  ( n2000 ) == ( bv_8_155_n97 )  ;
assign n2002 = in[7:0] ;
assign n2003 =  ( n2002 ) == ( bv_8_154_n370 )  ;
assign n2004 = in[7:0] ;
assign n2005 =  ( n2004 ) == ( bv_8_153_n30 )  ;
assign n2006 = in[7:0] ;
assign n2007 =  ( n2006 ) == ( bv_8_152_n120 )  ;
assign n2008 = in[7:0] ;
assign n2009 =  ( n2008 ) == ( bv_8_151_n378 )  ;
assign n2010 = in[7:0] ;
assign n2011 =  ( n2010 ) == ( bv_8_150_n382 )  ;
assign n2012 = in[7:0] ;
assign n2013 =  ( n2012 ) == ( bv_8_149_n307 )  ;
assign n2014 = in[7:0] ;
assign n2015 =  ( n2014 ) == ( bv_8_148_n101 )  ;
assign n2016 = in[7:0] ;
assign n2017 =  ( n2016 ) == ( bv_8_147_n392 )  ;
assign n2018 = in[7:0] ;
assign n2019 =  ( n2018 ) == ( bv_8_146_n395 )  ;
assign n2020 = in[7:0] ;
assign n2021 =  ( n2020 ) == ( bv_8_145_n311 )  ;
assign n2022 = in[7:0] ;
assign n2023 =  ( n2022 ) == ( bv_8_144_n384 )  ;
assign n2024 = in[7:0] ;
assign n2025 =  ( n2024 ) == ( bv_8_143_n405 )  ;
assign n2026 = in[7:0] ;
assign n2027 =  ( n2026 ) == ( bv_8_142_n104 )  ;
assign n2028 = in[7:0] ;
assign n2029 =  ( n2028 ) == ( bv_8_141_n284 )  ;
assign n2030 = in[7:0] ;
assign n2031 =  ( n2030 ) == ( bv_8_140_n66 )  ;
assign n2032 = in[7:0] ;
assign n2033 =  ( n2032 ) == ( bv_8_139_n194 )  ;
assign n2034 = in[7:0] ;
assign n2035 =  ( n2034 ) == ( bv_8_138_n191 )  ;
assign n2036 = in[7:0] ;
assign n2037 =  ( n2036 ) == ( bv_8_137_n58 )  ;
assign n2038 = in[7:0] ;
assign n2039 =  ( n2038 ) == ( bv_8_136_n380 )  ;
assign n2040 = in[7:0] ;
assign n2041 =  ( n2040 ) == ( bv_8_135_n90 )  ;
assign n2042 = in[7:0] ;
assign n2043 =  ( n2042 ) == ( bv_8_134_n141 )  ;
assign n2044 = in[7:0] ;
assign n2045 =  ( n2044 ) == ( bv_8_133_n434 )  ;
assign n2046 = in[7:0] ;
assign n2047 =  ( n2046 ) == ( bv_8_132_n437 )  ;
assign n2048 = in[7:0] ;
assign n2049 =  ( n2048 ) == ( bv_8_131_n441 )  ;
assign n2050 = in[7:0] ;
assign n2051 =  ( n2050 ) == ( bv_8_130_n444 )  ;
assign n2052 = in[7:0] ;
assign n2053 =  ( n2052 ) == ( bv_8_129_n400 )  ;
assign n2054 = in[7:0] ;
assign n2055 =  ( n2054 ) == ( bv_8_128_n451 )  ;
assign n2056 = in[7:0] ;
assign n2057 =  ( n2056 ) == ( bv_8_127_n454 )  ;
assign n2058 = in[7:0] ;
assign n2059 =  ( n2058 ) == ( bv_8_126_n422 )  ;
assign n2060 = in[7:0] ;
assign n2061 =  ( n2060 ) == ( bv_8_125_n459 )  ;
assign n2062 = in[7:0] ;
assign n2063 =  ( n2062 ) == ( bv_8_124_n462 )  ;
assign n2064 = in[7:0] ;
assign n2065 =  ( n2064 ) == ( bv_8_123_n466 )  ;
assign n2066 = in[7:0] ;
assign n2067 =  ( n2066 ) == ( bv_8_122_n256 )  ;
assign n2068 = in[7:0] ;
assign n2069 =  ( n2068 ) == ( bv_8_121_n301 )  ;
assign n2070 = in[7:0] ;
assign n2071 =  ( n2070 ) == ( bv_8_120_n242 )  ;
assign n2072 = in[7:0] ;
assign n2073 =  ( n2072 ) == ( bv_8_119_n476 )  ;
assign n2074 = in[7:0] ;
assign n2075 =  ( n2074 ) == ( bv_8_118_n479 )  ;
assign n2076 = in[7:0] ;
assign n2077 =  ( n2076 ) == ( bv_8_117_n483 )  ;
assign n2078 = in[7:0] ;
assign n2079 =  ( n2078 ) == ( bv_8_116_n210 )  ;
assign n2080 = in[7:0] ;
assign n2081 =  ( n2080 ) == ( bv_8_115_n407 )  ;
assign n2082 = in[7:0] ;
assign n2083 =  ( n2082 ) == ( bv_8_114_n490 )  ;
assign n2084 = in[7:0] ;
assign n2085 =  ( n2084 ) == ( bv_8_113_n494 )  ;
assign n2086 = in[7:0] ;
assign n2087 =  ( n2086 ) == ( bv_8_112_n187 )  ;
assign n2088 = in[7:0] ;
assign n2089 =  ( n2088 ) == ( bv_8_111_n500 )  ;
assign n2090 = in[7:0] ;
assign n2091 =  ( n2090 ) == ( bv_8_110_n503 )  ;
assign n2092 = in[7:0] ;
assign n2093 =  ( n2092 ) == ( bv_8_109_n288 )  ;
assign n2094 = in[7:0] ;
assign n2095 =  ( n2094 ) == ( bv_8_108_n271 )  ;
assign n2096 = in[7:0] ;
assign n2097 =  ( n2096 ) == ( bv_8_107_n512 )  ;
assign n2098 = in[7:0] ;
assign n2099 =  ( n2098 ) == ( bv_8_106_n515 )  ;
assign n2100 = in[7:0] ;
assign n2101 =  ( n2100 ) == ( bv_8_105_n112 )  ;
assign n2102 = in[7:0] ;
assign n2103 =  ( n2102 ) == ( bv_8_104_n38 )  ;
assign n2104 = in[7:0] ;
assign n2105 =  ( n2104 ) == ( bv_8_103_n524 )  ;
assign n2106 = in[7:0] ;
assign n2107 =  ( n2106 ) == ( bv_8_102_n175 )  ;
assign n2108 = in[7:0] ;
assign n2109 =  ( n2108 ) == ( bv_8_101_n260 )  ;
assign n2110 = in[7:0] ;
assign n2111 =  ( n2110 ) == ( bv_8_100_n416 )  ;
assign n2112 = in[7:0] ;
assign n2113 =  ( n2112 ) == ( bv_8_99_n536 )  ;
assign n2114 = in[7:0] ;
assign n2115 =  ( n2114 ) == ( bv_8_98_n315 )  ;
assign n2116 = in[7:0] ;
assign n2117 =  ( n2116 ) == ( bv_8_97_n156 )  ;
assign n2118 = in[7:0] ;
assign n2119 =  ( n2118 ) == ( bv_8_96_n403 )  ;
assign n2120 = in[7:0] ;
assign n2121 =  ( n2120 ) == ( bv_8_95_n439 )  ;
assign n2122 = in[7:0] ;
assign n2123 =  ( n2122 ) == ( bv_8_94_n362 )  ;
assign n2124 = in[7:0] ;
assign n2125 =  ( n2124 ) == ( bv_8_93_n413 )  ;
assign n2126 = in[7:0] ;
assign n2127 =  ( n2126 ) == ( bv_8_92_n327 )  ;
assign n2128 = in[7:0] ;
assign n2129 =  ( n2128 ) == ( bv_8_91_n556 )  ;
assign n2130 = in[7:0] ;
assign n2131 =  ( n2130 ) == ( bv_8_90_n560 )  ;
assign n2132 = in[7:0] ;
assign n2133 =  ( n2132 ) == ( bv_8_89_n563 )  ;
assign n2134 = in[7:0] ;
assign n2135 =  ( n2134 ) == ( bv_8_88_n548 )  ;
assign n2136 = in[7:0] ;
assign n2137 =  ( n2136 ) == ( bv_8_87_n149 )  ;
assign n2138 = in[7:0] ;
assign n2139 =  ( n2138 ) == ( bv_8_86_n267 )  ;
assign n2140 = in[7:0] ;
assign n2141 =  ( n2140 ) == ( bv_8_85_n78 )  ;
assign n2142 = in[7:0] ;
assign n2143 =  ( n2142 ) == ( bv_8_84_n14 )  ;
assign n2144 = in[7:0] ;
assign n2145 =  ( n2144 ) == ( bv_8_83_n577 )  ;
assign n2146 = in[7:0] ;
assign n2147 =  ( n2146 ) == ( bv_8_82_n580 )  ;
assign n2148 = in[7:0] ;
assign n2149 =  ( n2148 ) == ( bv_8_81_n498 )  ;
assign n2150 = in[7:0] ;
assign n2151 =  ( n2150 ) == ( bv_8_80_n510 )  ;
assign n2152 = in[7:0] ;
assign n2153 =  ( n2152 ) == ( bv_8_79_n397 )  ;
assign n2154 = in[7:0] ;
assign n2155 =  ( n2154 ) == ( bv_8_78_n279 )  ;
assign n2156 = in[7:0] ;
assign n2157 =  ( n2156 ) == ( bv_8_77_n531 )  ;
assign n2158 = in[7:0] ;
assign n2159 =  ( n2158 ) == ( bv_8_76_n551 )  ;
assign n2160 = in[7:0] ;
assign n2161 =  ( n2160 ) == ( bv_8_75_n202 )  ;
assign n2162 = in[7:0] ;
assign n2163 =  ( n2162 ) == ( bv_8_74_n554 )  ;
assign n2164 = in[7:0] ;
assign n2165 =  ( n2164 ) == ( bv_8_73_n338 )  ;
assign n2166 = in[7:0] ;
assign n2167 =  ( n2166 ) == ( bv_8_72_n171 )  ;
assign n2168 = in[7:0] ;
assign n2169 =  ( n2168 ) == ( bv_8_71_n607 )  ;
assign n2170 = in[7:0] ;
assign n2171 =  ( n2170 ) == ( bv_8_70_n376 )  ;
assign n2172 = in[7:0] ;
assign n2173 =  ( n2172 ) == ( bv_8_69_n522 )  ;
assign n2174 = in[7:0] ;
assign n2175 =  ( n2174 ) == ( bv_8_68_n432 )  ;
assign n2176 = in[7:0] ;
assign n2177 =  ( n2176 ) == ( bv_8_67_n534 )  ;
assign n2178 = in[7:0] ;
assign n2179 =  ( n2178 ) == ( bv_8_66_n42 )  ;
assign n2180 = in[7:0] ;
assign n2181 =  ( n2180 ) == ( bv_8_65_n34 )  ;
assign n2182 = in[7:0] ;
assign n2183 =  ( n2182 ) == ( bv_8_64_n492 )  ;
assign n2184 = in[7:0] ;
assign n2185 =  ( n2184 ) == ( bv_8_63_n628 )  ;
assign n2186 = in[7:0] ;
assign n2187 =  ( n2186 ) == ( bv_8_62_n183 )  ;
assign n2188 = in[7:0] ;
assign n2189 =  ( n2188 ) == ( bv_8_61_n419 )  ;
assign n2190 = in[7:0] ;
assign n2191 =  ( n2190 ) == ( bv_8_60_n507 )  ;
assign n2192 = in[7:0] ;
assign n2193 =  ( n2192 ) == ( bv_8_59_n603 )  ;
assign n2194 = in[7:0] ;
assign n2195 =  ( n2194 ) == ( bv_8_58_n346 )  ;
assign n2196 = in[7:0] ;
assign n2197 =  ( n2196 ) == ( bv_8_57_n558 )  ;
assign n2198 = in[7:0] ;
assign n2199 =  ( n2198 ) == ( bv_8_56_n481 )  ;
assign n2200 = in[7:0] ;
assign n2201 =  ( n2200 ) == ( bv_8_55_n292 )  ;
assign n2202 = in[7:0] ;
assign n2203 =  ( n2202 ) == ( bv_8_54_n650 )  ;
assign n2204 = in[7:0] ;
assign n2205 =  ( n2204 ) == ( bv_8_53_n152 )  ;
assign n2206 = in[7:0] ;
assign n2207 =  ( n2206 ) == ( bv_8_52_n656 )  ;
assign n2208 = in[7:0] ;
assign n2209 =  ( n2208 ) == ( bv_8_51_n528 )  ;
assign n2210 = in[7:0] ;
assign n2211 =  ( n2210 ) == ( bv_8_50_n349 )  ;
assign n2212 = in[7:0] ;
assign n2213 =  ( n2212 ) == ( bv_8_49_n665 )  ;
assign n2214 = in[7:0] ;
assign n2215 =  ( n2214 ) == ( bv_8_48_n668 )  ;
assign n2216 = in[7:0] ;
assign n2217 =  ( n2216 ) == ( bv_8_47_n591 )  ;
assign n2218 = in[7:0] ;
assign n2219 =  ( n2218 ) == ( bv_8_46_n235 )  ;
assign n2220 = in[7:0] ;
assign n2221 =  ( n2220 ) == ( bv_8_45_n26 )  ;
assign n2222 = in[7:0] ;
assign n2223 =  ( n2222 ) == ( bv_8_44_n621 )  ;
assign n2224 = in[7:0] ;
assign n2225 =  ( n2224 ) == ( bv_8_43_n681 )  ;
assign n2226 = in[7:0] ;
assign n2227 =  ( n2226 ) == ( bv_8_42_n387 )  ;
assign n2228 = in[7:0] ;
assign n2229 =  ( n2228 ) == ( bv_8_41_n596 )  ;
assign n2230 = in[7:0] ;
assign n2231 =  ( n2230 ) == ( bv_8_40_n74 )  ;
assign n2232 = in[7:0] ;
assign n2233 =  ( n2232 ) == ( bv_8_39_n634 )  ;
assign n2234 = in[7:0] ;
assign n2235 =  ( n2234 ) == ( bv_8_38_n692 )  ;
assign n2236 = in[7:0] ;
assign n2237 =  ( n2236 ) == ( bv_8_37_n239 )  ;
assign n2238 = in[7:0] ;
assign n2239 =  ( n2238 ) == ( bv_8_36_n330 )  ;
assign n2240 = in[7:0] ;
assign n2241 =  ( n2240 ) == ( bv_8_35_n663 )  ;
assign n2242 = in[7:0] ;
assign n2243 =  ( n2242 ) == ( bv_8_34_n390 )  ;
assign n2244 = in[7:0] ;
assign n2245 =  ( n2244 ) == ( bv_8_33_n468 )  ;
assign n2246 = in[7:0] ;
assign n2247 =  ( n2246 ) == ( bv_8_32_n575 )  ;
assign n2248 = in[7:0] ;
assign n2249 =  ( n2248 ) == ( bv_8_31_n206 )  ;
assign n2250 = in[7:0] ;
assign n2251 =  ( n2250 ) == ( bv_8_30_n93 )  ;
assign n2252 = in[7:0] ;
assign n2253 =  ( n2252 ) == ( bv_8_29_n133 )  ;
assign n2254 = in[7:0] ;
assign n2255 =  ( n2254 ) == ( bv_8_28_n231 )  ;
assign n2256 = in[7:0] ;
assign n2257 =  ( n2256 ) == ( bv_8_27_n615 )  ;
assign n2258 = in[7:0] ;
assign n2259 =  ( n2258 ) == ( bv_8_26_n618 )  ;
assign n2260 = in[7:0] ;
assign n2261 =  ( n2260 ) == ( bv_8_25_n410 )  ;
assign n2262 = in[7:0] ;
assign n2263 =  ( n2262 ) == ( bv_8_24_n658 )  ;
assign n2264 = in[7:0] ;
assign n2265 =  ( n2264 ) == ( bv_8_23_n429 )  ;
assign n2266 = in[7:0] ;
assign n2267 =  ( n2266 ) == ( bv_8_22_n6 )  ;
assign n2268 = in[7:0] ;
assign n2269 =  ( n2268 ) == ( bv_8_21_n673 )  ;
assign n2270 = in[7:0] ;
assign n2271 =  ( n2270 ) == ( bv_8_20_n368 )  ;
assign n2272 = in[7:0] ;
assign n2273 =  ( n2272 ) == ( bv_8_19_n446 )  ;
assign n2274 = in[7:0] ;
assign n2275 =  ( n2274 ) == ( bv_8_18_n643 )  ;
assign n2276 = in[7:0] ;
assign n2277 =  ( n2276 ) == ( bv_8_17_n116 )  ;
assign n2278 = in[7:0] ;
assign n2279 =  ( n2278 ) == ( bv_8_16_n464 )  ;
assign n2280 = in[7:0] ;
assign n2281 =  ( n2280 ) == ( bv_8_15_n22 )  ;
assign n2282 = in[7:0] ;
assign n2283 =  ( n2282 ) == ( bv_8_14_n160 )  ;
assign n2284 = in[7:0] ;
assign n2285 =  ( n2284 ) == ( bv_8_13_n54 )  ;
assign n2286 = in[7:0] ;
assign n2287 =  ( n2286 ) == ( bv_8_12_n449 )  ;
assign n2288 = in[7:0] ;
assign n2289 =  ( n2288 ) == ( bv_8_11_n358 )  ;
assign n2290 = in[7:0] ;
assign n2291 =  ( n2290 ) == ( bv_8_10_n342 )  ;
assign n2292 = in[7:0] ;
assign n2293 =  ( n2292 ) == ( bv_8_9_n626 )  ;
assign n2294 = in[7:0] ;
assign n2295 =  ( n2294 ) == ( bv_8_8_n249 )  ;
assign n2296 = in[7:0] ;
assign n2297 =  ( n2296 ) == ( bv_8_7_n646 )  ;
assign n2298 = in[7:0] ;
assign n2299 =  ( n2298 ) == ( bv_8_6_n334 )  ;
assign n2300 = in[7:0] ;
assign n2301 =  ( n2300 ) == ( bv_8_5_n652 )  ;
assign n2302 = in[7:0] ;
assign n2303 =  ( n2302 ) == ( bv_8_4_n670 )  ;
assign n2304 = in[7:0] ;
assign n2305 =  ( n2304 ) == ( bv_8_3_n167 )  ;
assign n2306 = in[7:0] ;
assign n2307 =  ( n2306 ) == ( bv_8_2_n517 )  ;
assign n2308 = in[7:0] ;
assign n2309 =  ( n2308 ) == ( bv_8_1_n752 )  ;
assign n2310 = in[7:0] ;
assign n2311 =  ( n2310 ) == ( bv_8_0_n582 )  ;
assign n2312 =  ( n2311 ) ? ( bv_8_99_n536 ) : ( bv_8_0_n582 ) ;
assign n2313 =  ( n2309 ) ? ( bv_8_124_n462 ) : ( n2312 ) ;
assign n2314 =  ( n2307 ) ? ( bv_8_119_n476 ) : ( n2313 ) ;
assign n2315 =  ( n2305 ) ? ( bv_8_123_n466 ) : ( n2314 ) ;
assign n2316 =  ( n2303 ) ? ( bv_8_242_n56 ) : ( n2315 ) ;
assign n2317 =  ( n2301 ) ? ( bv_8_107_n512 ) : ( n2316 ) ;
assign n2318 =  ( n2299 ) ? ( bv_8_111_n500 ) : ( n2317 ) ;
assign n2319 =  ( n2297 ) ? ( bv_8_197_n225 ) : ( n2318 ) ;
assign n2320 =  ( n2295 ) ? ( bv_8_48_n668 ) : ( n2319 ) ;
assign n2321 =  ( n2293 ) ? ( bv_8_1_n752 ) : ( n2320 ) ;
assign n2322 =  ( n2291 ) ? ( bv_8_103_n524 ) : ( n2321 ) ;
assign n2323 =  ( n2289 ) ? ( bv_8_43_n681 ) : ( n2322 ) ;
assign n2324 =  ( n2287 ) ? ( bv_8_254_n8 ) : ( n2323 ) ;
assign n2325 =  ( n2285 ) ? ( bv_8_215_n158 ) : ( n2324 ) ;
assign n2326 =  ( n2283 ) ? ( bv_8_171_n313 ) : ( n2325 ) ;
assign n2327 =  ( n2281 ) ? ( bv_8_118_n479 ) : ( n2326 ) ;
assign n2328 =  ( n2279 ) ? ( bv_8_202_n208 ) : ( n2327 ) ;
assign n2329 =  ( n2277 ) ? ( bv_8_130_n444 ) : ( n2328 ) ;
assign n2330 =  ( n2275 ) ? ( bv_8_201_n212 ) : ( n2329 ) ;
assign n2331 =  ( n2273 ) ? ( bv_8_125_n459 ) : ( n2330 ) ;
assign n2332 =  ( n2271 ) ? ( bv_8_250_n24 ) : ( n2331 ) ;
assign n2333 =  ( n2269 ) ? ( bv_8_89_n563 ) : ( n2332 ) ;
assign n2334 =  ( n2267 ) ? ( bv_8_71_n607 ) : ( n2333 ) ;
assign n2335 =  ( n2265 ) ? ( bv_8_240_n64 ) : ( n2334 ) ;
assign n2336 =  ( n2263 ) ? ( bv_8_173_n305 ) : ( n2335 ) ;
assign n2337 =  ( n2261 ) ? ( bv_8_212_n169 ) : ( n2336 ) ;
assign n2338 =  ( n2259 ) ? ( bv_8_162_n344 ) : ( n2337 ) ;
assign n2339 =  ( n2257 ) ? ( bv_8_175_n299 ) : ( n2338 ) ;
assign n2340 =  ( n2255 ) ? ( bv_8_156_n364 ) : ( n2339 ) ;
assign n2341 =  ( n2253 ) ? ( bv_8_164_n336 ) : ( n2340 ) ;
assign n2342 =  ( n2251 ) ? ( bv_8_114_n490 ) : ( n2341 ) ;
assign n2343 =  ( n2249 ) ? ( bv_8_192_n244 ) : ( n2342 ) ;
assign n2344 =  ( n2247 ) ? ( bv_8_183_n273 ) : ( n2343 ) ;
assign n2345 =  ( n2245 ) ? ( bv_8_253_n12 ) : ( n2344 ) ;
assign n2346 =  ( n2243 ) ? ( bv_8_147_n392 ) : ( n2345 ) ;
assign n2347 =  ( n2241 ) ? ( bv_8_38_n692 ) : ( n2346 ) ;
assign n2348 =  ( n2239 ) ? ( bv_8_54_n650 ) : ( n2347 ) ;
assign n2349 =  ( n2237 ) ? ( bv_8_63_n628 ) : ( n2348 ) ;
assign n2350 =  ( n2235 ) ? ( bv_8_247_n36 ) : ( n2349 ) ;
assign n2351 =  ( n2233 ) ? ( bv_8_204_n200 ) : ( n2350 ) ;
assign n2352 =  ( n2231 ) ? ( bv_8_52_n656 ) : ( n2351 ) ;
assign n2353 =  ( n2229 ) ? ( bv_8_165_n332 ) : ( n2352 ) ;
assign n2354 =  ( n2227 ) ? ( bv_8_229_n106 ) : ( n2353 ) ;
assign n2355 =  ( n2225 ) ? ( bv_8_241_n60 ) : ( n2354 ) ;
assign n2356 =  ( n2223 ) ? ( bv_8_113_n494 ) : ( n2355 ) ;
assign n2357 =  ( n2221 ) ? ( bv_8_216_n154 ) : ( n2356 ) ;
assign n2358 =  ( n2219 ) ? ( bv_8_49_n665 ) : ( n2357 ) ;
assign n2359 =  ( n2217 ) ? ( bv_8_21_n673 ) : ( n2358 ) ;
assign n2360 =  ( n2215 ) ? ( bv_8_4_n670 ) : ( n2359 ) ;
assign n2361 =  ( n2213 ) ? ( bv_8_199_n218 ) : ( n2360 ) ;
assign n2362 =  ( n2211 ) ? ( bv_8_35_n663 ) : ( n2361 ) ;
assign n2363 =  ( n2209 ) ? ( bv_8_195_n233 ) : ( n2362 ) ;
assign n2364 =  ( n2207 ) ? ( bv_8_24_n658 ) : ( n2363 ) ;
assign n2365 =  ( n2205 ) ? ( bv_8_150_n382 ) : ( n2364 ) ;
assign n2366 =  ( n2203 ) ? ( bv_8_5_n652 ) : ( n2365 ) ;
assign n2367 =  ( n2201 ) ? ( bv_8_154_n370 ) : ( n2366 ) ;
assign n2368 =  ( n2199 ) ? ( bv_8_7_n646 ) : ( n2367 ) ;
assign n2369 =  ( n2197 ) ? ( bv_8_18_n643 ) : ( n2368 ) ;
assign n2370 =  ( n2195 ) ? ( bv_8_128_n451 ) : ( n2369 ) ;
assign n2371 =  ( n2193 ) ? ( bv_8_226_n118 ) : ( n2370 ) ;
assign n2372 =  ( n2191 ) ? ( bv_8_235_n84 ) : ( n2371 ) ;
assign n2373 =  ( n2189 ) ? ( bv_8_39_n634 ) : ( n2372 ) ;
assign n2374 =  ( n2187 ) ? ( bv_8_178_n290 ) : ( n2373 ) ;
assign n2375 =  ( n2185 ) ? ( bv_8_117_n483 ) : ( n2374 ) ;
assign n2376 =  ( n2183 ) ? ( bv_8_9_n626 ) : ( n2375 ) ;
assign n2377 =  ( n2181 ) ? ( bv_8_131_n441 ) : ( n2376 ) ;
assign n2378 =  ( n2179 ) ? ( bv_8_44_n621 ) : ( n2377 ) ;
assign n2379 =  ( n2177 ) ? ( bv_8_26_n618 ) : ( n2378 ) ;
assign n2380 =  ( n2175 ) ? ( bv_8_27_n615 ) : ( n2379 ) ;
assign n2381 =  ( n2173 ) ? ( bv_8_110_n503 ) : ( n2380 ) ;
assign n2382 =  ( n2171 ) ? ( bv_8_90_n560 ) : ( n2381 ) ;
assign n2383 =  ( n2169 ) ? ( bv_8_160_n351 ) : ( n2382 ) ;
assign n2384 =  ( n2167 ) ? ( bv_8_82_n580 ) : ( n2383 ) ;
assign n2385 =  ( n2165 ) ? ( bv_8_59_n603 ) : ( n2384 ) ;
assign n2386 =  ( n2163 ) ? ( bv_8_214_n162 ) : ( n2385 ) ;
assign n2387 =  ( n2161 ) ? ( bv_8_179_n286 ) : ( n2386 ) ;
assign n2388 =  ( n2159 ) ? ( bv_8_41_n596 ) : ( n2387 ) ;
assign n2389 =  ( n2157 ) ? ( bv_8_227_n114 ) : ( n2388 ) ;
assign n2390 =  ( n2155 ) ? ( bv_8_47_n591 ) : ( n2389 ) ;
assign n2391 =  ( n2153 ) ? ( bv_8_132_n437 ) : ( n2390 ) ;
assign n2392 =  ( n2151 ) ? ( bv_8_83_n577 ) : ( n2391 ) ;
assign n2393 =  ( n2149 ) ? ( bv_8_209_n181 ) : ( n2392 ) ;
assign n2394 =  ( n2147 ) ? ( bv_8_0_n582 ) : ( n2393 ) ;
assign n2395 =  ( n2145 ) ? ( bv_8_237_n76 ) : ( n2394 ) ;
assign n2396 =  ( n2143 ) ? ( bv_8_32_n575 ) : ( n2395 ) ;
assign n2397 =  ( n2141 ) ? ( bv_8_252_n16 ) : ( n2396 ) ;
assign n2398 =  ( n2139 ) ? ( bv_8_177_n294 ) : ( n2397 ) ;
assign n2399 =  ( n2137 ) ? ( bv_8_91_n556 ) : ( n2398 ) ;
assign n2400 =  ( n2135 ) ? ( bv_8_106_n515 ) : ( n2399 ) ;
assign n2401 =  ( n2133 ) ? ( bv_8_203_n204 ) : ( n2400 ) ;
assign n2402 =  ( n2131 ) ? ( bv_8_190_n251 ) : ( n2401 ) ;
assign n2403 =  ( n2129 ) ? ( bv_8_57_n558 ) : ( n2402 ) ;
assign n2404 =  ( n2127 ) ? ( bv_8_74_n554 ) : ( n2403 ) ;
assign n2405 =  ( n2125 ) ? ( bv_8_76_n551 ) : ( n2404 ) ;
assign n2406 =  ( n2123 ) ? ( bv_8_88_n548 ) : ( n2405 ) ;
assign n2407 =  ( n2121 ) ? ( bv_8_207_n189 ) : ( n2406 ) ;
assign n2408 =  ( n2119 ) ? ( bv_8_208_n185 ) : ( n2407 ) ;
assign n2409 =  ( n2117 ) ? ( bv_8_239_n68 ) : ( n2408 ) ;
assign n2410 =  ( n2115 ) ? ( bv_8_170_n317 ) : ( n2409 ) ;
assign n2411 =  ( n2113 ) ? ( bv_8_251_n20 ) : ( n2410 ) ;
assign n2412 =  ( n2111 ) ? ( bv_8_67_n534 ) : ( n2411 ) ;
assign n2413 =  ( n2109 ) ? ( bv_8_77_n531 ) : ( n2412 ) ;
assign n2414 =  ( n2107 ) ? ( bv_8_51_n528 ) : ( n2413 ) ;
assign n2415 =  ( n2105 ) ? ( bv_8_133_n434 ) : ( n2414 ) ;
assign n2416 =  ( n2103 ) ? ( bv_8_69_n522 ) : ( n2415 ) ;
assign n2417 =  ( n2101 ) ? ( bv_8_249_n28 ) : ( n2416 ) ;
assign n2418 =  ( n2099 ) ? ( bv_8_2_n517 ) : ( n2417 ) ;
assign n2419 =  ( n2097 ) ? ( bv_8_127_n454 ) : ( n2418 ) ;
assign n2420 =  ( n2095 ) ? ( bv_8_80_n510 ) : ( n2419 ) ;
assign n2421 =  ( n2093 ) ? ( bv_8_60_n507 ) : ( n2420 ) ;
assign n2422 =  ( n2091 ) ? ( bv_8_159_n354 ) : ( n2421 ) ;
assign n2423 =  ( n2089 ) ? ( bv_8_168_n322 ) : ( n2422 ) ;
assign n2424 =  ( n2087 ) ? ( bv_8_81_n498 ) : ( n2423 ) ;
assign n2425 =  ( n2085 ) ? ( bv_8_163_n340 ) : ( n2424 ) ;
assign n2426 =  ( n2083 ) ? ( bv_8_64_n492 ) : ( n2425 ) ;
assign n2427 =  ( n2081 ) ? ( bv_8_143_n405 ) : ( n2426 ) ;
assign n2428 =  ( n2079 ) ? ( bv_8_146_n395 ) : ( n2427 ) ;
assign n2429 =  ( n2077 ) ? ( bv_8_157_n360 ) : ( n2428 ) ;
assign n2430 =  ( n2075 ) ? ( bv_8_56_n481 ) : ( n2429 ) ;
assign n2431 =  ( n2073 ) ? ( bv_8_245_n44 ) : ( n2430 ) ;
assign n2432 =  ( n2071 ) ? ( bv_8_188_n258 ) : ( n2431 ) ;
assign n2433 =  ( n2069 ) ? ( bv_8_182_n277 ) : ( n2432 ) ;
assign n2434 =  ( n2067 ) ? ( bv_8_218_n147 ) : ( n2433 ) ;
assign n2435 =  ( n2065 ) ? ( bv_8_33_n468 ) : ( n2434 ) ;
assign n2436 =  ( n2063 ) ? ( bv_8_16_n464 ) : ( n2435 ) ;
assign n2437 =  ( n2061 ) ? ( bv_8_255_n4 ) : ( n2436 ) ;
assign n2438 =  ( n2059 ) ? ( bv_8_243_n52 ) : ( n2437 ) ;
assign n2439 =  ( n2057 ) ? ( bv_8_210_n177 ) : ( n2438 ) ;
assign n2440 =  ( n2055 ) ? ( bv_8_205_n196 ) : ( n2439 ) ;
assign n2441 =  ( n2053 ) ? ( bv_8_12_n449 ) : ( n2440 ) ;
assign n2442 =  ( n2051 ) ? ( bv_8_19_n446 ) : ( n2441 ) ;
assign n2443 =  ( n2049 ) ? ( bv_8_236_n80 ) : ( n2442 ) ;
assign n2444 =  ( n2047 ) ? ( bv_8_95_n439 ) : ( n2443 ) ;
assign n2445 =  ( n2045 ) ? ( bv_8_151_n378 ) : ( n2444 ) ;
assign n2446 =  ( n2043 ) ? ( bv_8_68_n432 ) : ( n2445 ) ;
assign n2447 =  ( n2041 ) ? ( bv_8_23_n429 ) : ( n2446 ) ;
assign n2448 =  ( n2039 ) ? ( bv_8_196_n229 ) : ( n2447 ) ;
assign n2449 =  ( n2037 ) ? ( bv_8_167_n325 ) : ( n2448 ) ;
assign n2450 =  ( n2035 ) ? ( bv_8_126_n422 ) : ( n2449 ) ;
assign n2451 =  ( n2033 ) ? ( bv_8_61_n419 ) : ( n2450 ) ;
assign n2452 =  ( n2031 ) ? ( bv_8_100_n416 ) : ( n2451 ) ;
assign n2453 =  ( n2029 ) ? ( bv_8_93_n413 ) : ( n2452 ) ;
assign n2454 =  ( n2027 ) ? ( bv_8_25_n410 ) : ( n2453 ) ;
assign n2455 =  ( n2025 ) ? ( bv_8_115_n407 ) : ( n2454 ) ;
assign n2456 =  ( n2023 ) ? ( bv_8_96_n403 ) : ( n2455 ) ;
assign n2457 =  ( n2021 ) ? ( bv_8_129_n400 ) : ( n2456 ) ;
assign n2458 =  ( n2019 ) ? ( bv_8_79_n397 ) : ( n2457 ) ;
assign n2459 =  ( n2017 ) ? ( bv_8_220_n139 ) : ( n2458 ) ;
assign n2460 =  ( n2015 ) ? ( bv_8_34_n390 ) : ( n2459 ) ;
assign n2461 =  ( n2013 ) ? ( bv_8_42_n387 ) : ( n2460 ) ;
assign n2462 =  ( n2011 ) ? ( bv_8_144_n384 ) : ( n2461 ) ;
assign n2463 =  ( n2009 ) ? ( bv_8_136_n380 ) : ( n2462 ) ;
assign n2464 =  ( n2007 ) ? ( bv_8_70_n376 ) : ( n2463 ) ;
assign n2465 =  ( n2005 ) ? ( bv_8_238_n72 ) : ( n2464 ) ;
assign n2466 =  ( n2003 ) ? ( bv_8_184_n269 ) : ( n2465 ) ;
assign n2467 =  ( n2001 ) ? ( bv_8_20_n368 ) : ( n2466 ) ;
assign n2468 =  ( n1999 ) ? ( bv_8_222_n131 ) : ( n2467 ) ;
assign n2469 =  ( n1997 ) ? ( bv_8_94_n362 ) : ( n2468 ) ;
assign n2470 =  ( n1995 ) ? ( bv_8_11_n358 ) : ( n2469 ) ;
assign n2471 =  ( n1993 ) ? ( bv_8_219_n143 ) : ( n2470 ) ;
assign n2472 =  ( n1991 ) ? ( bv_8_224_n125 ) : ( n2471 ) ;
assign n2473 =  ( n1989 ) ? ( bv_8_50_n349 ) : ( n2472 ) ;
assign n2474 =  ( n1987 ) ? ( bv_8_58_n346 ) : ( n2473 ) ;
assign n2475 =  ( n1985 ) ? ( bv_8_10_n342 ) : ( n2474 ) ;
assign n2476 =  ( n1983 ) ? ( bv_8_73_n338 ) : ( n2475 ) ;
assign n2477 =  ( n1981 ) ? ( bv_8_6_n334 ) : ( n2476 ) ;
assign n2478 =  ( n1979 ) ? ( bv_8_36_n330 ) : ( n2477 ) ;
assign n2479 =  ( n1977 ) ? ( bv_8_92_n327 ) : ( n2478 ) ;
assign n2480 =  ( n1975 ) ? ( bv_8_194_n237 ) : ( n2479 ) ;
assign n2481 =  ( n1973 ) ? ( bv_8_211_n173 ) : ( n2480 ) ;
assign n2482 =  ( n1971 ) ? ( bv_8_172_n309 ) : ( n2481 ) ;
assign n2483 =  ( n1969 ) ? ( bv_8_98_n315 ) : ( n2482 ) ;
assign n2484 =  ( n1967 ) ? ( bv_8_145_n311 ) : ( n2483 ) ;
assign n2485 =  ( n1965 ) ? ( bv_8_149_n307 ) : ( n2484 ) ;
assign n2486 =  ( n1963 ) ? ( bv_8_228_n110 ) : ( n2485 ) ;
assign n2487 =  ( n1961 ) ? ( bv_8_121_n301 ) : ( n2486 ) ;
assign n2488 =  ( n1959 ) ? ( bv_8_231_n99 ) : ( n2487 ) ;
assign n2489 =  ( n1957 ) ? ( bv_8_200_n215 ) : ( n2488 ) ;
assign n2490 =  ( n1955 ) ? ( bv_8_55_n292 ) : ( n2489 ) ;
assign n2491 =  ( n1953 ) ? ( bv_8_109_n288 ) : ( n2490 ) ;
assign n2492 =  ( n1951 ) ? ( bv_8_141_n284 ) : ( n2491 ) ;
assign n2493 =  ( n1949 ) ? ( bv_8_213_n165 ) : ( n2492 ) ;
assign n2494 =  ( n1947 ) ? ( bv_8_78_n279 ) : ( n2493 ) ;
assign n2495 =  ( n1945 ) ? ( bv_8_169_n275 ) : ( n2494 ) ;
assign n2496 =  ( n1943 ) ? ( bv_8_108_n271 ) : ( n2495 ) ;
assign n2497 =  ( n1941 ) ? ( bv_8_86_n267 ) : ( n2496 ) ;
assign n2498 =  ( n1939 ) ? ( bv_8_244_n48 ) : ( n2497 ) ;
assign n2499 =  ( n1937 ) ? ( bv_8_234_n88 ) : ( n2498 ) ;
assign n2500 =  ( n1935 ) ? ( bv_8_101_n260 ) : ( n2499 ) ;
assign n2501 =  ( n1933 ) ? ( bv_8_122_n256 ) : ( n2500 ) ;
assign n2502 =  ( n1931 ) ? ( bv_8_174_n253 ) : ( n2501 ) ;
assign n2503 =  ( n1929 ) ? ( bv_8_8_n249 ) : ( n2502 ) ;
assign n2504 =  ( n1927 ) ? ( bv_8_186_n246 ) : ( n2503 ) ;
assign n2505 =  ( n1925 ) ? ( bv_8_120_n242 ) : ( n2504 ) ;
assign n2506 =  ( n1923 ) ? ( bv_8_37_n239 ) : ( n2505 ) ;
assign n2507 =  ( n1921 ) ? ( bv_8_46_n235 ) : ( n2506 ) ;
assign n2508 =  ( n1919 ) ? ( bv_8_28_n231 ) : ( n2507 ) ;
assign n2509 =  ( n1917 ) ? ( bv_8_166_n227 ) : ( n2508 ) ;
assign n2510 =  ( n1915 ) ? ( bv_8_180_n223 ) : ( n2509 ) ;
assign n2511 =  ( n1913 ) ? ( bv_8_198_n220 ) : ( n2510 ) ;
assign n2512 =  ( n1911 ) ? ( bv_8_232_n95 ) : ( n2511 ) ;
assign n2513 =  ( n1909 ) ? ( bv_8_221_n135 ) : ( n2512 ) ;
assign n2514 =  ( n1907 ) ? ( bv_8_116_n210 ) : ( n2513 ) ;
assign n2515 =  ( n1905 ) ? ( bv_8_31_n206 ) : ( n2514 ) ;
assign n2516 =  ( n1903 ) ? ( bv_8_75_n202 ) : ( n2515 ) ;
assign n2517 =  ( n1901 ) ? ( bv_8_189_n198 ) : ( n2516 ) ;
assign n2518 =  ( n1899 ) ? ( bv_8_139_n194 ) : ( n2517 ) ;
assign n2519 =  ( n1897 ) ? ( bv_8_138_n191 ) : ( n2518 ) ;
assign n2520 =  ( n1895 ) ? ( bv_8_112_n187 ) : ( n2519 ) ;
assign n2521 =  ( n1893 ) ? ( bv_8_62_n183 ) : ( n2520 ) ;
assign n2522 =  ( n1891 ) ? ( bv_8_181_n179 ) : ( n2521 ) ;
assign n2523 =  ( n1889 ) ? ( bv_8_102_n175 ) : ( n2522 ) ;
assign n2524 =  ( n1887 ) ? ( bv_8_72_n171 ) : ( n2523 ) ;
assign n2525 =  ( n1885 ) ? ( bv_8_3_n167 ) : ( n2524 ) ;
assign n2526 =  ( n1883 ) ? ( bv_8_246_n40 ) : ( n2525 ) ;
assign n2527 =  ( n1881 ) ? ( bv_8_14_n160 ) : ( n2526 ) ;
assign n2528 =  ( n1879 ) ? ( bv_8_97_n156 ) : ( n2527 ) ;
assign n2529 =  ( n1877 ) ? ( bv_8_53_n152 ) : ( n2528 ) ;
assign n2530 =  ( n1875 ) ? ( bv_8_87_n149 ) : ( n2529 ) ;
assign n2531 =  ( n1873 ) ? ( bv_8_185_n145 ) : ( n2530 ) ;
assign n2532 =  ( n1871 ) ? ( bv_8_134_n141 ) : ( n2531 ) ;
assign n2533 =  ( n1869 ) ? ( bv_8_193_n137 ) : ( n2532 ) ;
assign n2534 =  ( n1867 ) ? ( bv_8_29_n133 ) : ( n2533 ) ;
assign n2535 =  ( n1865 ) ? ( bv_8_158_n129 ) : ( n2534 ) ;
assign n2536 =  ( n1863 ) ? ( bv_8_225_n122 ) : ( n2535 ) ;
assign n2537 =  ( n1861 ) ? ( bv_8_248_n32 ) : ( n2536 ) ;
assign n2538 =  ( n1859 ) ? ( bv_8_152_n120 ) : ( n2537 ) ;
assign n2539 =  ( n1857 ) ? ( bv_8_17_n116 ) : ( n2538 ) ;
assign n2540 =  ( n1855 ) ? ( bv_8_105_n112 ) : ( n2539 ) ;
assign n2541 =  ( n1853 ) ? ( bv_8_217_n108 ) : ( n2540 ) ;
assign n2542 =  ( n1851 ) ? ( bv_8_142_n104 ) : ( n2541 ) ;
assign n2543 =  ( n1849 ) ? ( bv_8_148_n101 ) : ( n2542 ) ;
assign n2544 =  ( n1847 ) ? ( bv_8_155_n97 ) : ( n2543 ) ;
assign n2545 =  ( n1845 ) ? ( bv_8_30_n93 ) : ( n2544 ) ;
assign n2546 =  ( n1843 ) ? ( bv_8_135_n90 ) : ( n2545 ) ;
assign n2547 =  ( n1841 ) ? ( bv_8_233_n86 ) : ( n2546 ) ;
assign n2548 =  ( n1839 ) ? ( bv_8_206_n82 ) : ( n2547 ) ;
assign n2549 =  ( n1837 ) ? ( bv_8_85_n78 ) : ( n2548 ) ;
assign n2550 =  ( n1835 ) ? ( bv_8_40_n74 ) : ( n2549 ) ;
assign n2551 =  ( n1833 ) ? ( bv_8_223_n70 ) : ( n2550 ) ;
assign n2552 =  ( n1831 ) ? ( bv_8_140_n66 ) : ( n2551 ) ;
assign n2553 =  ( n1829 ) ? ( bv_8_161_n62 ) : ( n2552 ) ;
assign n2554 =  ( n1827 ) ? ( bv_8_137_n58 ) : ( n2553 ) ;
assign n2555 =  ( n1825 ) ? ( bv_8_13_n54 ) : ( n2554 ) ;
assign n2556 =  ( n1823 ) ? ( bv_8_191_n50 ) : ( n2555 ) ;
assign n2557 =  ( n1821 ) ? ( bv_8_230_n46 ) : ( n2556 ) ;
assign n2558 =  ( n1819 ) ? ( bv_8_66_n42 ) : ( n2557 ) ;
assign n2559 =  ( n1817 ) ? ( bv_8_104_n38 ) : ( n2558 ) ;
assign n2560 =  ( n1815 ) ? ( bv_8_65_n34 ) : ( n2559 ) ;
assign n2561 =  ( n1813 ) ? ( bv_8_153_n30 ) : ( n2560 ) ;
assign n2562 =  ( n1811 ) ? ( bv_8_45_n26 ) : ( n2561 ) ;
assign n2563 =  ( n1809 ) ? ( bv_8_15_n22 ) : ( n2562 ) ;
assign n2564 =  ( n1807 ) ? ( bv_8_176_n18 ) : ( n2563 ) ;
assign n2565 =  ( n1805 ) ? ( bv_8_84_n14 ) : ( n2564 ) ;
assign n2566 =  ( n1803 ) ? ( bv_8_187_n10 ) : ( n2565 ) ;
assign n2567 =  ( n1801 ) ? ( bv_8_22_n6 ) : ( n2566 ) ;
assign n2568 =  ( n1799 ) ^ ( n2567 )  ;
assign n2569 =  { ( n1798 ) , ( n2568 ) }  ;
assign n2570 = in[103:96] ;
assign n2571 = in[31:24] ;
assign n2572 =  ( n2571 ) == ( bv_8_255_n4 )  ;
assign n2573 = in[31:24] ;
assign n2574 =  ( n2573 ) == ( bv_8_254_n8 )  ;
assign n2575 = in[31:24] ;
assign n2576 =  ( n2575 ) == ( bv_8_253_n12 )  ;
assign n2577 = in[31:24] ;
assign n2578 =  ( n2577 ) == ( bv_8_252_n16 )  ;
assign n2579 = in[31:24] ;
assign n2580 =  ( n2579 ) == ( bv_8_251_n20 )  ;
assign n2581 = in[31:24] ;
assign n2582 =  ( n2581 ) == ( bv_8_250_n24 )  ;
assign n2583 = in[31:24] ;
assign n2584 =  ( n2583 ) == ( bv_8_249_n28 )  ;
assign n2585 = in[31:24] ;
assign n2586 =  ( n2585 ) == ( bv_8_248_n32 )  ;
assign n2587 = in[31:24] ;
assign n2588 =  ( n2587 ) == ( bv_8_247_n36 )  ;
assign n2589 = in[31:24] ;
assign n2590 =  ( n2589 ) == ( bv_8_246_n40 )  ;
assign n2591 = in[31:24] ;
assign n2592 =  ( n2591 ) == ( bv_8_245_n44 )  ;
assign n2593 = in[31:24] ;
assign n2594 =  ( n2593 ) == ( bv_8_244_n48 )  ;
assign n2595 = in[31:24] ;
assign n2596 =  ( n2595 ) == ( bv_8_243_n52 )  ;
assign n2597 = in[31:24] ;
assign n2598 =  ( n2597 ) == ( bv_8_242_n56 )  ;
assign n2599 = in[31:24] ;
assign n2600 =  ( n2599 ) == ( bv_8_241_n60 )  ;
assign n2601 = in[31:24] ;
assign n2602 =  ( n2601 ) == ( bv_8_240_n64 )  ;
assign n2603 = in[31:24] ;
assign n2604 =  ( n2603 ) == ( bv_8_239_n68 )  ;
assign n2605 = in[31:24] ;
assign n2606 =  ( n2605 ) == ( bv_8_238_n72 )  ;
assign n2607 = in[31:24] ;
assign n2608 =  ( n2607 ) == ( bv_8_237_n76 )  ;
assign n2609 = in[31:24] ;
assign n2610 =  ( n2609 ) == ( bv_8_236_n80 )  ;
assign n2611 = in[31:24] ;
assign n2612 =  ( n2611 ) == ( bv_8_235_n84 )  ;
assign n2613 = in[31:24] ;
assign n2614 =  ( n2613 ) == ( bv_8_234_n88 )  ;
assign n2615 = in[31:24] ;
assign n2616 =  ( n2615 ) == ( bv_8_233_n86 )  ;
assign n2617 = in[31:24] ;
assign n2618 =  ( n2617 ) == ( bv_8_232_n95 )  ;
assign n2619 = in[31:24] ;
assign n2620 =  ( n2619 ) == ( bv_8_231_n99 )  ;
assign n2621 = in[31:24] ;
assign n2622 =  ( n2621 ) == ( bv_8_230_n46 )  ;
assign n2623 = in[31:24] ;
assign n2624 =  ( n2623 ) == ( bv_8_229_n106 )  ;
assign n2625 = in[31:24] ;
assign n2626 =  ( n2625 ) == ( bv_8_228_n110 )  ;
assign n2627 = in[31:24] ;
assign n2628 =  ( n2627 ) == ( bv_8_227_n114 )  ;
assign n2629 = in[31:24] ;
assign n2630 =  ( n2629 ) == ( bv_8_226_n118 )  ;
assign n2631 = in[31:24] ;
assign n2632 =  ( n2631 ) == ( bv_8_225_n122 )  ;
assign n2633 = in[31:24] ;
assign n2634 =  ( n2633 ) == ( bv_8_224_n125 )  ;
assign n2635 = in[31:24] ;
assign n2636 =  ( n2635 ) == ( bv_8_223_n70 )  ;
assign n2637 = in[31:24] ;
assign n2638 =  ( n2637 ) == ( bv_8_222_n131 )  ;
assign n2639 = in[31:24] ;
assign n2640 =  ( n2639 ) == ( bv_8_221_n135 )  ;
assign n2641 = in[31:24] ;
assign n2642 =  ( n2641 ) == ( bv_8_220_n139 )  ;
assign n2643 = in[31:24] ;
assign n2644 =  ( n2643 ) == ( bv_8_219_n143 )  ;
assign n2645 = in[31:24] ;
assign n2646 =  ( n2645 ) == ( bv_8_218_n147 )  ;
assign n2647 = in[31:24] ;
assign n2648 =  ( n2647 ) == ( bv_8_217_n108 )  ;
assign n2649 = in[31:24] ;
assign n2650 =  ( n2649 ) == ( bv_8_216_n154 )  ;
assign n2651 = in[31:24] ;
assign n2652 =  ( n2651 ) == ( bv_8_215_n158 )  ;
assign n2653 = in[31:24] ;
assign n2654 =  ( n2653 ) == ( bv_8_214_n162 )  ;
assign n2655 = in[31:24] ;
assign n2656 =  ( n2655 ) == ( bv_8_213_n165 )  ;
assign n2657 = in[31:24] ;
assign n2658 =  ( n2657 ) == ( bv_8_212_n169 )  ;
assign n2659 = in[31:24] ;
assign n2660 =  ( n2659 ) == ( bv_8_211_n173 )  ;
assign n2661 = in[31:24] ;
assign n2662 =  ( n2661 ) == ( bv_8_210_n177 )  ;
assign n2663 = in[31:24] ;
assign n2664 =  ( n2663 ) == ( bv_8_209_n181 )  ;
assign n2665 = in[31:24] ;
assign n2666 =  ( n2665 ) == ( bv_8_208_n185 )  ;
assign n2667 = in[31:24] ;
assign n2668 =  ( n2667 ) == ( bv_8_207_n189 )  ;
assign n2669 = in[31:24] ;
assign n2670 =  ( n2669 ) == ( bv_8_206_n82 )  ;
assign n2671 = in[31:24] ;
assign n2672 =  ( n2671 ) == ( bv_8_205_n196 )  ;
assign n2673 = in[31:24] ;
assign n2674 =  ( n2673 ) == ( bv_8_204_n200 )  ;
assign n2675 = in[31:24] ;
assign n2676 =  ( n2675 ) == ( bv_8_203_n204 )  ;
assign n2677 = in[31:24] ;
assign n2678 =  ( n2677 ) == ( bv_8_202_n208 )  ;
assign n2679 = in[31:24] ;
assign n2680 =  ( n2679 ) == ( bv_8_201_n212 )  ;
assign n2681 = in[31:24] ;
assign n2682 =  ( n2681 ) == ( bv_8_200_n215 )  ;
assign n2683 = in[31:24] ;
assign n2684 =  ( n2683 ) == ( bv_8_199_n218 )  ;
assign n2685 = in[31:24] ;
assign n2686 =  ( n2685 ) == ( bv_8_198_n220 )  ;
assign n2687 = in[31:24] ;
assign n2688 =  ( n2687 ) == ( bv_8_197_n225 )  ;
assign n2689 = in[31:24] ;
assign n2690 =  ( n2689 ) == ( bv_8_196_n229 )  ;
assign n2691 = in[31:24] ;
assign n2692 =  ( n2691 ) == ( bv_8_195_n233 )  ;
assign n2693 = in[31:24] ;
assign n2694 =  ( n2693 ) == ( bv_8_194_n237 )  ;
assign n2695 = in[31:24] ;
assign n2696 =  ( n2695 ) == ( bv_8_193_n137 )  ;
assign n2697 = in[31:24] ;
assign n2698 =  ( n2697 ) == ( bv_8_192_n244 )  ;
assign n2699 = in[31:24] ;
assign n2700 =  ( n2699 ) == ( bv_8_191_n50 )  ;
assign n2701 = in[31:24] ;
assign n2702 =  ( n2701 ) == ( bv_8_190_n251 )  ;
assign n2703 = in[31:24] ;
assign n2704 =  ( n2703 ) == ( bv_8_189_n198 )  ;
assign n2705 = in[31:24] ;
assign n2706 =  ( n2705 ) == ( bv_8_188_n258 )  ;
assign n2707 = in[31:24] ;
assign n2708 =  ( n2707 ) == ( bv_8_187_n10 )  ;
assign n2709 = in[31:24] ;
assign n2710 =  ( n2709 ) == ( bv_8_186_n246 )  ;
assign n2711 = in[31:24] ;
assign n2712 =  ( n2711 ) == ( bv_8_185_n145 )  ;
assign n2713 = in[31:24] ;
assign n2714 =  ( n2713 ) == ( bv_8_184_n269 )  ;
assign n2715 = in[31:24] ;
assign n2716 =  ( n2715 ) == ( bv_8_183_n273 )  ;
assign n2717 = in[31:24] ;
assign n2718 =  ( n2717 ) == ( bv_8_182_n277 )  ;
assign n2719 = in[31:24] ;
assign n2720 =  ( n2719 ) == ( bv_8_181_n179 )  ;
assign n2721 = in[31:24] ;
assign n2722 =  ( n2721 ) == ( bv_8_180_n223 )  ;
assign n2723 = in[31:24] ;
assign n2724 =  ( n2723 ) == ( bv_8_179_n286 )  ;
assign n2725 = in[31:24] ;
assign n2726 =  ( n2725 ) == ( bv_8_178_n290 )  ;
assign n2727 = in[31:24] ;
assign n2728 =  ( n2727 ) == ( bv_8_177_n294 )  ;
assign n2729 = in[31:24] ;
assign n2730 =  ( n2729 ) == ( bv_8_176_n18 )  ;
assign n2731 = in[31:24] ;
assign n2732 =  ( n2731 ) == ( bv_8_175_n299 )  ;
assign n2733 = in[31:24] ;
assign n2734 =  ( n2733 ) == ( bv_8_174_n253 )  ;
assign n2735 = in[31:24] ;
assign n2736 =  ( n2735 ) == ( bv_8_173_n305 )  ;
assign n2737 = in[31:24] ;
assign n2738 =  ( n2737 ) == ( bv_8_172_n309 )  ;
assign n2739 = in[31:24] ;
assign n2740 =  ( n2739 ) == ( bv_8_171_n313 )  ;
assign n2741 = in[31:24] ;
assign n2742 =  ( n2741 ) == ( bv_8_170_n317 )  ;
assign n2743 = in[31:24] ;
assign n2744 =  ( n2743 ) == ( bv_8_169_n275 )  ;
assign n2745 = in[31:24] ;
assign n2746 =  ( n2745 ) == ( bv_8_168_n322 )  ;
assign n2747 = in[31:24] ;
assign n2748 =  ( n2747 ) == ( bv_8_167_n325 )  ;
assign n2749 = in[31:24] ;
assign n2750 =  ( n2749 ) == ( bv_8_166_n227 )  ;
assign n2751 = in[31:24] ;
assign n2752 =  ( n2751 ) == ( bv_8_165_n332 )  ;
assign n2753 = in[31:24] ;
assign n2754 =  ( n2753 ) == ( bv_8_164_n336 )  ;
assign n2755 = in[31:24] ;
assign n2756 =  ( n2755 ) == ( bv_8_163_n340 )  ;
assign n2757 = in[31:24] ;
assign n2758 =  ( n2757 ) == ( bv_8_162_n344 )  ;
assign n2759 = in[31:24] ;
assign n2760 =  ( n2759 ) == ( bv_8_161_n62 )  ;
assign n2761 = in[31:24] ;
assign n2762 =  ( n2761 ) == ( bv_8_160_n351 )  ;
assign n2763 = in[31:24] ;
assign n2764 =  ( n2763 ) == ( bv_8_159_n354 )  ;
assign n2765 = in[31:24] ;
assign n2766 =  ( n2765 ) == ( bv_8_158_n129 )  ;
assign n2767 = in[31:24] ;
assign n2768 =  ( n2767 ) == ( bv_8_157_n360 )  ;
assign n2769 = in[31:24] ;
assign n2770 =  ( n2769 ) == ( bv_8_156_n364 )  ;
assign n2771 = in[31:24] ;
assign n2772 =  ( n2771 ) == ( bv_8_155_n97 )  ;
assign n2773 = in[31:24] ;
assign n2774 =  ( n2773 ) == ( bv_8_154_n370 )  ;
assign n2775 = in[31:24] ;
assign n2776 =  ( n2775 ) == ( bv_8_153_n30 )  ;
assign n2777 = in[31:24] ;
assign n2778 =  ( n2777 ) == ( bv_8_152_n120 )  ;
assign n2779 = in[31:24] ;
assign n2780 =  ( n2779 ) == ( bv_8_151_n378 )  ;
assign n2781 = in[31:24] ;
assign n2782 =  ( n2781 ) == ( bv_8_150_n382 )  ;
assign n2783 = in[31:24] ;
assign n2784 =  ( n2783 ) == ( bv_8_149_n307 )  ;
assign n2785 = in[31:24] ;
assign n2786 =  ( n2785 ) == ( bv_8_148_n101 )  ;
assign n2787 = in[31:24] ;
assign n2788 =  ( n2787 ) == ( bv_8_147_n392 )  ;
assign n2789 = in[31:24] ;
assign n2790 =  ( n2789 ) == ( bv_8_146_n395 )  ;
assign n2791 = in[31:24] ;
assign n2792 =  ( n2791 ) == ( bv_8_145_n311 )  ;
assign n2793 = in[31:24] ;
assign n2794 =  ( n2793 ) == ( bv_8_144_n384 )  ;
assign n2795 = in[31:24] ;
assign n2796 =  ( n2795 ) == ( bv_8_143_n405 )  ;
assign n2797 = in[31:24] ;
assign n2798 =  ( n2797 ) == ( bv_8_142_n104 )  ;
assign n2799 = in[31:24] ;
assign n2800 =  ( n2799 ) == ( bv_8_141_n284 )  ;
assign n2801 = in[31:24] ;
assign n2802 =  ( n2801 ) == ( bv_8_140_n66 )  ;
assign n2803 = in[31:24] ;
assign n2804 =  ( n2803 ) == ( bv_8_139_n194 )  ;
assign n2805 = in[31:24] ;
assign n2806 =  ( n2805 ) == ( bv_8_138_n191 )  ;
assign n2807 = in[31:24] ;
assign n2808 =  ( n2807 ) == ( bv_8_137_n58 )  ;
assign n2809 = in[31:24] ;
assign n2810 =  ( n2809 ) == ( bv_8_136_n380 )  ;
assign n2811 = in[31:24] ;
assign n2812 =  ( n2811 ) == ( bv_8_135_n90 )  ;
assign n2813 = in[31:24] ;
assign n2814 =  ( n2813 ) == ( bv_8_134_n141 )  ;
assign n2815 = in[31:24] ;
assign n2816 =  ( n2815 ) == ( bv_8_133_n434 )  ;
assign n2817 = in[31:24] ;
assign n2818 =  ( n2817 ) == ( bv_8_132_n437 )  ;
assign n2819 = in[31:24] ;
assign n2820 =  ( n2819 ) == ( bv_8_131_n441 )  ;
assign n2821 = in[31:24] ;
assign n2822 =  ( n2821 ) == ( bv_8_130_n444 )  ;
assign n2823 = in[31:24] ;
assign n2824 =  ( n2823 ) == ( bv_8_129_n400 )  ;
assign n2825 = in[31:24] ;
assign n2826 =  ( n2825 ) == ( bv_8_128_n451 )  ;
assign n2827 = in[31:24] ;
assign n2828 =  ( n2827 ) == ( bv_8_127_n454 )  ;
assign n2829 = in[31:24] ;
assign n2830 =  ( n2829 ) == ( bv_8_126_n422 )  ;
assign n2831 = in[31:24] ;
assign n2832 =  ( n2831 ) == ( bv_8_125_n459 )  ;
assign n2833 = in[31:24] ;
assign n2834 =  ( n2833 ) == ( bv_8_124_n462 )  ;
assign n2835 = in[31:24] ;
assign n2836 =  ( n2835 ) == ( bv_8_123_n466 )  ;
assign n2837 = in[31:24] ;
assign n2838 =  ( n2837 ) == ( bv_8_122_n256 )  ;
assign n2839 = in[31:24] ;
assign n2840 =  ( n2839 ) == ( bv_8_121_n301 )  ;
assign n2841 = in[31:24] ;
assign n2842 =  ( n2841 ) == ( bv_8_120_n242 )  ;
assign n2843 = in[31:24] ;
assign n2844 =  ( n2843 ) == ( bv_8_119_n476 )  ;
assign n2845 = in[31:24] ;
assign n2846 =  ( n2845 ) == ( bv_8_118_n479 )  ;
assign n2847 = in[31:24] ;
assign n2848 =  ( n2847 ) == ( bv_8_117_n483 )  ;
assign n2849 = in[31:24] ;
assign n2850 =  ( n2849 ) == ( bv_8_116_n210 )  ;
assign n2851 = in[31:24] ;
assign n2852 =  ( n2851 ) == ( bv_8_115_n407 )  ;
assign n2853 = in[31:24] ;
assign n2854 =  ( n2853 ) == ( bv_8_114_n490 )  ;
assign n2855 = in[31:24] ;
assign n2856 =  ( n2855 ) == ( bv_8_113_n494 )  ;
assign n2857 = in[31:24] ;
assign n2858 =  ( n2857 ) == ( bv_8_112_n187 )  ;
assign n2859 = in[31:24] ;
assign n2860 =  ( n2859 ) == ( bv_8_111_n500 )  ;
assign n2861 = in[31:24] ;
assign n2862 =  ( n2861 ) == ( bv_8_110_n503 )  ;
assign n2863 = in[31:24] ;
assign n2864 =  ( n2863 ) == ( bv_8_109_n288 )  ;
assign n2865 = in[31:24] ;
assign n2866 =  ( n2865 ) == ( bv_8_108_n271 )  ;
assign n2867 = in[31:24] ;
assign n2868 =  ( n2867 ) == ( bv_8_107_n512 )  ;
assign n2869 = in[31:24] ;
assign n2870 =  ( n2869 ) == ( bv_8_106_n515 )  ;
assign n2871 = in[31:24] ;
assign n2872 =  ( n2871 ) == ( bv_8_105_n112 )  ;
assign n2873 = in[31:24] ;
assign n2874 =  ( n2873 ) == ( bv_8_104_n38 )  ;
assign n2875 = in[31:24] ;
assign n2876 =  ( n2875 ) == ( bv_8_103_n524 )  ;
assign n2877 = in[31:24] ;
assign n2878 =  ( n2877 ) == ( bv_8_102_n175 )  ;
assign n2879 = in[31:24] ;
assign n2880 =  ( n2879 ) == ( bv_8_101_n260 )  ;
assign n2881 = in[31:24] ;
assign n2882 =  ( n2881 ) == ( bv_8_100_n416 )  ;
assign n2883 = in[31:24] ;
assign n2884 =  ( n2883 ) == ( bv_8_99_n536 )  ;
assign n2885 = in[31:24] ;
assign n2886 =  ( n2885 ) == ( bv_8_98_n315 )  ;
assign n2887 = in[31:24] ;
assign n2888 =  ( n2887 ) == ( bv_8_97_n156 )  ;
assign n2889 = in[31:24] ;
assign n2890 =  ( n2889 ) == ( bv_8_96_n403 )  ;
assign n2891 = in[31:24] ;
assign n2892 =  ( n2891 ) == ( bv_8_95_n439 )  ;
assign n2893 = in[31:24] ;
assign n2894 =  ( n2893 ) == ( bv_8_94_n362 )  ;
assign n2895 = in[31:24] ;
assign n2896 =  ( n2895 ) == ( bv_8_93_n413 )  ;
assign n2897 = in[31:24] ;
assign n2898 =  ( n2897 ) == ( bv_8_92_n327 )  ;
assign n2899 = in[31:24] ;
assign n2900 =  ( n2899 ) == ( bv_8_91_n556 )  ;
assign n2901 = in[31:24] ;
assign n2902 =  ( n2901 ) == ( bv_8_90_n560 )  ;
assign n2903 = in[31:24] ;
assign n2904 =  ( n2903 ) == ( bv_8_89_n563 )  ;
assign n2905 = in[31:24] ;
assign n2906 =  ( n2905 ) == ( bv_8_88_n548 )  ;
assign n2907 = in[31:24] ;
assign n2908 =  ( n2907 ) == ( bv_8_87_n149 )  ;
assign n2909 = in[31:24] ;
assign n2910 =  ( n2909 ) == ( bv_8_86_n267 )  ;
assign n2911 = in[31:24] ;
assign n2912 =  ( n2911 ) == ( bv_8_85_n78 )  ;
assign n2913 = in[31:24] ;
assign n2914 =  ( n2913 ) == ( bv_8_84_n14 )  ;
assign n2915 = in[31:24] ;
assign n2916 =  ( n2915 ) == ( bv_8_83_n577 )  ;
assign n2917 = in[31:24] ;
assign n2918 =  ( n2917 ) == ( bv_8_82_n580 )  ;
assign n2919 = in[31:24] ;
assign n2920 =  ( n2919 ) == ( bv_8_81_n498 )  ;
assign n2921 = in[31:24] ;
assign n2922 =  ( n2921 ) == ( bv_8_80_n510 )  ;
assign n2923 = in[31:24] ;
assign n2924 =  ( n2923 ) == ( bv_8_79_n397 )  ;
assign n2925 = in[31:24] ;
assign n2926 =  ( n2925 ) == ( bv_8_78_n279 )  ;
assign n2927 = in[31:24] ;
assign n2928 =  ( n2927 ) == ( bv_8_77_n531 )  ;
assign n2929 = in[31:24] ;
assign n2930 =  ( n2929 ) == ( bv_8_76_n551 )  ;
assign n2931 = in[31:24] ;
assign n2932 =  ( n2931 ) == ( bv_8_75_n202 )  ;
assign n2933 = in[31:24] ;
assign n2934 =  ( n2933 ) == ( bv_8_74_n554 )  ;
assign n2935 = in[31:24] ;
assign n2936 =  ( n2935 ) == ( bv_8_73_n338 )  ;
assign n2937 = in[31:24] ;
assign n2938 =  ( n2937 ) == ( bv_8_72_n171 )  ;
assign n2939 = in[31:24] ;
assign n2940 =  ( n2939 ) == ( bv_8_71_n607 )  ;
assign n2941 = in[31:24] ;
assign n2942 =  ( n2941 ) == ( bv_8_70_n376 )  ;
assign n2943 = in[31:24] ;
assign n2944 =  ( n2943 ) == ( bv_8_69_n522 )  ;
assign n2945 = in[31:24] ;
assign n2946 =  ( n2945 ) == ( bv_8_68_n432 )  ;
assign n2947 = in[31:24] ;
assign n2948 =  ( n2947 ) == ( bv_8_67_n534 )  ;
assign n2949 = in[31:24] ;
assign n2950 =  ( n2949 ) == ( bv_8_66_n42 )  ;
assign n2951 = in[31:24] ;
assign n2952 =  ( n2951 ) == ( bv_8_65_n34 )  ;
assign n2953 = in[31:24] ;
assign n2954 =  ( n2953 ) == ( bv_8_64_n492 )  ;
assign n2955 = in[31:24] ;
assign n2956 =  ( n2955 ) == ( bv_8_63_n628 )  ;
assign n2957 = in[31:24] ;
assign n2958 =  ( n2957 ) == ( bv_8_62_n183 )  ;
assign n2959 = in[31:24] ;
assign n2960 =  ( n2959 ) == ( bv_8_61_n419 )  ;
assign n2961 = in[31:24] ;
assign n2962 =  ( n2961 ) == ( bv_8_60_n507 )  ;
assign n2963 = in[31:24] ;
assign n2964 =  ( n2963 ) == ( bv_8_59_n603 )  ;
assign n2965 = in[31:24] ;
assign n2966 =  ( n2965 ) == ( bv_8_58_n346 )  ;
assign n2967 = in[31:24] ;
assign n2968 =  ( n2967 ) == ( bv_8_57_n558 )  ;
assign n2969 = in[31:24] ;
assign n2970 =  ( n2969 ) == ( bv_8_56_n481 )  ;
assign n2971 = in[31:24] ;
assign n2972 =  ( n2971 ) == ( bv_8_55_n292 )  ;
assign n2973 = in[31:24] ;
assign n2974 =  ( n2973 ) == ( bv_8_54_n650 )  ;
assign n2975 = in[31:24] ;
assign n2976 =  ( n2975 ) == ( bv_8_53_n152 )  ;
assign n2977 = in[31:24] ;
assign n2978 =  ( n2977 ) == ( bv_8_52_n656 )  ;
assign n2979 = in[31:24] ;
assign n2980 =  ( n2979 ) == ( bv_8_51_n528 )  ;
assign n2981 = in[31:24] ;
assign n2982 =  ( n2981 ) == ( bv_8_50_n349 )  ;
assign n2983 = in[31:24] ;
assign n2984 =  ( n2983 ) == ( bv_8_49_n665 )  ;
assign n2985 = in[31:24] ;
assign n2986 =  ( n2985 ) == ( bv_8_48_n668 )  ;
assign n2987 = in[31:24] ;
assign n2988 =  ( n2987 ) == ( bv_8_47_n591 )  ;
assign n2989 = in[31:24] ;
assign n2990 =  ( n2989 ) == ( bv_8_46_n235 )  ;
assign n2991 = in[31:24] ;
assign n2992 =  ( n2991 ) == ( bv_8_45_n26 )  ;
assign n2993 = in[31:24] ;
assign n2994 =  ( n2993 ) == ( bv_8_44_n621 )  ;
assign n2995 = in[31:24] ;
assign n2996 =  ( n2995 ) == ( bv_8_43_n681 )  ;
assign n2997 = in[31:24] ;
assign n2998 =  ( n2997 ) == ( bv_8_42_n387 )  ;
assign n2999 = in[31:24] ;
assign n3000 =  ( n2999 ) == ( bv_8_41_n596 )  ;
assign n3001 = in[31:24] ;
assign n3002 =  ( n3001 ) == ( bv_8_40_n74 )  ;
assign n3003 = in[31:24] ;
assign n3004 =  ( n3003 ) == ( bv_8_39_n634 )  ;
assign n3005 = in[31:24] ;
assign n3006 =  ( n3005 ) == ( bv_8_38_n692 )  ;
assign n3007 = in[31:24] ;
assign n3008 =  ( n3007 ) == ( bv_8_37_n239 )  ;
assign n3009 = in[31:24] ;
assign n3010 =  ( n3009 ) == ( bv_8_36_n330 )  ;
assign n3011 = in[31:24] ;
assign n3012 =  ( n3011 ) == ( bv_8_35_n663 )  ;
assign n3013 = in[31:24] ;
assign n3014 =  ( n3013 ) == ( bv_8_34_n390 )  ;
assign n3015 = in[31:24] ;
assign n3016 =  ( n3015 ) == ( bv_8_33_n468 )  ;
assign n3017 = in[31:24] ;
assign n3018 =  ( n3017 ) == ( bv_8_32_n575 )  ;
assign n3019 = in[31:24] ;
assign n3020 =  ( n3019 ) == ( bv_8_31_n206 )  ;
assign n3021 = in[31:24] ;
assign n3022 =  ( n3021 ) == ( bv_8_30_n93 )  ;
assign n3023 = in[31:24] ;
assign n3024 =  ( n3023 ) == ( bv_8_29_n133 )  ;
assign n3025 = in[31:24] ;
assign n3026 =  ( n3025 ) == ( bv_8_28_n231 )  ;
assign n3027 = in[31:24] ;
assign n3028 =  ( n3027 ) == ( bv_8_27_n615 )  ;
assign n3029 = in[31:24] ;
assign n3030 =  ( n3029 ) == ( bv_8_26_n618 )  ;
assign n3031 = in[31:24] ;
assign n3032 =  ( n3031 ) == ( bv_8_25_n410 )  ;
assign n3033 = in[31:24] ;
assign n3034 =  ( n3033 ) == ( bv_8_24_n658 )  ;
assign n3035 = in[31:24] ;
assign n3036 =  ( n3035 ) == ( bv_8_23_n429 )  ;
assign n3037 = in[31:24] ;
assign n3038 =  ( n3037 ) == ( bv_8_22_n6 )  ;
assign n3039 = in[31:24] ;
assign n3040 =  ( n3039 ) == ( bv_8_21_n673 )  ;
assign n3041 = in[31:24] ;
assign n3042 =  ( n3041 ) == ( bv_8_20_n368 )  ;
assign n3043 = in[31:24] ;
assign n3044 =  ( n3043 ) == ( bv_8_19_n446 )  ;
assign n3045 = in[31:24] ;
assign n3046 =  ( n3045 ) == ( bv_8_18_n643 )  ;
assign n3047 = in[31:24] ;
assign n3048 =  ( n3047 ) == ( bv_8_17_n116 )  ;
assign n3049 = in[31:24] ;
assign n3050 =  ( n3049 ) == ( bv_8_16_n464 )  ;
assign n3051 = in[31:24] ;
assign n3052 =  ( n3051 ) == ( bv_8_15_n22 )  ;
assign n3053 = in[31:24] ;
assign n3054 =  ( n3053 ) == ( bv_8_14_n160 )  ;
assign n3055 = in[31:24] ;
assign n3056 =  ( n3055 ) == ( bv_8_13_n54 )  ;
assign n3057 = in[31:24] ;
assign n3058 =  ( n3057 ) == ( bv_8_12_n449 )  ;
assign n3059 = in[31:24] ;
assign n3060 =  ( n3059 ) == ( bv_8_11_n358 )  ;
assign n3061 = in[31:24] ;
assign n3062 =  ( n3061 ) == ( bv_8_10_n342 )  ;
assign n3063 = in[31:24] ;
assign n3064 =  ( n3063 ) == ( bv_8_9_n626 )  ;
assign n3065 = in[31:24] ;
assign n3066 =  ( n3065 ) == ( bv_8_8_n249 )  ;
assign n3067 = in[31:24] ;
assign n3068 =  ( n3067 ) == ( bv_8_7_n646 )  ;
assign n3069 = in[31:24] ;
assign n3070 =  ( n3069 ) == ( bv_8_6_n334 )  ;
assign n3071 = in[31:24] ;
assign n3072 =  ( n3071 ) == ( bv_8_5_n652 )  ;
assign n3073 = in[31:24] ;
assign n3074 =  ( n3073 ) == ( bv_8_4_n670 )  ;
assign n3075 = in[31:24] ;
assign n3076 =  ( n3075 ) == ( bv_8_3_n167 )  ;
assign n3077 = in[31:24] ;
assign n3078 =  ( n3077 ) == ( bv_8_2_n517 )  ;
assign n3079 = in[31:24] ;
assign n3080 =  ( n3079 ) == ( bv_8_1_n752 )  ;
assign n3081 = in[31:24] ;
assign n3082 =  ( n3081 ) == ( bv_8_0_n582 )  ;
assign n3083 =  ( n3082 ) ? ( bv_8_99_n536 ) : ( bv_8_0_n582 ) ;
assign n3084 =  ( n3080 ) ? ( bv_8_124_n462 ) : ( n3083 ) ;
assign n3085 =  ( n3078 ) ? ( bv_8_119_n476 ) : ( n3084 ) ;
assign n3086 =  ( n3076 ) ? ( bv_8_123_n466 ) : ( n3085 ) ;
assign n3087 =  ( n3074 ) ? ( bv_8_242_n56 ) : ( n3086 ) ;
assign n3088 =  ( n3072 ) ? ( bv_8_107_n512 ) : ( n3087 ) ;
assign n3089 =  ( n3070 ) ? ( bv_8_111_n500 ) : ( n3088 ) ;
assign n3090 =  ( n3068 ) ? ( bv_8_197_n225 ) : ( n3089 ) ;
assign n3091 =  ( n3066 ) ? ( bv_8_48_n668 ) : ( n3090 ) ;
assign n3092 =  ( n3064 ) ? ( bv_8_1_n752 ) : ( n3091 ) ;
assign n3093 =  ( n3062 ) ? ( bv_8_103_n524 ) : ( n3092 ) ;
assign n3094 =  ( n3060 ) ? ( bv_8_43_n681 ) : ( n3093 ) ;
assign n3095 =  ( n3058 ) ? ( bv_8_254_n8 ) : ( n3094 ) ;
assign n3096 =  ( n3056 ) ? ( bv_8_215_n158 ) : ( n3095 ) ;
assign n3097 =  ( n3054 ) ? ( bv_8_171_n313 ) : ( n3096 ) ;
assign n3098 =  ( n3052 ) ? ( bv_8_118_n479 ) : ( n3097 ) ;
assign n3099 =  ( n3050 ) ? ( bv_8_202_n208 ) : ( n3098 ) ;
assign n3100 =  ( n3048 ) ? ( bv_8_130_n444 ) : ( n3099 ) ;
assign n3101 =  ( n3046 ) ? ( bv_8_201_n212 ) : ( n3100 ) ;
assign n3102 =  ( n3044 ) ? ( bv_8_125_n459 ) : ( n3101 ) ;
assign n3103 =  ( n3042 ) ? ( bv_8_250_n24 ) : ( n3102 ) ;
assign n3104 =  ( n3040 ) ? ( bv_8_89_n563 ) : ( n3103 ) ;
assign n3105 =  ( n3038 ) ? ( bv_8_71_n607 ) : ( n3104 ) ;
assign n3106 =  ( n3036 ) ? ( bv_8_240_n64 ) : ( n3105 ) ;
assign n3107 =  ( n3034 ) ? ( bv_8_173_n305 ) : ( n3106 ) ;
assign n3108 =  ( n3032 ) ? ( bv_8_212_n169 ) : ( n3107 ) ;
assign n3109 =  ( n3030 ) ? ( bv_8_162_n344 ) : ( n3108 ) ;
assign n3110 =  ( n3028 ) ? ( bv_8_175_n299 ) : ( n3109 ) ;
assign n3111 =  ( n3026 ) ? ( bv_8_156_n364 ) : ( n3110 ) ;
assign n3112 =  ( n3024 ) ? ( bv_8_164_n336 ) : ( n3111 ) ;
assign n3113 =  ( n3022 ) ? ( bv_8_114_n490 ) : ( n3112 ) ;
assign n3114 =  ( n3020 ) ? ( bv_8_192_n244 ) : ( n3113 ) ;
assign n3115 =  ( n3018 ) ? ( bv_8_183_n273 ) : ( n3114 ) ;
assign n3116 =  ( n3016 ) ? ( bv_8_253_n12 ) : ( n3115 ) ;
assign n3117 =  ( n3014 ) ? ( bv_8_147_n392 ) : ( n3116 ) ;
assign n3118 =  ( n3012 ) ? ( bv_8_38_n692 ) : ( n3117 ) ;
assign n3119 =  ( n3010 ) ? ( bv_8_54_n650 ) : ( n3118 ) ;
assign n3120 =  ( n3008 ) ? ( bv_8_63_n628 ) : ( n3119 ) ;
assign n3121 =  ( n3006 ) ? ( bv_8_247_n36 ) : ( n3120 ) ;
assign n3122 =  ( n3004 ) ? ( bv_8_204_n200 ) : ( n3121 ) ;
assign n3123 =  ( n3002 ) ? ( bv_8_52_n656 ) : ( n3122 ) ;
assign n3124 =  ( n3000 ) ? ( bv_8_165_n332 ) : ( n3123 ) ;
assign n3125 =  ( n2998 ) ? ( bv_8_229_n106 ) : ( n3124 ) ;
assign n3126 =  ( n2996 ) ? ( bv_8_241_n60 ) : ( n3125 ) ;
assign n3127 =  ( n2994 ) ? ( bv_8_113_n494 ) : ( n3126 ) ;
assign n3128 =  ( n2992 ) ? ( bv_8_216_n154 ) : ( n3127 ) ;
assign n3129 =  ( n2990 ) ? ( bv_8_49_n665 ) : ( n3128 ) ;
assign n3130 =  ( n2988 ) ? ( bv_8_21_n673 ) : ( n3129 ) ;
assign n3131 =  ( n2986 ) ? ( bv_8_4_n670 ) : ( n3130 ) ;
assign n3132 =  ( n2984 ) ? ( bv_8_199_n218 ) : ( n3131 ) ;
assign n3133 =  ( n2982 ) ? ( bv_8_35_n663 ) : ( n3132 ) ;
assign n3134 =  ( n2980 ) ? ( bv_8_195_n233 ) : ( n3133 ) ;
assign n3135 =  ( n2978 ) ? ( bv_8_24_n658 ) : ( n3134 ) ;
assign n3136 =  ( n2976 ) ? ( bv_8_150_n382 ) : ( n3135 ) ;
assign n3137 =  ( n2974 ) ? ( bv_8_5_n652 ) : ( n3136 ) ;
assign n3138 =  ( n2972 ) ? ( bv_8_154_n370 ) : ( n3137 ) ;
assign n3139 =  ( n2970 ) ? ( bv_8_7_n646 ) : ( n3138 ) ;
assign n3140 =  ( n2968 ) ? ( bv_8_18_n643 ) : ( n3139 ) ;
assign n3141 =  ( n2966 ) ? ( bv_8_128_n451 ) : ( n3140 ) ;
assign n3142 =  ( n2964 ) ? ( bv_8_226_n118 ) : ( n3141 ) ;
assign n3143 =  ( n2962 ) ? ( bv_8_235_n84 ) : ( n3142 ) ;
assign n3144 =  ( n2960 ) ? ( bv_8_39_n634 ) : ( n3143 ) ;
assign n3145 =  ( n2958 ) ? ( bv_8_178_n290 ) : ( n3144 ) ;
assign n3146 =  ( n2956 ) ? ( bv_8_117_n483 ) : ( n3145 ) ;
assign n3147 =  ( n2954 ) ? ( bv_8_9_n626 ) : ( n3146 ) ;
assign n3148 =  ( n2952 ) ? ( bv_8_131_n441 ) : ( n3147 ) ;
assign n3149 =  ( n2950 ) ? ( bv_8_44_n621 ) : ( n3148 ) ;
assign n3150 =  ( n2948 ) ? ( bv_8_26_n618 ) : ( n3149 ) ;
assign n3151 =  ( n2946 ) ? ( bv_8_27_n615 ) : ( n3150 ) ;
assign n3152 =  ( n2944 ) ? ( bv_8_110_n503 ) : ( n3151 ) ;
assign n3153 =  ( n2942 ) ? ( bv_8_90_n560 ) : ( n3152 ) ;
assign n3154 =  ( n2940 ) ? ( bv_8_160_n351 ) : ( n3153 ) ;
assign n3155 =  ( n2938 ) ? ( bv_8_82_n580 ) : ( n3154 ) ;
assign n3156 =  ( n2936 ) ? ( bv_8_59_n603 ) : ( n3155 ) ;
assign n3157 =  ( n2934 ) ? ( bv_8_214_n162 ) : ( n3156 ) ;
assign n3158 =  ( n2932 ) ? ( bv_8_179_n286 ) : ( n3157 ) ;
assign n3159 =  ( n2930 ) ? ( bv_8_41_n596 ) : ( n3158 ) ;
assign n3160 =  ( n2928 ) ? ( bv_8_227_n114 ) : ( n3159 ) ;
assign n3161 =  ( n2926 ) ? ( bv_8_47_n591 ) : ( n3160 ) ;
assign n3162 =  ( n2924 ) ? ( bv_8_132_n437 ) : ( n3161 ) ;
assign n3163 =  ( n2922 ) ? ( bv_8_83_n577 ) : ( n3162 ) ;
assign n3164 =  ( n2920 ) ? ( bv_8_209_n181 ) : ( n3163 ) ;
assign n3165 =  ( n2918 ) ? ( bv_8_0_n582 ) : ( n3164 ) ;
assign n3166 =  ( n2916 ) ? ( bv_8_237_n76 ) : ( n3165 ) ;
assign n3167 =  ( n2914 ) ? ( bv_8_32_n575 ) : ( n3166 ) ;
assign n3168 =  ( n2912 ) ? ( bv_8_252_n16 ) : ( n3167 ) ;
assign n3169 =  ( n2910 ) ? ( bv_8_177_n294 ) : ( n3168 ) ;
assign n3170 =  ( n2908 ) ? ( bv_8_91_n556 ) : ( n3169 ) ;
assign n3171 =  ( n2906 ) ? ( bv_8_106_n515 ) : ( n3170 ) ;
assign n3172 =  ( n2904 ) ? ( bv_8_203_n204 ) : ( n3171 ) ;
assign n3173 =  ( n2902 ) ? ( bv_8_190_n251 ) : ( n3172 ) ;
assign n3174 =  ( n2900 ) ? ( bv_8_57_n558 ) : ( n3173 ) ;
assign n3175 =  ( n2898 ) ? ( bv_8_74_n554 ) : ( n3174 ) ;
assign n3176 =  ( n2896 ) ? ( bv_8_76_n551 ) : ( n3175 ) ;
assign n3177 =  ( n2894 ) ? ( bv_8_88_n548 ) : ( n3176 ) ;
assign n3178 =  ( n2892 ) ? ( bv_8_207_n189 ) : ( n3177 ) ;
assign n3179 =  ( n2890 ) ? ( bv_8_208_n185 ) : ( n3178 ) ;
assign n3180 =  ( n2888 ) ? ( bv_8_239_n68 ) : ( n3179 ) ;
assign n3181 =  ( n2886 ) ? ( bv_8_170_n317 ) : ( n3180 ) ;
assign n3182 =  ( n2884 ) ? ( bv_8_251_n20 ) : ( n3181 ) ;
assign n3183 =  ( n2882 ) ? ( bv_8_67_n534 ) : ( n3182 ) ;
assign n3184 =  ( n2880 ) ? ( bv_8_77_n531 ) : ( n3183 ) ;
assign n3185 =  ( n2878 ) ? ( bv_8_51_n528 ) : ( n3184 ) ;
assign n3186 =  ( n2876 ) ? ( bv_8_133_n434 ) : ( n3185 ) ;
assign n3187 =  ( n2874 ) ? ( bv_8_69_n522 ) : ( n3186 ) ;
assign n3188 =  ( n2872 ) ? ( bv_8_249_n28 ) : ( n3187 ) ;
assign n3189 =  ( n2870 ) ? ( bv_8_2_n517 ) : ( n3188 ) ;
assign n3190 =  ( n2868 ) ? ( bv_8_127_n454 ) : ( n3189 ) ;
assign n3191 =  ( n2866 ) ? ( bv_8_80_n510 ) : ( n3190 ) ;
assign n3192 =  ( n2864 ) ? ( bv_8_60_n507 ) : ( n3191 ) ;
assign n3193 =  ( n2862 ) ? ( bv_8_159_n354 ) : ( n3192 ) ;
assign n3194 =  ( n2860 ) ? ( bv_8_168_n322 ) : ( n3193 ) ;
assign n3195 =  ( n2858 ) ? ( bv_8_81_n498 ) : ( n3194 ) ;
assign n3196 =  ( n2856 ) ? ( bv_8_163_n340 ) : ( n3195 ) ;
assign n3197 =  ( n2854 ) ? ( bv_8_64_n492 ) : ( n3196 ) ;
assign n3198 =  ( n2852 ) ? ( bv_8_143_n405 ) : ( n3197 ) ;
assign n3199 =  ( n2850 ) ? ( bv_8_146_n395 ) : ( n3198 ) ;
assign n3200 =  ( n2848 ) ? ( bv_8_157_n360 ) : ( n3199 ) ;
assign n3201 =  ( n2846 ) ? ( bv_8_56_n481 ) : ( n3200 ) ;
assign n3202 =  ( n2844 ) ? ( bv_8_245_n44 ) : ( n3201 ) ;
assign n3203 =  ( n2842 ) ? ( bv_8_188_n258 ) : ( n3202 ) ;
assign n3204 =  ( n2840 ) ? ( bv_8_182_n277 ) : ( n3203 ) ;
assign n3205 =  ( n2838 ) ? ( bv_8_218_n147 ) : ( n3204 ) ;
assign n3206 =  ( n2836 ) ? ( bv_8_33_n468 ) : ( n3205 ) ;
assign n3207 =  ( n2834 ) ? ( bv_8_16_n464 ) : ( n3206 ) ;
assign n3208 =  ( n2832 ) ? ( bv_8_255_n4 ) : ( n3207 ) ;
assign n3209 =  ( n2830 ) ? ( bv_8_243_n52 ) : ( n3208 ) ;
assign n3210 =  ( n2828 ) ? ( bv_8_210_n177 ) : ( n3209 ) ;
assign n3211 =  ( n2826 ) ? ( bv_8_205_n196 ) : ( n3210 ) ;
assign n3212 =  ( n2824 ) ? ( bv_8_12_n449 ) : ( n3211 ) ;
assign n3213 =  ( n2822 ) ? ( bv_8_19_n446 ) : ( n3212 ) ;
assign n3214 =  ( n2820 ) ? ( bv_8_236_n80 ) : ( n3213 ) ;
assign n3215 =  ( n2818 ) ? ( bv_8_95_n439 ) : ( n3214 ) ;
assign n3216 =  ( n2816 ) ? ( bv_8_151_n378 ) : ( n3215 ) ;
assign n3217 =  ( n2814 ) ? ( bv_8_68_n432 ) : ( n3216 ) ;
assign n3218 =  ( n2812 ) ? ( bv_8_23_n429 ) : ( n3217 ) ;
assign n3219 =  ( n2810 ) ? ( bv_8_196_n229 ) : ( n3218 ) ;
assign n3220 =  ( n2808 ) ? ( bv_8_167_n325 ) : ( n3219 ) ;
assign n3221 =  ( n2806 ) ? ( bv_8_126_n422 ) : ( n3220 ) ;
assign n3222 =  ( n2804 ) ? ( bv_8_61_n419 ) : ( n3221 ) ;
assign n3223 =  ( n2802 ) ? ( bv_8_100_n416 ) : ( n3222 ) ;
assign n3224 =  ( n2800 ) ? ( bv_8_93_n413 ) : ( n3223 ) ;
assign n3225 =  ( n2798 ) ? ( bv_8_25_n410 ) : ( n3224 ) ;
assign n3226 =  ( n2796 ) ? ( bv_8_115_n407 ) : ( n3225 ) ;
assign n3227 =  ( n2794 ) ? ( bv_8_96_n403 ) : ( n3226 ) ;
assign n3228 =  ( n2792 ) ? ( bv_8_129_n400 ) : ( n3227 ) ;
assign n3229 =  ( n2790 ) ? ( bv_8_79_n397 ) : ( n3228 ) ;
assign n3230 =  ( n2788 ) ? ( bv_8_220_n139 ) : ( n3229 ) ;
assign n3231 =  ( n2786 ) ? ( bv_8_34_n390 ) : ( n3230 ) ;
assign n3232 =  ( n2784 ) ? ( bv_8_42_n387 ) : ( n3231 ) ;
assign n3233 =  ( n2782 ) ? ( bv_8_144_n384 ) : ( n3232 ) ;
assign n3234 =  ( n2780 ) ? ( bv_8_136_n380 ) : ( n3233 ) ;
assign n3235 =  ( n2778 ) ? ( bv_8_70_n376 ) : ( n3234 ) ;
assign n3236 =  ( n2776 ) ? ( bv_8_238_n72 ) : ( n3235 ) ;
assign n3237 =  ( n2774 ) ? ( bv_8_184_n269 ) : ( n3236 ) ;
assign n3238 =  ( n2772 ) ? ( bv_8_20_n368 ) : ( n3237 ) ;
assign n3239 =  ( n2770 ) ? ( bv_8_222_n131 ) : ( n3238 ) ;
assign n3240 =  ( n2768 ) ? ( bv_8_94_n362 ) : ( n3239 ) ;
assign n3241 =  ( n2766 ) ? ( bv_8_11_n358 ) : ( n3240 ) ;
assign n3242 =  ( n2764 ) ? ( bv_8_219_n143 ) : ( n3241 ) ;
assign n3243 =  ( n2762 ) ? ( bv_8_224_n125 ) : ( n3242 ) ;
assign n3244 =  ( n2760 ) ? ( bv_8_50_n349 ) : ( n3243 ) ;
assign n3245 =  ( n2758 ) ? ( bv_8_58_n346 ) : ( n3244 ) ;
assign n3246 =  ( n2756 ) ? ( bv_8_10_n342 ) : ( n3245 ) ;
assign n3247 =  ( n2754 ) ? ( bv_8_73_n338 ) : ( n3246 ) ;
assign n3248 =  ( n2752 ) ? ( bv_8_6_n334 ) : ( n3247 ) ;
assign n3249 =  ( n2750 ) ? ( bv_8_36_n330 ) : ( n3248 ) ;
assign n3250 =  ( n2748 ) ? ( bv_8_92_n327 ) : ( n3249 ) ;
assign n3251 =  ( n2746 ) ? ( bv_8_194_n237 ) : ( n3250 ) ;
assign n3252 =  ( n2744 ) ? ( bv_8_211_n173 ) : ( n3251 ) ;
assign n3253 =  ( n2742 ) ? ( bv_8_172_n309 ) : ( n3252 ) ;
assign n3254 =  ( n2740 ) ? ( bv_8_98_n315 ) : ( n3253 ) ;
assign n3255 =  ( n2738 ) ? ( bv_8_145_n311 ) : ( n3254 ) ;
assign n3256 =  ( n2736 ) ? ( bv_8_149_n307 ) : ( n3255 ) ;
assign n3257 =  ( n2734 ) ? ( bv_8_228_n110 ) : ( n3256 ) ;
assign n3258 =  ( n2732 ) ? ( bv_8_121_n301 ) : ( n3257 ) ;
assign n3259 =  ( n2730 ) ? ( bv_8_231_n99 ) : ( n3258 ) ;
assign n3260 =  ( n2728 ) ? ( bv_8_200_n215 ) : ( n3259 ) ;
assign n3261 =  ( n2726 ) ? ( bv_8_55_n292 ) : ( n3260 ) ;
assign n3262 =  ( n2724 ) ? ( bv_8_109_n288 ) : ( n3261 ) ;
assign n3263 =  ( n2722 ) ? ( bv_8_141_n284 ) : ( n3262 ) ;
assign n3264 =  ( n2720 ) ? ( bv_8_213_n165 ) : ( n3263 ) ;
assign n3265 =  ( n2718 ) ? ( bv_8_78_n279 ) : ( n3264 ) ;
assign n3266 =  ( n2716 ) ? ( bv_8_169_n275 ) : ( n3265 ) ;
assign n3267 =  ( n2714 ) ? ( bv_8_108_n271 ) : ( n3266 ) ;
assign n3268 =  ( n2712 ) ? ( bv_8_86_n267 ) : ( n3267 ) ;
assign n3269 =  ( n2710 ) ? ( bv_8_244_n48 ) : ( n3268 ) ;
assign n3270 =  ( n2708 ) ? ( bv_8_234_n88 ) : ( n3269 ) ;
assign n3271 =  ( n2706 ) ? ( bv_8_101_n260 ) : ( n3270 ) ;
assign n3272 =  ( n2704 ) ? ( bv_8_122_n256 ) : ( n3271 ) ;
assign n3273 =  ( n2702 ) ? ( bv_8_174_n253 ) : ( n3272 ) ;
assign n3274 =  ( n2700 ) ? ( bv_8_8_n249 ) : ( n3273 ) ;
assign n3275 =  ( n2698 ) ? ( bv_8_186_n246 ) : ( n3274 ) ;
assign n3276 =  ( n2696 ) ? ( bv_8_120_n242 ) : ( n3275 ) ;
assign n3277 =  ( n2694 ) ? ( bv_8_37_n239 ) : ( n3276 ) ;
assign n3278 =  ( n2692 ) ? ( bv_8_46_n235 ) : ( n3277 ) ;
assign n3279 =  ( n2690 ) ? ( bv_8_28_n231 ) : ( n3278 ) ;
assign n3280 =  ( n2688 ) ? ( bv_8_166_n227 ) : ( n3279 ) ;
assign n3281 =  ( n2686 ) ? ( bv_8_180_n223 ) : ( n3280 ) ;
assign n3282 =  ( n2684 ) ? ( bv_8_198_n220 ) : ( n3281 ) ;
assign n3283 =  ( n2682 ) ? ( bv_8_232_n95 ) : ( n3282 ) ;
assign n3284 =  ( n2680 ) ? ( bv_8_221_n135 ) : ( n3283 ) ;
assign n3285 =  ( n2678 ) ? ( bv_8_116_n210 ) : ( n3284 ) ;
assign n3286 =  ( n2676 ) ? ( bv_8_31_n206 ) : ( n3285 ) ;
assign n3287 =  ( n2674 ) ? ( bv_8_75_n202 ) : ( n3286 ) ;
assign n3288 =  ( n2672 ) ? ( bv_8_189_n198 ) : ( n3287 ) ;
assign n3289 =  ( n2670 ) ? ( bv_8_139_n194 ) : ( n3288 ) ;
assign n3290 =  ( n2668 ) ? ( bv_8_138_n191 ) : ( n3289 ) ;
assign n3291 =  ( n2666 ) ? ( bv_8_112_n187 ) : ( n3290 ) ;
assign n3292 =  ( n2664 ) ? ( bv_8_62_n183 ) : ( n3291 ) ;
assign n3293 =  ( n2662 ) ? ( bv_8_181_n179 ) : ( n3292 ) ;
assign n3294 =  ( n2660 ) ? ( bv_8_102_n175 ) : ( n3293 ) ;
assign n3295 =  ( n2658 ) ? ( bv_8_72_n171 ) : ( n3294 ) ;
assign n3296 =  ( n2656 ) ? ( bv_8_3_n167 ) : ( n3295 ) ;
assign n3297 =  ( n2654 ) ? ( bv_8_246_n40 ) : ( n3296 ) ;
assign n3298 =  ( n2652 ) ? ( bv_8_14_n160 ) : ( n3297 ) ;
assign n3299 =  ( n2650 ) ? ( bv_8_97_n156 ) : ( n3298 ) ;
assign n3300 =  ( n2648 ) ? ( bv_8_53_n152 ) : ( n3299 ) ;
assign n3301 =  ( n2646 ) ? ( bv_8_87_n149 ) : ( n3300 ) ;
assign n3302 =  ( n2644 ) ? ( bv_8_185_n145 ) : ( n3301 ) ;
assign n3303 =  ( n2642 ) ? ( bv_8_134_n141 ) : ( n3302 ) ;
assign n3304 =  ( n2640 ) ? ( bv_8_193_n137 ) : ( n3303 ) ;
assign n3305 =  ( n2638 ) ? ( bv_8_29_n133 ) : ( n3304 ) ;
assign n3306 =  ( n2636 ) ? ( bv_8_158_n129 ) : ( n3305 ) ;
assign n3307 =  ( n2634 ) ? ( bv_8_225_n122 ) : ( n3306 ) ;
assign n3308 =  ( n2632 ) ? ( bv_8_248_n32 ) : ( n3307 ) ;
assign n3309 =  ( n2630 ) ? ( bv_8_152_n120 ) : ( n3308 ) ;
assign n3310 =  ( n2628 ) ? ( bv_8_17_n116 ) : ( n3309 ) ;
assign n3311 =  ( n2626 ) ? ( bv_8_105_n112 ) : ( n3310 ) ;
assign n3312 =  ( n2624 ) ? ( bv_8_217_n108 ) : ( n3311 ) ;
assign n3313 =  ( n2622 ) ? ( bv_8_142_n104 ) : ( n3312 ) ;
assign n3314 =  ( n2620 ) ? ( bv_8_148_n101 ) : ( n3313 ) ;
assign n3315 =  ( n2618 ) ? ( bv_8_155_n97 ) : ( n3314 ) ;
assign n3316 =  ( n2616 ) ? ( bv_8_30_n93 ) : ( n3315 ) ;
assign n3317 =  ( n2614 ) ? ( bv_8_135_n90 ) : ( n3316 ) ;
assign n3318 =  ( n2612 ) ? ( bv_8_233_n86 ) : ( n3317 ) ;
assign n3319 =  ( n2610 ) ? ( bv_8_206_n82 ) : ( n3318 ) ;
assign n3320 =  ( n2608 ) ? ( bv_8_85_n78 ) : ( n3319 ) ;
assign n3321 =  ( n2606 ) ? ( bv_8_40_n74 ) : ( n3320 ) ;
assign n3322 =  ( n2604 ) ? ( bv_8_223_n70 ) : ( n3321 ) ;
assign n3323 =  ( n2602 ) ? ( bv_8_140_n66 ) : ( n3322 ) ;
assign n3324 =  ( n2600 ) ? ( bv_8_161_n62 ) : ( n3323 ) ;
assign n3325 =  ( n2598 ) ? ( bv_8_137_n58 ) : ( n3324 ) ;
assign n3326 =  ( n2596 ) ? ( bv_8_13_n54 ) : ( n3325 ) ;
assign n3327 =  ( n2594 ) ? ( bv_8_191_n50 ) : ( n3326 ) ;
assign n3328 =  ( n2592 ) ? ( bv_8_230_n46 ) : ( n3327 ) ;
assign n3329 =  ( n2590 ) ? ( bv_8_66_n42 ) : ( n3328 ) ;
assign n3330 =  ( n2588 ) ? ( bv_8_104_n38 ) : ( n3329 ) ;
assign n3331 =  ( n2586 ) ? ( bv_8_65_n34 ) : ( n3330 ) ;
assign n3332 =  ( n2584 ) ? ( bv_8_153_n30 ) : ( n3331 ) ;
assign n3333 =  ( n2582 ) ? ( bv_8_45_n26 ) : ( n3332 ) ;
assign n3334 =  ( n2580 ) ? ( bv_8_15_n22 ) : ( n3333 ) ;
assign n3335 =  ( n2578 ) ? ( bv_8_176_n18 ) : ( n3334 ) ;
assign n3336 =  ( n2576 ) ? ( bv_8_84_n14 ) : ( n3335 ) ;
assign n3337 =  ( n2574 ) ? ( bv_8_187_n10 ) : ( n3336 ) ;
assign n3338 =  ( n2572 ) ? ( bv_8_22_n6 ) : ( n3337 ) ;
assign n3339 =  ( n2570 ) ^ ( n3338 )  ;
assign n3340 =  { ( n2569 ) , ( n3339 ) }  ;
assign n3341 = in[127:120] ;
assign n3342 =  ( n3341 ) ^ ( rcon )  ;
assign n3343 = in[95:88] ;
assign n3344 =  ( n3342 ) ^ ( n3343 )  ;
assign n3345 =  ( n3344 ) ^ ( n1026 )  ;
assign n3346 =  { ( n3340 ) , ( n3345 ) }  ;
assign n3347 = in[119:112] ;
assign n3348 = in[87:80] ;
assign n3349 =  ( n3347 ) ^ ( n3348 )  ;
assign n3350 =  ( n3349 ) ^ ( n1796 )  ;
assign n3351 =  { ( n3346 ) , ( n3350 ) }  ;
assign n3352 = in[111:104] ;
assign n3353 = in[79:72] ;
assign n3354 =  ( n3352 ) ^ ( n3353 )  ;
assign n3355 =  ( n3354 ) ^ ( n2567 )  ;
assign n3356 =  { ( n3351 ) , ( n3355 ) }  ;
assign n3357 = in[103:96] ;
assign n3358 = in[71:64] ;
assign n3359 =  ( n3357 ) ^ ( n3358 )  ;
assign n3360 =  ( n3359 ) ^ ( n3338 )  ;
assign n3361 =  { ( n3356 ) , ( n3360 ) }  ;
assign n3362 = in[127:120] ;
assign n3363 =  ( n3362 ) ^ ( rcon )  ;
assign n3364 = in[95:88] ;
assign n3365 =  ( n3363 ) ^ ( n3364 )  ;
assign n3366 = in[63:56] ;
assign n3367 =  ( n3365 ) ^ ( n3366 )  ;
assign n3368 =  ( n3367 ) ^ ( n1026 )  ;
assign n3369 =  { ( n3361 ) , ( n3368 ) }  ;
assign n3370 = in[119:112] ;
assign n3371 = in[87:80] ;
assign n3372 =  ( n3370 ) ^ ( n3371 )  ;
assign n3373 = in[55:48] ;
assign n3374 =  ( n3372 ) ^ ( n3373 )  ;
assign n3375 =  ( n3374 ) ^ ( n1796 )  ;
assign n3376 =  { ( n3369 ) , ( n3375 ) }  ;
assign n3377 = in[111:104] ;
assign n3378 = in[79:72] ;
assign n3379 =  ( n3377 ) ^ ( n3378 )  ;
assign n3380 = in[47:40] ;
assign n3381 =  ( n3379 ) ^ ( n3380 )  ;
assign n3382 =  ( n3381 ) ^ ( n2567 )  ;
assign n3383 =  { ( n3376 ) , ( n3382 ) }  ;
assign n3384 = in[103:96] ;
assign n3385 = in[71:64] ;
assign n3386 =  ( n3384 ) ^ ( n3385 )  ;
assign n3387 = in[39:32] ;
assign n3388 =  ( n3386 ) ^ ( n3387 )  ;
assign n3389 =  ( n3388 ) ^ ( n3338 )  ;
assign n3390 =  { ( n3383 ) , ( n3389 ) }  ;
assign n3391 = in[127:120] ;
assign n3392 =  ( n3391 ) ^ ( rcon )  ;
assign n3393 = in[95:88] ;
assign n3394 =  ( n3392 ) ^ ( n3393 )  ;
assign n3395 = in[63:56] ;
assign n3396 =  ( n3394 ) ^ ( n3395 )  ;
assign n3397 = in[31:24] ;
assign n3398 =  ( n3396 ) ^ ( n3397 )  ;
assign n3399 =  ( n3398 ) ^ ( n1026 )  ;
assign n3400 =  { ( n3390 ) , ( n3399 ) }  ;
assign n3401 = in[119:112] ;
assign n3402 = in[87:80] ;
assign n3403 =  ( n3401 ) ^ ( n3402 )  ;
assign n3404 = in[55:48] ;
assign n3405 =  ( n3403 ) ^ ( n3404 )  ;
assign n3406 = in[23:16] ;
assign n3407 =  ( n3405 ) ^ ( n3406 )  ;
assign n3408 =  ( n3407 ) ^ ( n1796 )  ;
assign n3409 =  { ( n3400 ) , ( n3408 ) }  ;
assign n3410 = in[111:104] ;
assign n3411 = in[79:72] ;
assign n3412 =  ( n3410 ) ^ ( n3411 )  ;
assign n3413 = in[47:40] ;
assign n3414 =  ( n3412 ) ^ ( n3413 )  ;
assign n3415 = in[15:8] ;
assign n3416 =  ( n3414 ) ^ ( n3415 )  ;
assign n3417 =  ( n3416 ) ^ ( n2567 )  ;
assign n3418 =  { ( n3409 ) , ( n3417 ) }  ;
assign n3419 = in[103:96] ;
assign n3420 = in[71:64] ;
assign n3421 =  ( n3419 ) ^ ( n3420 )  ;
assign n3422 = in[39:32] ;
assign n3423 =  ( n3421 ) ^ ( n3422 )  ;
assign n3424 = in[7:0] ;
assign n3425 =  ( n3423 ) ^ ( n3424 )  ;
assign n3426 =  ( n3425 ) ^ ( n3338 )  ;
assign n3427 =  { ( n3418 ) , ( n3426 ) }  ;
always @(posedge clk) begin
   if(rst) begin
       in <= in_randinit ;
       rcon <= rcon_randinit ;
       out_1 <= out_1_randinit ;
       __COUNTER_start__n0 <= 0;
   end
   else if(__START__ && __ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           in <= in ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           rcon <= rcon ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           out_1 <= n3427 ;
       end
   end
end
endmodule
