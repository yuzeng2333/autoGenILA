module SDP_C_chn_out_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:318" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_c.v:319" *)
  output outsig;
  assign outsig = in_0;
endmodule
