module \$paramod\SDP_X_mgc_in_wire_v1\rscid=16\width=16 (d, z);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:109" *)
  output [15:0] d;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_x.v:110" *)
  input [15:0] z;
  assign d = z;
endmodule
