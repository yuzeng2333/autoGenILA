module top(clk_i, rst_i, mem_d_data_rd_i, mem_d_accept_i, mem_d_ack_i, mem_d_error_i, mem_d_resp_tag_i, mem_i_accept_i, mem_i_valid_i, mem_i_error_i, mem_i_inst_i, intr_i, reset_vector_i, cpu_id_i, mem_d_addr_o_fifo, mem_d_data_wr_o_fifo, mem_d_rd_o_fifo, mem_d_wr_o_fifo, mem_d_cacheable_o_fifo, mem_d_req_tag_o_fifo, mem_d_invalidate_o_fifo, mem_d_writeback_o_fifo, mem_d_flush_o_fifo, mem_i_rd_o_fifo, mem_i_flush_o_fifo, mem_i_invalidate_o_fifo, mem_i_pc_o_fifo);
  wire _0000_;
  wire _0001_;
  wire _0002_;
  wire _0003_;
  wire _0004_;
  wire _0005_;
  wire [31:0] _0006_;
  wire [31:0] _0007_;
  wire [31:0] _0008_;
  wire [31:0] _0009_;
  wire [31:0] _0010_;
  wire [31:0] _0011_;
  wire [31:0] _0012_;
  wire [31:0] _0013_;
  wire _0014_;
  wire _0015_;
  wire _0016_;
  wire _0017_;
  wire [3:0] _0018_;
  wire [3:0] _0019_;
  wire [3:0] _0020_;
  wire [3:0] _0021_;
  wire [31:0] _0022_;
  wire [31:0] _0023_;
  wire [31:0] _0024_;
  wire [31:0] _0025_;
  wire _0026_;
  wire _0027_;
  wire _0028_;
  wire _0029_;
  wire _0030_;
  wire [31:0] _0031_;
  wire [31:0] _0032_;
  wire [5:0] _0033_;
  wire [31:0] _0034_;
  wire _0035_;
  wire _0036_;
  wire _0037_;
  wire [5:0] _0038_;
  wire [31:0] _0039_;
  wire [31:0] _0040_;
  wire [31:0] _0041_;
  wire [31:0] _0042_;
  wire [31:0] _0043_;
  wire _0044_;
  wire _0045_;
  wire _0046_;
  wire _0047_;
  wire _0048_;
  wire _0049_;
  wire _0050_;
  wire _0051_;
  wire _0052_;
  wire _0053_;
  wire _0054_;
  wire _0055_;
  wire _0056_;
  wire _0057_;
  wire _0058_;
  wire _0059_;
  wire _0060_;
  wire _0061_;
  wire _0062_;
  wire _0063_;
  wire [31:0] _0064_;
  wire _0065_;
  wire _0066_;
  wire _0067_;
  wire _0068_;
  wire _0069_;
  wire _0070_;
  wire _0071_;
  wire _0072_;
  wire [31:0] _0073_;
  wire _0074_;
  wire [31:0] _0075_;
  wire [5:0] _0076_;
  wire [5:0] _0077_;
  wire [5:0] _0078_;
  wire [5:0] _0079_;
  wire [5:0] _0080_;
  wire [5:0] _0081_;
  wire [31:0] _0082_;
  wire [31:0] _0083_;
  wire _0084_;
  wire [31:0] _0085_;
  wire [31:0] _0086_;
  wire [31:0] _0087_;
  wire [31:0] _0088_;
  wire _0089_;
  wire [31:0] _0090_;
  wire [31:0] _0091_;
  wire [31:0] _0092_;
  wire [31:0] _0093_;
  wire [31:0] _0094_;
  wire [31:0] _0095_;
  wire _0096_;
  wire [31:0] _0097_;
  wire _0098_;
  wire [31:0] _0099_;
  wire [31:0] _0100_;
  wire [31:0] _0101_;
  wire [31:0] _0102_;
  wire [1:0] _0103_;
  wire _0104_;
  wire [1:0] _0105_;
  wire [1:0] _0106_;
  wire [31:0] _0107_;
  wire [31:0] _0108_;
  wire [31:0] _0109_;
  wire _0110_;
  wire _0111_;
  wire [31:0] _0112_;
  wire [31:0] _0113_;
  wire [31:0] _0114_;
  wire [31:0] _0115_;
  wire [31:0] _0116_;
  wire [31:0] _0117_;
  wire _0118_;
  wire [31:0] _0119_;
  wire [31:0] _0120_;
  wire [31:0] _0121_;
  wire _0122_;
  wire [31:0] _0123_;
  wire [31:0] _0124_;
  wire [31:0] _0125_;
  wire [31:0] _0126_;
  wire [31:0] _0127_;
  wire [31:0] _0128_;
  wire _0129_;
  wire [31:0] _0130_;
  wire [31:0] _0131_;
  wire [31:0] _0132_;
  wire _0133_;
  wire _0134_;
  wire [31:0] _0135_;
  wire [31:0] _0136_;
  wire [31:0] _0137_;
  wire _0138_;
  wire [31:0] _0139_;
  wire _0140_;
  wire [31:0] _0141_;
  wire [31:0] _0142_;
  wire [31:0] _0143_;
  wire [31:0] _0144_;
  wire _0145_;
  wire [31:0] _0146_;
  wire [31:0] _0147_;
  wire [1:0] _0148_;
  wire _0149_;
  wire [31:0] _0150_;
  wire [31:0] _0151_;
  wire [31:0] _0152_;
  wire [31:0] _0153_;
  wire [1:0] _0154_;
  wire [31:0] _0155_;
  wire [31:0] _0156_;
  wire [31:0] _0157_;
  wire _0158_;
  wire [31:0] _0159_;
  wire _0160_;
  wire [31:0] _0161_;
  wire [31:0] _0162_;
  wire [31:0] _0163_;
  wire [31:0] _0164_;
  wire [31:0] _0165_;
  wire [31:0] _0166_;
  wire [31:0] _0167_;
  wire [31:0] _0168_;
  wire [31:0] _0169_;
  wire [5:0] _0170_;
  wire [31:0] _0171_;
  wire [31:0] _0172_;
  wire [31:0] _0173_;
  wire [31:0] _0174_;
  wire [31:0] _0175_;
  wire [31:0] _0176_;
  wire [31:0] _0177_;
  wire [31:0] _0178_;
  wire _0179_;
  wire _0180_;
  wire _0181_;
  wire _0182_;
  wire _0183_;
  wire _0184_;
  wire _0185_;
  wire _0186_;
  wire _0187_;
  wire _0188_;
  wire _0189_;
  wire _0190_;
  wire _0191_;
  wire _0192_;
  wire _0193_;
  wire _0194_;
  wire _0195_;
  wire _0196_;
  wire _0197_;
  wire [31:0] _0198_;
  wire [31:0] _0199_;
  wire [31:0] _0200_;
  wire _0201_;
  wire _0202_;
  wire _0203_;
  wire _0204_;
  wire _0205_;
  wire _0206_;
  wire _0207_;
  wire _0208_;
  wire _0209_;
  wire _0210_;
  wire [6:0] _0211_;
  wire _0212_;
  wire [2:0] _0213_;
  wire _0214_;
  wire _0215_;
  wire _0216_;
  wire _0217_;
  wire [1:0] _0218_;
  wire _0219_;
  wire _0220_;
  wire _0221_;
  wire _0222_;
  wire _0223_;
  wire _0224_;
  wire _0225_;
  wire _0226_;
  wire _0227_;
  wire _0228_;
  wire [1:0] _0229_;
  wire _0230_;
  wire _0231_;
  wire [31:0] _0232_;
  wire [31:0] _0233_;
  wire [31:0] _0234_;
  wire [31:0] _0235_;
  wire [31:0] _0236_;
  wire [31:0] _0237_;
  wire [31:0] _0238_;
  wire [31:0] _0239_;
  wire [31:0] _0240_;
  wire [31:0] _0241_;
  wire _0242_;
  wire _0243_;
  wire _0244_;
  wire _0245_;
  wire _0246_;
  wire _0247_;
  wire _0248_;
  wire _0249_;
  wire _0250_;
  wire _0251_;
  wire _0252_;
  wire _0253_;
  wire _0254_;
  wire _0255_;
  wire _0256_;
  wire _0257_;
  wire _0258_;
  wire _0259_;
  wire _0260_;
  wire _0261_;
  wire _0262_;
  wire _0263_;
  wire _0264_;
  wire _0265_;
  wire _0266_;
  wire _0267_;
  wire _0268_;
  wire _0269_;
  wire _0270_;
  wire _0271_;
  wire _0272_;
  wire _0273_;
  wire _0274_;
  wire _0275_;
  wire _0276_;
  wire _0277_;
  wire _0278_;
  wire _0279_;
  wire _0280_;
  wire _0281_;
  wire _0282_;
  wire _0283_;
  wire _0284_;
  wire _0285_;
  wire _0286_;
  wire _0287_;
  wire _0288_;
  wire _0289_;
  wire _0290_;
  wire _0291_;
  wire _0292_;
  wire _0293_;
  wire _0294_;
  wire _0295_;
  wire _0296_;
  wire _0297_;
  wire _0298_;
  wire _0299_;
  wire _0300_;
  wire _0301_;
  wire _0302_;
  wire _0303_;
  wire _0304_;
  wire _0305_;
  wire _0306_;
  wire _0307_;
  wire _0308_;
  wire _0309_;
  wire _0310_;
  wire _0311_;
  wire _0312_;
  wire _0313_;
  wire _0314_;
  wire _0315_;
  wire _0316_;
  wire _0317_;
  wire _0318_;
  wire _0319_;
  wire _0320_;
  wire _0321_;
  wire _0322_;
  wire _0323_;
  wire _0324_;
  wire _0325_;
  wire _0326_;
  wire _0327_;
  wire _0328_;
  wire _0329_;
  wire _0330_;
  wire _0331_;
  wire _0332_;
  wire _0333_;
  wire _0334_;
  wire _0335_;
  wire _0336_;
  wire _0337_;
  wire _0338_;
  wire _0339_;
  wire _0340_;
  wire _0341_;
  wire _0342_;
  wire _0343_;
  wire _0344_;
  wire _0345_;
  wire _0346_;
  wire _0347_;
  wire _0348_;
  wire _0349_;
  wire _0350_;
  wire _0351_;
  wire _0352_;
  wire _0353_;
  wire _0354_;
  wire _0355_;
  wire _0356_;
  wire _0357_;
  wire _0358_;
  wire _0359_;
  wire _0360_;
  wire _0361_;
  wire _0362_;
  wire _0363_;
  wire _0364_;
  wire _0365_;
  wire _0366_;
  wire _0367_;
  wire _0368_;
  wire _0369_;
  wire _0370_;
  wire _0371_;
  wire _0372_;
  wire _0373_;
  wire _0374_;
  wire _0375_;
  wire _0376_;
  wire _0377_;
  wire _0378_;
  wire _0379_;
  wire _0380_;
  wire _0381_;
  wire _0382_;
  wire _0383_;
  wire _0384_;
  wire _0385_;
  wire _0386_;
  wire _0387_;
  wire _0388_;
  wire _0389_;
  wire _0390_;
  wire _0391_;
  wire _0392_;
  wire _0393_;
  wire _0394_;
  wire _0395_;
  wire _0396_;
  wire _0397_;
  wire _0398_;
  wire _0399_;
  wire _0400_;
  wire _0401_;
  wire _0402_;
  wire _0403_;
  wire _0404_;
  wire _0405_;
  wire _0406_;
  wire _0407_;
  wire _0408_;
  wire _0409_;
  wire _0410_;
  wire _0411_;
  wire _0412_;
  wire _0413_;
  wire _0414_;
  wire _0415_;
  wire _0416_;
  wire _0417_;
  wire _0418_;
  wire _0419_;
  wire _0420_;
  wire _0421_;
  wire _0422_;
  wire _0423_;
  wire _0424_;
  wire _0425_;
  wire _0426_;
  wire _0427_;
  wire _0428_;
  wire _0429_;
  wire _0430_;
  wire _0431_;
  wire _0432_;
  wire _0433_;
  wire _0434_;
  wire _0435_;
  wire _0436_;
  wire _0437_;
  wire _0438_;
  wire _0439_;
  wire _0440_;
  wire [31:0] _0441_;
  wire [62:0] _0442_;
  wire _0443_;
  wire [31:0] _0444_;
  wire [31:0] _0445_;
  wire _0446_;
  wire [31:0] _0447_;
  wire [31:0] _0448_;
  wire _0449_;
  wire _0450_;
  wire _0451_;
  wire _0452_;
  wire _0453_;
  wire _0454_;
  wire _0455_;
  wire _0456_;
  wire _0457_;
  wire _0458_;
  wire _0459_;
  wire _0460_;
  wire _0461_;
  wire _0462_;
  wire [31:0] _0463_;
  wire [31:0] _0464_;
  wire [31:0] _0465_;
  wire [31:0] _0466_;
  wire [31:0] _0467_;
  wire [31:0] _0468_;
  wire _0469_;
  wire _0470_;
  wire _0471_;
  wire _0472_;
  wire [31:0] _0473_;
  wire [31:0] _0474_;
  wire [31:0] _0475_;
  wire [31:0] _0476_;
  wire [31:0] _0477_;
  wire [31:0] _0478_;
  wire [31:0] _0479_;
  wire [62:0] _0480_;
  wire [62:0] _0481_;
  wire [62:0] _0482_;
  wire [62:0] _0483_;
  wire [31:0] _0484_;
  wire [31:0] _0485_;
  wire [31:0] _0486_;
  wire [31:0] _0487_;
  wire [31:0] _0488_;
  wire _0489_;
  wire _0490_;
  wire [31:0] _0491_;
  wire [31:0] _0492_;
  wire [31:0] _0493_;
  wire [31:0] _0494_;
  wire [3:0] _0495_;
  wire [31:0] _0496_;
  wire [31:0] _0497_;
  wire [3:0] _0498_;
  wire [31:0] _0499_;
  wire [31:0] _0500_;
  wire [3:0] _0501_;
  wire [31:0] _0502_;
  wire [31:0] _0503_;
  wire [3:0] _0504_;
  wire [31:0] _0505_;
  wire [31:0] _0506_;
  wire [3:0] _0507_;
  wire [31:0] _0508_;
  wire [31:0] _0509_;
  wire [3:0] _0510_;
  wire [31:0] _0511_;
  wire [31:0] _0512_;
  wire [3:0] _0513_;
  wire [31:0] _0514_;
  wire [31:0] _0515_;
  wire [2:0] _0516_;
  wire [31:0] _0517_;
  wire [31:0] _0518_;
  wire [2:0] _0519_;
  wire [31:0] _0520_;
  wire [31:0] _0521_;
  wire [2:0] _0522_;
  wire [31:0] _0523_;
  wire [31:0] _0524_;
  wire [2:0] _0525_;
  wire [31:0] _0526_;
  wire [31:0] _0527_;
  wire [2:0] _0528_;
  wire [31:0] _0529_;
  wire [31:0] _0530_;
  wire [2:0] _0531_;
  wire [31:0] _0532_;
  wire [3:0] _0533_;
  wire [31:0] _0534_;
  wire [31:0] _0535_;
  wire _0536_;
  wire _0537_;
  wire [31:0] _0538_;
  wire [3:0] _0539_;
  wire [31:0] _0540_;
  wire [31:0] _0541_;
  wire _0542_;
  wire _0543_;
  wire [3:0] _0544_;
  wire [31:0] _0545_;
  wire [31:0] _0546_;
  wire _0547_;
  wire _0548_;
  wire [3:0] _0549_;
  wire [31:0] _0550_;
  wire [31:0] _0551_;
  wire _0552_;
  wire _0553_;
  wire [3:0] _0554_;
  wire [31:0] _0555_;
  wire [31:0] _0556_;
  wire _0557_;
  wire _0558_;
  wire _0559_;
  wire [3:0] _0560_;
  wire [31:0] _0561_;
  wire [31:0] _0562_;
  wire _0563_;
  wire _0564_;
  wire _0565_;
  wire [3:0] _0566_;
  wire [31:0] _0567_;
  wire [31:0] _0568_;
  wire _0569_;
  wire _0570_;
  wire [3:0] _0571_;
  wire [31:0] _0572_;
  wire [31:0] _0573_;
  wire [31:0] _0574_;
  wire [31:0] _0575_;
  wire [31:0] _0576_;
  wire [31:0] _0577_;
  wire [31:0] _0578_;
  wire [31:0] _0579_;
  wire [31:0] _0580_;
  wire _0581_;
  wire _0582_;
  wire _0583_;
  wire _0584_;
  wire _0585_;
  wire _0586_;
  wire _0587_;
  wire _0588_;
  wire _0589_;
  wire _0590_;
  wire _0591_;
  wire _0592_;
  wire _0593_;
  wire _0594_;
  wire _0595_;
  wire _0596_;
  wire _0597_;
  wire _0598_;
  wire _0599_;
  wire _0600_;
  wire _0601_;
  wire _0602_;
  wire _0603_;
  wire _0604_;
  wire _0605_;
  wire _0606_;
  wire _0607_;
  wire _0608_;
  wire _0609_;
  wire _0610_;
  wire _0611_;
  wire _0612_;
  wire _0613_;
  wire _0614_;
  wire _0615_;
  wire _0616_;
  wire _0617_;
  wire _0618_;
  wire _0619_;
  wire _0620_;
  wire _0621_;
  wire _0622_;
  wire _0623_;
  wire [31:0] _0624_;
  wire [31:0] _0625_;
  wire [31:0] _0626_;
  wire [31:0] _0627_;
  wire [31:0] _0628_;
  wire [31:0] _0629_;
  wire [31:0] _0630_;
  wire [31:0] _0631_;
  wire [31:0] _0632_;
  wire [31:0] _0633_;
  wire [31:0] _0634_;
  wire [31:0] _0635_;
  wire [15:0] _0636_;
  wire [31:0] _0637_;
  wire _0638_;
  wire [31:0] _0639_;
  wire [31:0] _0640_;
  wire [31:0] _0641_;
  wire _0642_;
  wire _0643_;
  wire _0644_;
  wire _0645_;
  wire [31:0] _0646_;
  wire _0647_;
  wire [1:0] _0648_;
  wire _0649_;
  wire _0650_;
  wire _0651_;
  wire _0652_;
  wire _0653_;
  wire _0654_;
  wire _0655_;
  wire _0656_;
  wire [31:0] _0657_;
  wire [31:0] _0658_;
  wire [31:0] _0659_;
  wire _0660_;
  wire _0661_;
  wire [31:0] _0662_;
  wire _0663_;
  wire _0664_;
  wire [31:0] _0665_;
  wire [31:0] _0666_;
  wire [65:0] _0667_;
  wire _0668_;
  wire [31:0] _0669_;
  wire _0670_;
  wire _0671_;
  wire _0672_;
  wire _0673_;
  wire _0674_;
  wire _0675_;
  wire _0676_;
  wire _0677_;
  wire _0678_;
  wire _0679_;
  wire _0680_;
  wire _0681_;
  wire _0682_;
  wire [65:0] _0683_;
  wire [31:0] _0684_;
  wire _0685_;
  wire _0686_;
  wire [31:0] _0687_;
  wire [31:0] _0688_;
  wire _0689_;
  wire _0690_;
  wire _0691_;
  wire [31:0] _0692_;
  wire [31:0] _0693_;
  wire _0694_;
  wire _0695_;
  wire _0696_;
  wire _0697_;
  wire [31:0] _0698_;
  wire [31:0] _0699_;
  wire [31:0] _0700_;
  wire [31:0] _0701_;
  wire [31:0] _0702_;
  wire _0703_;
  wire [31:0] _0704_;
  wire [31:0] _0705_;
  wire [31:0] _0706_;
  wire [31:0] _0707_;
  wire _0708_;
  wire [5:0] _0709_;
  wire _0710_;
  wire _0711_;
  wire _0712_;
  wire _0713_;
  wire _0714_;
  wire _0715_;
  wire _0716_;
  wire _0717_;
  wire _0718_;
  wire _0719_;
  wire _0720_;
  wire _0721_;
  wire _0722_;
  wire _0723_;
  wire _0724_;
  wire _0725_;
  wire _0726_;
  wire _0727_;
  wire _0728_;
  wire _0729_;
  wire _0730_;
  wire _0731_;
  wire [31:0] _0732_;
  wire _0733_;
  wire _0734_;
  wire _0735_;
  wire [31:0] _0736_;
  wire _0737_;
  wire _0738_;
  wire _0739_;
  wire _0740_;
  wire _0741_;
  wire _0742_;
  wire _0743_;
  wire _0744_;
  wire _0745_;
  wire [31:0] _0746_;
  wire [31:0] _0747_;
  wire [31:0] _0748_;
  wire _0749_;
  wire _0750_;
  wire [9:0] _0751_;
  wire [9:0] _0752_;
  wire [9:0] _0753_;
  wire [5:0] _0754_;
  wire [5:0] _0755_;
  wire [5:0] _0756_;
  wire [31:0] _0757_;
  wire [31:0] _0758_;
  wire [31:0] _0759_;
  wire [31:0] _0760_;
  wire [31:0] _0761_;
  wire [31:0] _0762_;
  wire [31:0] _0763_;
  wire [31:0] _0764_;
  wire _0765_;
  wire _0766_;
  wire _0767_;
  wire _0768_;
  wire [31:0] _0769_;
  wire _0770_;
  wire _0771_;
  wire _0772_;
  wire _0773_;
  wire _0774_;
  wire _0775_;
  wire _0776_;
  wire _0777_;
  wire _0778_;
  wire _0779_;
  wire [9:0] _0780_;
  wire [5:0] _0781_;
  wire _0782_;
  wire _0783_;
  wire _0784_;
  wire _0785_;
  wire _0786_;
  wire _0787_;
  wire _0788_;
  wire _0789_;
  wire _0790_;
  wire _0791_;
  wire _0792_;
  wire _0793_;
  wire _0794_;
  wire _0795_;
  wire _0796_;
  wire _0797_;
  wire _0798_;
  wire _0799_;
  wire _0800_;
  wire _0801_;
  wire _0802_;
  wire _0803_;
  wire _0804_;
  wire _0805_;
  wire _0806_;
  wire _0807_;
  wire _0808_;
  wire _0809_;
  wire _0810_;
  wire [5:0] _0811_;
  wire [5:0] _0812_;
  wire [31:0] _0813_;
  wire [31:0] _0814_;
  wire [31:0] _0815_;
  wire [31:0] _0816_;
  wire [31:0] _0817_;
  wire [31:0] _0818_;
  wire [31:0] _0819_;
  wire [31:0] _0820_;
  wire [31:0] _0821_;
  wire [31:0] _0822_;
  wire _0823_;
  wire _0824_;
  wire [9:0] _0825_;
  wire [9:0] _0826_;
  wire [9:0] _0827_;
  wire _0828_;
  wire [5:0] _0829_;
  wire _0830_;
  wire _0831_;
  wire _0832_;
  wire _0833_;
  wire [5:0] _0834_;
  wire _0835_;
  wire [5:0] _0836_;
  wire [5:0] _0837_;
  wire [5:0] _0838_;
  wire [31:0] _0839_;
  wire [31:0] _0840_;
  wire [31:0] _0841_;
  wire [31:0] _0842_;
  wire [31:0] _0843_;
  wire [31:0] _0844_;
  wire _0845_;
  wire _0846_;
  wire [9:0] _0847_;
  wire [9:0] _0848_;
  wire _0849_;
  wire _0850_;
  wire _0851_;
  wire _0852_;
  wire [31:0] _0853_;
  wire [31:0] _0854_;
  wire [31:0] _0855_;
  wire [31:0] _0856_;
  wire _0857_;
  wire _0858_;
  wire _0859_;
  wire _0860_;
  wire _0861_;
  wire _0862_;
  wire _0863_;
  wire _0864_;
  wire _0865_;
  wire _0866_;
  wire _0867_;
  wire _0868_;
  wire _0869_;
  wire _0870_;
  wire _0871_;
  wire _0872_;
  wire _0873_;
  wire _0874_;
  wire _0875_;
  wire _0876_;
  wire [31:0] _0877_;
  wire [31:0] _0878_;
  wire [31:0] _0879_;
  wire [31:0] _0880_;
  wire _0881_;
  wire [5:0] _0882_;
  wire [5:0] _0883_;
  wire _0884_;
  wire [5:0] _0885_;
  wire [31:0] _0886_;
  wire [31:0] _0887_;
  wire [31:0] _0888_;
  wire [31:0] _0889_;
  wire [31:0] _0890_;
  wire [31:0] _0891_;
  wire [31:0] _0892_;
  wire [31:0] _0893_;
  wire [31:0] _0894_;
  wire [31:0] _0895_;
  wire [31:0] _0896_;
  wire [31:0] _0897_;
  wire [31:0] _0898_;
  wire [31:0] _0899_;
  wire [31:0] _0900_;
  wire [31:0] _0901_;
  wire [31:0] _0902_;
  wire [31:0] _0903_;
  wire [31:0] _0904_;
  wire [31:0] _0905_;
  wire [31:0] _0906_;
  wire [31:0] _0907_;
  wire [31:0] _0908_;
  wire [31:0] _0909_;
  wire [31:0] _0910_;
  wire [31:0] _0911_;
  wire [31:0] _0912_;
  wire [31:0] _0913_;
  wire [31:0] _0914_;
  wire [31:0] _0915_;
  wire [31:0] _0916_;
  wire _0917_;
  wire _0918_;
  wire _0919_;
  wire _0920_;
  wire _0921_;
  wire _0922_;
  wire _0923_;
  wire _0924_;
  wire _0925_;
  wire _0926_;
  wire _0927_;
  wire _0928_;
  wire _0929_;
  wire _0930_;
  wire _0931_;
  wire _0932_;
  wire _0933_;
  wire _0934_;
  wire _0935_;
  wire _0936_;
  wire _0937_;
  wire _0938_;
  wire _0939_;
  wire _0940_;
  wire _0941_;
  wire _0942_;
  wire _0943_;
  wire _0944_;
  wire _0945_;
  wire _0946_;
  wire _0947_;
  wire _0948_;
  wire _0949_;
  wire _0950_;
  wire _0951_;
  wire _0952_;
  wire _0953_;
  wire _0954_;
  wire _0955_;
  wire _0956_;
  wire _0957_;
  wire _0958_;
  wire _0959_;
  wire _0960_;
  wire _0961_;
  wire _0962_;
  wire _0963_;
  wire _0964_;
  wire _0965_;
  wire _0966_;
  wire _0967_;
  wire _0968_;
  wire _0969_;
  wire _0970_;
  wire _0971_;
  wire _0972_;
  wire _0973_;
  wire _0974_;
  wire _0975_;
  wire _0976_;
  wire _0977_;
  wire _0978_;
  wire _0979_;
  wire _0980_;
  wire _0981_;
  wire _0982_;
  wire _0983_;
  wire _0984_;
  wire _0985_;
  wire _0986_;
  wire _0987_;
  wire _0988_;
  wire _0989_;
  wire _0990_;
  wire _0991_;
  wire _0992_;
  wire _0993_;
  wire _0994_;
  wire _0995_;
  wire _0996_;
  wire _0997_;
  wire _0998_;
  wire _0999_;
  wire _1000_;
  wire _1001_;
  wire _1002_;
  wire _1003_;
  wire _1004_;
  wire _1005_;
  wire _1006_;
  wire _1007_;
  wire _1008_;
  wire _1009_;
  wire [31:0] _1010_;
  wire [31:0] _1011_;
  wire [31:0] _1012_;
  wire [31:0] _1013_;
  wire [31:0] _1014_;
  wire [31:0] _1015_;
  wire [31:0] _1016_;
  wire [31:0] _1017_;
  wire [31:0] _1018_;
  wire [31:0] _1019_;
  wire [31:0] _1020_;
  wire [31:0] _1021_;
  wire [31:0] _1022_;
  wire [31:0] _1023_;
  wire [31:0] _1024_;
  wire [31:0] _1025_;
  wire [31:0] _1026_;
  wire [31:0] _1027_;
  wire [31:0] _1028_;
  wire [31:0] _1029_;
  wire [31:0] _1030_;
  wire [31:0] _1031_;
  wire [31:0] _1032_;
  wire [31:0] _1033_;
  wire [31:0] _1034_;
  wire [31:0] _1035_;
  wire [31:0] _1036_;
  wire [31:0] _1037_;
  wire [31:0] _1038_;
  wire [31:0] _1039_;
  wire [31:0] _1040_;
  wire [31:0] _1041_;
  wire [31:0] _1042_;
  wire _1043_;
  wire _1044_;
  wire _1045_;
  wire _1046_;
  wire _1047_;
  wire _1048_;
  wire _1049_;
  wire [3:0] _1050_;
  wire _1051_;
  wire _1052_;
  wire _1053_;
  wire _1054_;
  wire [31:0] _1055_;
  wire [31:0] _1056_;
  wire _1057_;
  wire [3:0] _1058_;
  wire [31:0] _1059_;
  wire [31:0] _1060_;
  wire [3:0] _1061_;
  wire [31:0] _1062_;
  wire [31:0] _1063_;
  wire [3:0] _1064_;
  wire [31:0] _1065_;
  wire [31:0] _1066_;
  wire [3:0] _1067_;
  wire [31:0] _1068_;
  wire [31:0] _1069_;
  wire [31:0] _1070_;
  wire [31:0] _1071_;
  wire [31:0] _1072_;
  wire [31:0] _1073_;
  wire _1074_;
  wire [31:0] _1075_;
  wire _1076_;
  wire _1077_;
  wire _1078_;
  wire [31:0] _1079_;
  wire [5:0] _1080_;
  wire [5:0] _1081_;
  wire [5:0] _1082_;
  wire [5:0] _1083_;
  wire [5:0] _1084_;
  wire _1085_;
  wire _1086_;
  wire _1087_;
  wire _1088_;
  wire _1089_;
  wire _1090_;
  wire _1091_;
  wire _1092_;
  wire _1093_;
  wire _1094_;
  wire _1095_;
  wire _1096_;
  wire _1097_;
  wire _1098_;
  wire _1099_;
  wire _1100_;
  wire _1101_;
  wire _1102_;
  wire _1103_;
  wire _1104_;
  wire _1105_;
  wire _1106_;
  wire _1107_;
  wire _1108_;
  wire _1109_;
  wire _1110_;
  wire _1111_;
  wire _1112_;
  wire _1113_;
  wire _1114_;
  wire _1115_;
  wire _1116_;
  wire _1117_;
  wire _1118_;
  wire _1119_;
  wire _1120_;
  wire _1121_;
  wire _1122_;
  wire _1123_;
  wire _1124_;
  wire _1125_;
  wire _1126_;
  wire _1127_;
  wire _1128_;
  wire _1129_;
  wire _1130_;
  wire _1131_;
  wire _1132_;
  wire _1133_;
  wire _1134_;
  wire _1135_;
  wire _1136_;
  wire _1137_;
  wire [3:0] _1138_;
  wire _1139_;
  wire _1140_;
  wire _1141_;
  wire [31:0] _1142_;
  wire [31:0] _1143_;
  wire [31:0] _1144_;
  wire [31:0] _1145_;
  wire _1146_;
  wire _1147_;
  wire _1148_;
  wire _1149_;
  wire [31:0] _1150_;
  wire [31:0] _1151_;
  wire _1152_;
  wire _1153_;
  wire _1154_;
  wire _1155_;
  wire _1156_;
  wire _1157_;
  wire _1158_;
  wire _1159_;
  wire _1160_;
  wire _1161_;
  wire _1162_;
  wire _1163_;
  wire _1164_;
  wire _1165_;
  wire _1166_;
  wire _1167_;
  wire _1168_;
  wire _1169_;
  wire _1170_;
  wire _1171_;
  wire _1172_;
  wire _1173_;
  wire _1174_;
  wire _1175_;
  wire [3:0] _1176_;
  wire [3:0] _1177_;
  wire [3:0] _1178_;
  wire _1179_;
  wire _1180_;
  wire _1181_;
  wire [31:0] _1182_;
  wire [31:0] _1183_;
  wire [31:0] _1184_;
  wire [31:0] _1185_;
  wire [31:0] _1186_;
  wire [31:0] _1187_;
  wire _1188_;
  wire _1189_;
  wire _1190_;
  wire _1191_;
  wire _1192_;
  wire _1193_;
  wire _1194_;
  wire _1195_;
  wire [35:0] _1196_;
  wire _1197_;
  wire [35:0] _1198_;
  wire [35:0] _1199_;
  wire [1:0] _1200_;
  wire _1201_;
  wire _1202_;
  wire _1203_;
  wire [31:0] _1204_;
  wire [31:0] _1205_;
  wire _1206_;
  wire _1207_;
  wire _1208_;
  wire _1209_;
  wire _1210_;
  wire _1211_;
  wire [35:0] _1212_;
  wire [35:0] _1213_;
  wire _1214_;
  wire [1:0] _1215_;
  wire [1:0] _1216_;
  wire _1217_;
  wire _1218_;
  wire [31:0] _1219_;
  wire _1220_;
  wire [32:0] _1221_;
  wire [32:0] _1222_;
  wire [31:0] _1223_;
  wire [32:0] _1224_;
  wire [32:0] _1225_;
  wire [31:0] _1226_;
  wire _1227_;
  wire _1228_;
  wire _1229_;
  wire _1230_;
  wire _1231_;
  wire _1232_;
  wire _1233_;
  wire _1234_;
  wire [31:0] _1235_;
  wire _1236_;
  wire _1237_;
  wire [32:0] _1238_;
  wire [32:0] _1239_;
  wire [32:0] _1240_;
  wire [32:0] _1241_;
  wire _1242_;
  wire _1243_;
  wire _1244_;
  wire _1245_;
  wire _1246_;
  wire _1247_;
  wire [35:0] _1248_;
  wire [35:0] _1249_;
  wire [35:0] _1250_;
  wire [35:0] _1251_;
  wire [35:0] _1252_;
  wire [35:0] _1253_;
  input clk_i;
  input [31:0] cpu_id_i;
  wire \fifo_d_addr.clk ;
  wire [31:0] \fifo_d_addr.in ;
  wire [31:0] \fifo_d_addr.out ;
  reg [31:0] \fifo_d_addr.r0 ;
  reg [31:0] \fifo_d_addr.r1 ;
  wire \fifo_d_addr.rst ;
  wire \fifo_d_addr.wr ;
  wire \fifo_d_data_wr.clk ;
  wire [31:0] \fifo_d_data_wr.in ;
  wire [31:0] \fifo_d_data_wr.out ;
  reg [31:0] \fifo_d_data_wr.r0 ;
  reg [31:0] \fifo_d_data_wr.r1 ;
  wire \fifo_d_data_wr.rst ;
  wire \fifo_d_data_wr.wr ;
  wire \fifo_d_rd.clk ;
  wire \fifo_d_rd.in ;
  wire \fifo_d_rd.out ;
  reg \fifo_d_rd.r0 ;
  reg \fifo_d_rd.r1 ;
  wire \fifo_d_rd.rst ;
  wire \fifo_d_rd.wr ;
  wire \fifo_d_wr.clk ;
  wire [3:0] \fifo_d_wr.in ;
  wire [3:0] \fifo_d_wr.out ;
  reg [3:0] \fifo_d_wr.r0 ;
  reg [3:0] \fifo_d_wr.r1 ;
  wire \fifo_d_wr.rst ;
  wire \fifo_d_wr.wr ;
  wire \fifo_i_pc.clk ;
  wire [31:0] \fifo_i_pc.in ;
  wire [31:0] \fifo_i_pc.out ;
  reg [31:0] \fifo_i_pc.r0 ;
  reg [31:0] \fifo_i_pc.r1 ;
  wire \fifo_i_pc.rst ;
  wire \fifo_i_pc.wr ;
  wire \fifo_i_rd.clk ;
  wire \fifo_i_rd.in ;
  wire \fifo_i_rd.out ;
  reg \fifo_i_rd.r0 ;
  reg \fifo_i_rd.r1 ;
  wire \fifo_i_rd.rst ;
  wire \fifo_i_rd.wr ;
  input intr_i;
  input mem_d_accept_i;
  input mem_d_ack_i;
  wire mem_d_addr_o;
  output [31:0] mem_d_addr_o_fifo;
  wire mem_d_cacheable_o;
  output mem_d_cacheable_o_fifo;
  input [31:0] mem_d_data_rd_i;
  wire mem_d_data_wr_o;
  output [31:0] mem_d_data_wr_o_fifo;
  input mem_d_error_i;
  wire mem_d_flush_o;
  output mem_d_flush_o_fifo;
  wire mem_d_invalidate_o;
  output mem_d_invalidate_o_fifo;
  wire mem_d_rd_o;
  output mem_d_rd_o_fifo;
  wire mem_d_req_tag_o;
  output [10:0] mem_d_req_tag_o_fifo;
  input [10:0] mem_d_resp_tag_i;
  wire mem_d_wr_o;
  output [3:0] mem_d_wr_o_fifo;
  wire mem_d_writeback_o;
  output mem_d_writeback_o_fifo;
  input mem_i_accept_i;
  input mem_i_error_i;
  wire mem_i_flush_o;
  output mem_i_flush_o_fifo;
  input [31:0] mem_i_inst_i;
  wire mem_i_invalidate_o;
  output mem_i_invalidate_o_fifo;
  wire mem_i_pc_o;
  output [31:0] mem_i_pc_o_fifo;
  wire mem_i_rd_o;
  output mem_i_rd_o_fifo;
  input mem_i_valid_i;
  input [31:0] reset_vector_i;
  input rst_i;
  wire [31:0] \u0.branch_csr_pc_w ;
  wire \u0.branch_csr_request_w ;
  wire [31:0] \u0.branch_d_exec_pc_w ;
  wire [1:0] \u0.branch_d_exec_priv_w ;
  wire \u0.branch_d_exec_request_w ;
  wire [31:0] \u0.branch_pc_w ;
  wire \u0.branch_request_w ;
  wire \u0.clk_i ;
  wire [31:0] \u0.cpu_id_i ;
  wire \u0.csr_opcode_invalid_w ;
  wire [31:0] \u0.csr_opcode_opcode_w ;
  wire [31:0] \u0.csr_opcode_pc_w ;
  wire [4:0] \u0.csr_opcode_ra_idx_w ;
  wire [31:0] \u0.csr_opcode_ra_operand_w ;
  wire [4:0] \u0.csr_opcode_rb_idx_w ;
  wire [31:0] \u0.csr_opcode_rb_operand_w ;
  wire [4:0] \u0.csr_opcode_rd_idx_w ;
  wire \u0.csr_opcode_valid_w ;
  wire [5:0] \u0.csr_result_e1_exception_w ;
  wire [31:0] \u0.csr_result_e1_value_w ;
  wire [31:0] \u0.csr_result_e1_wdata_w ;
  wire \u0.csr_result_e1_write_w ;
  wire [31:0] \u0.csr_writeback_exception_addr_w ;
  wire [31:0] \u0.csr_writeback_exception_pc_w ;
  wire [5:0] \u0.csr_writeback_exception_w ;
  wire [11:0] \u0.csr_writeback_waddr_w ;
  wire [31:0] \u0.csr_writeback_wdata_w ;
  wire \u0.csr_writeback_write_w ;
  wire \u0.div_opcode_valid_w ;
  wire \u0.exec_hold_w ;
  wire \u0.exec_opcode_valid_w ;
  wire \u0.fetch_accept_w ;
  wire \u0.fetch_dec_accept_w ;
  wire \u0.fetch_dec_fault_fetch_w ;
  wire \u0.fetch_dec_fault_page_w ;
  wire [31:0] \u0.fetch_dec_instr_w ;
  wire [31:0] \u0.fetch_dec_pc_w ;
  wire \u0.fetch_dec_valid_w ;
  wire \u0.fetch_fault_fetch_w ;
  wire \u0.fetch_fault_page_w ;
  wire \u0.fetch_in_fault_w ;
  wire \u0.fetch_instr_branch_w ;
  wire \u0.fetch_instr_csr_w ;
  wire \u0.fetch_instr_div_w ;
  wire \u0.fetch_instr_exec_w ;
  wire \u0.fetch_instr_invalid_w ;
  wire \u0.fetch_instr_lsu_w ;
  wire \u0.fetch_instr_mul_w ;
  wire \u0.fetch_instr_rd_valid_w ;
  wire [31:0] \u0.fetch_instr_w ;
  wire [31:0] \u0.fetch_pc_w ;
  wire \u0.fetch_valid_w ;
  wire \u0.ifence_w ;
  wire \u0.interrupt_inhibit_w ;
  wire \u0.intr_i ;
  wire \u0.lsu_opcode_invalid_w ;
  wire [31:0] \u0.lsu_opcode_opcode_w ;
  wire [31:0] \u0.lsu_opcode_pc_w ;
  wire [4:0] \u0.lsu_opcode_ra_idx_w ;
  wire [31:0] \u0.lsu_opcode_ra_operand_w ;
  wire [4:0] \u0.lsu_opcode_rb_idx_w ;
  wire [31:0] \u0.lsu_opcode_rb_operand_w ;
  wire [4:0] \u0.lsu_opcode_rd_idx_w ;
  wire \u0.lsu_opcode_valid_w ;
  wire \u0.lsu_stall_w ;
  wire \u0.mem_d_accept_i ;
  wire \u0.mem_d_ack_i ;
  wire [31:0] \u0.mem_d_addr_o ;
  wire \u0.mem_d_cacheable_o ;
  wire [31:0] \u0.mem_d_data_rd_i ;
  wire [31:0] \u0.mem_d_data_wr_o ;
  wire \u0.mem_d_error_i ;
  wire \u0.mem_d_flush_o ;
  wire \u0.mem_d_invalidate_o ;
  wire \u0.mem_d_rd_o ;
  wire [10:0] \u0.mem_d_req_tag_o ;
  wire [10:0] \u0.mem_d_resp_tag_i ;
  wire [3:0] \u0.mem_d_wr_o ;
  wire \u0.mem_d_writeback_o ;
  wire \u0.mem_i_accept_i ;
  wire \u0.mem_i_error_i ;
  wire \u0.mem_i_flush_o ;
  wire [31:0] \u0.mem_i_inst_i ;
  wire \u0.mem_i_invalidate_o ;
  wire [31:0] \u0.mem_i_pc_o ;
  wire \u0.mem_i_rd_o ;
  wire \u0.mem_i_valid_i ;
  wire \u0.mmu_ifetch_accept_w ;
  wire \u0.mmu_ifetch_error_w ;
  wire \u0.mmu_ifetch_flush_w ;
  wire [31:0] \u0.mmu_ifetch_inst_w ;
  wire \u0.mmu_ifetch_invalidate_w ;
  wire [31:0] \u0.mmu_ifetch_pc_w ;
  wire \u0.mmu_ifetch_rd_w ;
  wire \u0.mmu_ifetch_valid_w ;
  wire \u0.mmu_load_fault_w ;
  wire \u0.mmu_lsu_accept_w ;
  wire \u0.mmu_lsu_ack_w ;
  wire [31:0] \u0.mmu_lsu_addr_w ;
  wire \u0.mmu_lsu_cacheable_w ;
  wire [31:0] \u0.mmu_lsu_data_rd_w ;
  wire [31:0] \u0.mmu_lsu_data_wr_w ;
  wire \u0.mmu_lsu_error_w ;
  wire \u0.mmu_lsu_flush_w ;
  wire \u0.mmu_lsu_invalidate_w ;
  wire \u0.mmu_lsu_rd_w ;
  wire [10:0] \u0.mmu_lsu_req_tag_w ;
  wire [10:0] \u0.mmu_lsu_resp_tag_w ;
  wire [3:0] \u0.mmu_lsu_wr_w ;
  wire \u0.mmu_lsu_writeback_w ;
  wire \u0.mmu_mxr_w ;
  wire [31:0] \u0.mmu_satp_w ;
  wire \u0.mmu_store_fault_w ;
  wire \u0.mmu_sum_w ;
  wire \u0.mul_hold_w ;
  wire \u0.mul_opcode_invalid_w ;
  wire [31:0] \u0.mul_opcode_opcode_w ;
  wire [31:0] \u0.mul_opcode_pc_w ;
  wire [4:0] \u0.mul_opcode_ra_idx_w ;
  wire [31:0] \u0.mul_opcode_ra_operand_w ;
  wire [4:0] \u0.mul_opcode_rb_idx_w ;
  wire [31:0] \u0.mul_opcode_rb_operand_w ;
  wire [4:0] \u0.mul_opcode_rd_idx_w ;
  wire \u0.mul_opcode_valid_w ;
  wire \u0.opcode_invalid_w ;
  wire [31:0] \u0.opcode_opcode_w ;
  wire [31:0] \u0.opcode_pc_w ;
  wire [4:0] \u0.opcode_ra_idx_w ;
  wire [31:0] \u0.opcode_ra_operand_w ;
  wire [4:0] \u0.opcode_rb_idx_w ;
  wire [31:0] \u0.opcode_rb_operand_w ;
  wire [4:0] \u0.opcode_rd_idx_w ;
  wire [31:0] \u0.reset_vector_i ;
  wire \u0.rst_i ;
  wire \u0.squash_decode_w ;
  wire \u0.take_interrupt_w ;
  wire [31:0] \u0.u_csr.branch_csr_pc_o ;
  wire \u0.u_csr.branch_csr_request_o ;
  reg \u0.u_csr.branch_q ;
  reg [31:0] \u0.u_csr.branch_target_q ;
  wire \u0.u_csr.clk_i ;
  wire \u0.u_csr.clr_r ;
  wire [31:0] \u0.u_csr.cpu_id_i ;
  wire \u0.u_csr.csr_branch_w ;
  wire \u0.u_csr.csr_fault_r ;
  wire [1:0] \u0.u_csr.csr_priv_r ;
  wire [31:0] \u0.u_csr.csr_rdata_w ;
  wire [5:0] \u0.u_csr.csr_result_e1_exception_o ;
  wire [31:0] \u0.u_csr.csr_result_e1_value_o ;
  wire [31:0] \u0.u_csr.csr_result_e1_wdata_o ;
  wire \u0.u_csr.csr_result_e1_write_o ;
  wire [31:0] \u0.u_csr.csr_target_w ;
  reg [31:0] \u0.u_csr.csr_wdata_e1_q ;
  wire \u0.u_csr.csr_write_r ;
  wire [31:0] \u0.u_csr.csr_writeback_exception_addr_i ;
  wire [5:0] \u0.u_csr.csr_writeback_exception_i ;
  wire [31:0] \u0.u_csr.csr_writeback_exception_pc_i ;
  wire [11:0] \u0.u_csr.csr_writeback_waddr_i ;
  wire [31:0] \u0.u_csr.csr_writeback_wdata_i ;
  wire \u0.u_csr.csr_writeback_write_i ;
  wire \u0.u_csr.csrrc_w ;
  wire \u0.u_csr.csrrci_w ;
  wire \u0.u_csr.csrrs_w ;
  wire \u0.u_csr.csrrsi_w ;
  wire \u0.u_csr.csrrw_w ;
  wire \u0.u_csr.csrrwi_w ;
  wire [1:0] \u0.u_csr.current_priv_w ;
  wire [31:0] \u0.u_csr.data_r ;
  reg [5:0] \u0.u_csr.exception_e1_q ;
  wire \u0.u_csr.ifence_o ;
  wire \u0.u_csr.ifence_q ;
  wire \u0.u_csr.ifence_w ;
  wire \u0.u_csr.interrupt_inhibit_i ;
  wire [31:0] \u0.u_csr.interrupt_w ;
  wire \u0.u_csr.intr_i ;
  wire [31:0] \u0.u_csr.misa_w ;
  wire \u0.u_csr.mmu_mxr_o ;
  wire [31:0] \u0.u_csr.mmu_satp_o ;
  wire \u0.u_csr.mmu_sum_o ;
  wire \u0.u_csr.opcode_invalid_i ;
  wire [31:0] \u0.u_csr.opcode_opcode_i ;
  wire [31:0] \u0.u_csr.opcode_pc_i ;
  wire [4:0] \u0.u_csr.opcode_ra_idx_i ;
  wire [31:0] \u0.u_csr.opcode_ra_operand_i ;
  wire [4:0] \u0.u_csr.opcode_rb_idx_i ;
  wire [31:0] \u0.u_csr.opcode_rb_operand_i ;
  wire [4:0] \u0.u_csr.opcode_rd_idx_i ;
  wire \u0.u_csr.opcode_valid_i ;
  reg [31:0] \u0.u_csr.rd_result_e1_q ;
  reg \u0.u_csr.rd_valid_e1_q ;
  reg \u0.u_csr.reset_q ;
  wire [31:0] \u0.u_csr.reset_vector_i ;
  wire \u0.u_csr.rst_i ;
  wire [31:0] \u0.u_csr.satp_reg_w ;
  wire \u0.u_csr.satp_update_w ;
  wire \u0.u_csr.set_r ;
  wire \u0.u_csr.sfence_w ;
  wire [31:0] \u0.u_csr.status_reg_w ;
  wire \u0.u_csr.take_interrupt_o ;
  reg \u0.u_csr.take_interrupt_q ;
  wire \u0.u_csr.timer_irq_w ;
  wire \u0.u_csr.u_csrfile.branch_r ;
  wire [31:0] \u0.u_csr.u_csrfile.branch_target_r ;
  wire \u0.u_csr.u_csrfile.buffer_mip_w ;
  wire \u0.u_csr.u_csrfile.clk_i ;
  wire [31:0] \u0.u_csr.u_csrfile.cpu_id_i ;
  wire \u0.u_csr.u_csrfile.csr_branch_o ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mcause_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mcause_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mcycle_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mcycle_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mepc_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mepc_r ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mideleg_q ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mie_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mie_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mip_next_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mip_next_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mip_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mip_r ;
  reg \u0.u_csr.u_csrfile.csr_mip_upd_q ;
  wire [1:0] \u0.u_csr.u_csrfile.csr_mpriv_q ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mscratch_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mscratch_r ;
  reg \u0.u_csr.u_csrfile.csr_mtime_ie_q ;
  wire \u0.u_csr.u_csrfile.csr_mtime_ie_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mtimecmp_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mtimecmp_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mtval_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mtval_r ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_mtvec_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_mtvec_r ;
  wire [11:0] \u0.u_csr.u_csrfile.csr_raddr_i ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_rdata_o ;
  wire \u0.u_csr.u_csrfile.csr_ren_i ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_satp_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_sepc_q ;
  reg [31:0] \u0.u_csr.u_csrfile.csr_sr_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_sr_r ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_stvec_q ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_target_o ;
  wire [11:0] \u0.u_csr.u_csrfile.csr_waddr_i ;
  wire [31:0] \u0.u_csr.u_csrfile.csr_wdata_i ;
  wire [31:0] \u0.u_csr.u_csrfile.exception_addr_i ;
  wire [5:0] \u0.u_csr.u_csrfile.exception_i ;
  wire [31:0] \u0.u_csr.u_csrfile.exception_pc_i ;
  wire \u0.u_csr.u_csrfile.exception_s_w ;
  wire \u0.u_csr.u_csrfile.ext_intr_i ;
  wire [31:0] \u0.u_csr.u_csrfile.interrupt_o ;
  wire [31:0] \u0.u_csr.u_csrfile.irq_masked_r ;
  wire [31:0] \u0.u_csr.u_csrfile.irq_pending_r ;
  reg [1:0] \u0.u_csr.u_csrfile.irq_priv_q ;
  wire [1:0] \u0.u_csr.u_csrfile.irq_priv_r ;
  wire \u0.u_csr.u_csrfile.is_exception_w ;
  wire [31:0] \u0.u_csr.u_csrfile.misa_i ;
  wire [1:0] \u0.u_csr.u_csrfile.priv_o ;
  wire [31:0] \u0.u_csr.u_csrfile.rdata_r ;
  wire \u0.u_csr.u_csrfile.rst_i ;
  wire [31:0] \u0.u_csr.u_csrfile.satp_o ;
  wire [31:0] \u0.u_csr.u_csrfile.status_o ;
  wire \u0.u_csr.u_csrfile.timer_intr_i ;
  wire \u0.u_decode.clk_i ;
  wire \u0.u_decode.enable_muldiv_w ;
  wire \u0.u_decode.fetch_in_accept_o ;
  wire \u0.u_decode.fetch_in_fault_fetch_i ;
  wire \u0.u_decode.fetch_in_fault_page_i ;
  wire [31:0] \u0.u_decode.fetch_in_instr_i ;
  wire [31:0] \u0.u_decode.fetch_in_pc_i ;
  wire \u0.u_decode.fetch_in_valid_i ;
  wire \u0.u_decode.fetch_out_accept_i ;
  wire \u0.u_decode.fetch_out_fault_fetch_o ;
  wire \u0.u_decode.fetch_out_fault_page_o ;
  wire \u0.u_decode.fetch_out_instr_branch_o ;
  wire \u0.u_decode.fetch_out_instr_csr_o ;
  wire \u0.u_decode.fetch_out_instr_div_o ;
  wire \u0.u_decode.fetch_out_instr_exec_o ;
  wire \u0.u_decode.fetch_out_instr_invalid_o ;
  wire \u0.u_decode.fetch_out_instr_lsu_o ;
  wire \u0.u_decode.fetch_out_instr_mul_o ;
  wire [31:0] \u0.u_decode.fetch_out_instr_o ;
  wire \u0.u_decode.fetch_out_instr_rd_valid_o ;
  wire [31:0] \u0.u_decode.fetch_out_pc_o ;
  wire \u0.u_decode.fetch_out_valid_o ;
  wire [31:0] \u0.u_decode.genblk1.fetch_in_instr_w ;
  wire \u0.u_decode.genblk1.u_dec.branch_o ;
  wire \u0.u_decode.genblk1.u_dec.csr_o ;
  wire \u0.u_decode.genblk1.u_dec.div_o ;
  wire \u0.u_decode.genblk1.u_dec.enable_muldiv_i ;
  wire \u0.u_decode.genblk1.u_dec.exec_o ;
  wire \u0.u_decode.genblk1.u_dec.fetch_fault_i ;
  wire \u0.u_decode.genblk1.u_dec.invalid_o ;
  wire \u0.u_decode.genblk1.u_dec.invalid_w ;
  wire \u0.u_decode.genblk1.u_dec.lsu_o ;
  wire \u0.u_decode.genblk1.u_dec.mul_o ;
  wire [31:0] \u0.u_decode.genblk1.u_dec.opcode_i ;
  wire \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  wire \u0.u_decode.genblk1.u_dec.valid_i ;
  wire \u0.u_decode.rst_i ;
  wire \u0.u_decode.squash_decode_i ;
  wire \u0.u_div.clk_i ;
  reg \u0.u_div.div_busy_q ;
  wire \u0.u_div.div_complete_w ;
  reg \u0.u_div.div_inst_q ;
  wire \u0.u_div.div_operation_w ;
  wire \u0.u_div.div_rem_inst_w ;
  wire [31:0] \u0.u_div.div_result_r ;
  wire \u0.u_div.div_start_w ;
  reg [31:0] \u0.u_div.dividend_q ;
  reg [62:0] \u0.u_div.divisor_q ;
  reg \u0.u_div.invert_res_q ;
  wire \u0.u_div.opcode_invalid_i ;
  wire [31:0] \u0.u_div.opcode_opcode_i ;
  wire [31:0] \u0.u_div.opcode_pc_i ;
  wire [4:0] \u0.u_div.opcode_ra_idx_i ;
  wire [31:0] \u0.u_div.opcode_ra_operand_i ;
  wire [4:0] \u0.u_div.opcode_rb_idx_i ;
  wire [31:0] \u0.u_div.opcode_rb_operand_i ;
  wire [4:0] \u0.u_div.opcode_rd_idx_i ;
  wire \u0.u_div.opcode_valid_i ;
  reg [31:0] \u0.u_div.q_mask_q ;
  reg [31:0] \u0.u_div.quotient_q ;
  wire \u0.u_div.rst_i ;
  wire \u0.u_div.signed_operation_w ;
  reg \u0.u_div.valid_q ;
  reg [31:0] \u0.u_div.wb_result_q ;
  wire \u0.u_div.writeback_valid_o ;
  wire [31:0] \u0.u_div.writeback_value_o ;
  wire [3:0] \u0.u_exec.alu_func_r ;
  wire [31:0] \u0.u_exec.alu_input_a_r ;
  wire [31:0] \u0.u_exec.alu_input_b_r ;
  wire [31:0] \u0.u_exec.alu_p_w ;
  wire [31:0] \u0.u_exec.bimm_r ;
  wire [31:0] \u0.u_exec.branch_d_pc_o ;
  wire [1:0] \u0.u_exec.branch_d_priv_o ;
  wire \u0.u_exec.branch_d_request_o ;
  wire \u0.u_exec.branch_r ;
  wire \u0.u_exec.branch_taken_r ;
  wire [31:0] \u0.u_exec.branch_target_r ;
  wire \u0.u_exec.clk_i ;
  wire [31:0] \u0.u_exec.greater_than_signed$func$../../core/riscv/riscv_exec.v:362$760.v ;
  wire [31:0] \u0.u_exec.greater_than_signed$func$../../core/riscv/riscv_exec.v:362$760.x ;
  wire [31:0] \u0.u_exec.greater_than_signed$func$../../core/riscv/riscv_exec.v:362$760.y ;
  wire \u0.u_exec.hold_i ;
  wire [31:0] \u0.u_exec.imm12_r ;
  wire [31:0] \u0.u_exec.imm20_r ;
  wire [31:0] \u0.u_exec.jimm20_r ;
  wire [31:0] \u0.u_exec.less_than_signed$func$../../core/riscv/riscv_exec.v:357$759.v ;
  wire [31:0] \u0.u_exec.less_than_signed$func$../../core/riscv/riscv_exec.v:357$759.x ;
  wire [31:0] \u0.u_exec.less_than_signed$func$../../core/riscv/riscv_exec.v:357$759.y ;
  wire \u0.u_exec.opcode_invalid_i ;
  wire [31:0] \u0.u_exec.opcode_opcode_i ;
  wire [31:0] \u0.u_exec.opcode_pc_i ;
  wire [4:0] \u0.u_exec.opcode_ra_idx_i ;
  wire [31:0] \u0.u_exec.opcode_ra_operand_i ;
  wire [4:0] \u0.u_exec.opcode_rb_idx_i ;
  wire [31:0] \u0.u_exec.opcode_rb_operand_i ;
  wire [4:0] \u0.u_exec.opcode_rd_idx_i ;
  wire \u0.u_exec.opcode_valid_i ;
  reg [31:0] \u0.u_exec.result_q ;
  wire \u0.u_exec.rst_i ;
  wire [4:0] \u0.u_exec.shamt_r ;
  wire [31:0] \u0.u_exec.u_alu.alu_a_i ;
  wire [31:0] \u0.u_exec.u_alu.alu_b_i ;
  wire [3:0] \u0.u_exec.u_alu.alu_op_i ;
  wire [31:0] \u0.u_exec.u_alu.alu_p_o ;
  wire [31:0] \u0.u_exec.u_alu.result_r ;
  wire [31:0] \u0.u_exec.u_alu.sub_res_w ;
  wire [31:0] \u0.u_exec.writeback_value_o ;
  reg \u0.u_fetch.active_q ;
  reg \u0.u_fetch.branch_d_q ;
  wire [31:0] \u0.u_fetch.branch_pc_i ;
  reg [31:0] \u0.u_fetch.branch_pc_q ;
  wire [31:0] \u0.u_fetch.branch_pc_w ;
  reg \u0.u_fetch.branch_q ;
  wire \u0.u_fetch.branch_request_i ;
  wire \u0.u_fetch.branch_w ;
  wire \u0.u_fetch.clk_i ;
  wire \u0.u_fetch.fetch_accept_i ;
  wire \u0.u_fetch.fetch_fault_fetch_o ;
  wire \u0.u_fetch.fetch_fault_page_o ;
  wire [31:0] \u0.u_fetch.fetch_instr_o ;
  wire \u0.u_fetch.fetch_invalidate_i ;
  wire [31:0] \u0.u_fetch.fetch_pc_o ;
  wire \u0.u_fetch.fetch_resp_drop_w ;
  wire \u0.u_fetch.fetch_valid_o ;
  wire \u0.u_fetch.icache_accept_i ;
  wire \u0.u_fetch.icache_busy_w ;
  wire \u0.u_fetch.icache_error_i ;
  reg \u0.u_fetch.icache_fetch_q ;
  wire \u0.u_fetch.icache_flush_o ;
  wire [31:0] \u0.u_fetch.icache_inst_i ;
  wire \u0.u_fetch.icache_invalidate_o ;
  wire \u0.u_fetch.icache_invalidate_q ;
  wire \u0.u_fetch.icache_page_fault_i ;
  wire [31:0] \u0.u_fetch.icache_pc_o ;
  wire [31:0] \u0.u_fetch.icache_pc_w ;
  wire \u0.u_fetch.icache_rd_o ;
  wire \u0.u_fetch.icache_valid_i ;
  reg [31:0] \u0.u_fetch.pc_d_q ;
  reg [31:0] \u0.u_fetch.pc_f_q ;
  wire \u0.u_fetch.rst_i ;
  reg [65:0] \u0.u_fetch.skid_buffer_q ;
  reg \u0.u_fetch.skid_valid_q ;
  wire \u0.u_fetch.squash_decode_o ;
  wire \u0.u_fetch.stall_w ;
  wire [31:0] \u0.u_issue.branch_csr_pc_i ;
  wire \u0.u_issue.branch_csr_request_i ;
  wire [31:0] \u0.u_issue.branch_d_exec_pc_i ;
  wire [1:0] \u0.u_issue.branch_d_exec_priv_i ;
  wire \u0.u_issue.branch_d_exec_request_i ;
  wire [31:0] \u0.u_issue.branch_pc_o ;
  wire \u0.u_issue.branch_request_o ;
  wire \u0.u_issue.clk_i ;
  wire \u0.u_issue.csr_opcode_invalid_o ;
  wire [31:0] \u0.u_issue.csr_opcode_opcode_o ;
  wire [31:0] \u0.u_issue.csr_opcode_pc_o ;
  wire [4:0] \u0.u_issue.csr_opcode_ra_idx_o ;
  wire [31:0] \u0.u_issue.csr_opcode_ra_operand_o ;
  wire [4:0] \u0.u_issue.csr_opcode_rb_idx_o ;
  wire [31:0] \u0.u_issue.csr_opcode_rb_operand_o ;
  wire [4:0] \u0.u_issue.csr_opcode_rd_idx_o ;
  wire \u0.u_issue.csr_opcode_valid_o ;
  reg \u0.u_issue.csr_pending_q ;
  wire [5:0] \u0.u_issue.csr_result_e1_exception_i ;
  wire [31:0] \u0.u_issue.csr_result_e1_value_i ;
  wire [31:0] \u0.u_issue.csr_result_e1_wdata_i ;
  wire \u0.u_issue.csr_result_e1_write_i ;
  wire [31:0] \u0.u_issue.csr_writeback_exception_addr_o ;
  wire [5:0] \u0.u_issue.csr_writeback_exception_o ;
  wire [31:0] \u0.u_issue.csr_writeback_exception_pc_o ;
  wire [11:0] \u0.u_issue.csr_writeback_waddr_o ;
  wire [31:0] \u0.u_issue.csr_writeback_wdata_o ;
  wire \u0.u_issue.csr_writeback_write_o ;
  wire \u0.u_issue.div_opcode_valid_o ;
  reg \u0.u_issue.div_pending_q ;
  wire \u0.u_issue.enable_mul_bypass_w ;
  wire \u0.u_issue.enable_muldiv_w ;
  wire \u0.u_issue.exec_hold_o ;
  wire \u0.u_issue.exec_opcode_valid_o ;
  wire \u0.u_issue.fetch_accept_o ;
  wire \u0.u_issue.fetch_fault_fetch_i ;
  wire \u0.u_issue.fetch_fault_page_i ;
  wire \u0.u_issue.fetch_instr_branch_i ;
  wire \u0.u_issue.fetch_instr_csr_i ;
  wire \u0.u_issue.fetch_instr_div_i ;
  wire \u0.u_issue.fetch_instr_exec_i ;
  wire [31:0] \u0.u_issue.fetch_instr_i ;
  wire \u0.u_issue.fetch_instr_invalid_i ;
  wire \u0.u_issue.fetch_instr_lsu_i ;
  wire \u0.u_issue.fetch_instr_mul_i ;
  wire \u0.u_issue.fetch_instr_rd_valid_i ;
  wire [31:0] \u0.u_issue.fetch_pc_i ;
  wire \u0.u_issue.fetch_valid_i ;
  wire \u0.u_issue.interrupt_inhibit_o ;
  wire \u0.u_issue.issue_branch_w ;
  wire \u0.u_issue.issue_csr_w ;
  wire \u0.u_issue.issue_div_w ;
  wire \u0.u_issue.issue_exec_w ;
  wire [4:0] \u0.u_issue.issue_fault_w ;
  wire \u0.u_issue.issue_invalid_w ;
  wire \u0.u_issue.issue_lsu_w ;
  wire \u0.u_issue.issue_mul_w ;
  wire [4:0] \u0.u_issue.issue_ra_idx_w ;
  wire [31:0] \u0.u_issue.issue_ra_value_r ;
  wire [31:0] \u0.u_issue.issue_ra_value_w ;
  wire [4:0] \u0.u_issue.issue_rb_idx_w ;
  wire [31:0] \u0.u_issue.issue_rb_value_r ;
  wire [31:0] \u0.u_issue.issue_rb_value_w ;
  wire [4:0] \u0.u_issue.issue_rd_idx_w ;
  wire \u0.u_issue.issue_sb_alloc_w ;
  wire \u0.u_issue.lsu_opcode_invalid_o ;
  wire [31:0] \u0.u_issue.lsu_opcode_opcode_o ;
  wire [31:0] \u0.u_issue.lsu_opcode_pc_o ;
  wire [4:0] \u0.u_issue.lsu_opcode_ra_idx_o ;
  wire [31:0] \u0.u_issue.lsu_opcode_ra_operand_o ;
  wire [4:0] \u0.u_issue.lsu_opcode_rb_idx_o ;
  wire [31:0] \u0.u_issue.lsu_opcode_rb_operand_o ;
  wire [4:0] \u0.u_issue.lsu_opcode_rd_idx_o ;
  wire \u0.u_issue.lsu_opcode_valid_o ;
  wire \u0.u_issue.lsu_stall_i ;
  wire \u0.u_issue.mul_hold_o ;
  wire \u0.u_issue.mul_opcode_invalid_o ;
  wire [31:0] \u0.u_issue.mul_opcode_opcode_o ;
  wire [31:0] \u0.u_issue.mul_opcode_pc_o ;
  wire [4:0] \u0.u_issue.mul_opcode_ra_idx_o ;
  wire [31:0] \u0.u_issue.mul_opcode_ra_operand_o ;
  wire [4:0] \u0.u_issue.mul_opcode_rb_idx_o ;
  wire [31:0] \u0.u_issue.mul_opcode_rb_operand_o ;
  wire [4:0] \u0.u_issue.mul_opcode_rd_idx_o ;
  wire \u0.u_issue.mul_opcode_valid_o ;
  wire \u0.u_issue.opcode_accept_r ;
  wire \u0.u_issue.opcode_invalid_o ;
  wire \u0.u_issue.opcode_issue_r ;
  wire [31:0] \u0.u_issue.opcode_opcode_o ;
  wire [31:0] \u0.u_issue.opcode_pc_o ;
  wire [4:0] \u0.u_issue.opcode_ra_idx_o ;
  wire [31:0] \u0.u_issue.opcode_ra_operand_o ;
  wire [4:0] \u0.u_issue.opcode_rb_idx_o ;
  wire [31:0] \u0.u_issue.opcode_rb_operand_o ;
  wire [4:0] \u0.u_issue.opcode_rd_idx_o ;
  wire \u0.u_issue.opcode_valid_w ;
  wire \u0.u_issue.pipe_branch_e1_w ;
  wire \u0.u_issue.pipe_csr_wb_w ;
  wire [5:0] \u0.u_issue.pipe_exception_wb_w ;
  wire \u0.u_issue.pipe_load_e1_w ;
  wire \u0.u_issue.pipe_load_e2_w ;
  wire \u0.u_issue.pipe_mul_e1_w ;
  wire \u0.u_issue.pipe_mul_e2_w ;
  wire [31:0] \u0.u_issue.pipe_opc_wb_w ;
  wire [31:0] \u0.u_issue.pipe_opcode_e1_w ;
  wire [31:0] \u0.u_issue.pipe_pc_e1_w ;
  wire [31:0] \u0.u_issue.pipe_pc_wb_w ;
  wire [4:0] \u0.u_issue.pipe_rd_e1_w ;
  wire [4:0] \u0.u_issue.pipe_rd_e2_w ;
  wire [4:0] \u0.u_issue.pipe_rd_wb_w ;
  wire [31:0] \u0.u_issue.pipe_result_e2_w ;
  wire [31:0] \u0.u_issue.pipe_result_wb_w ;
  wire \u0.u_issue.pipe_squash_e1_e2_w ;
  wire \u0.u_issue.pipe_stall_raw_w ;
  wire \u0.u_issue.pipe_store_e1_w ;
  wire \u0.u_issue.pipe_valid_wb_w ;
  wire \u0.u_issue.rst_i ;
  wire \u0.u_issue.squash_w ;
  wire \u0.u_issue.stall_w ;
  wire \u0.u_issue.take_interrupt_i ;
  wire \u0.u_issue.u_pipe_ctrl.alu_e1_w ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.alu_result_e1_i ;
  wire \u0.u_issue.u_pipe_ctrl.branch_e1_o ;
  wire \u0.u_issue.u_pipe_ctrl.branch_misaligned_w ;
  wire \u0.u_issue.u_pipe_ctrl.clk_i ;
  wire \u0.u_issue.u_pipe_ctrl.csr_e1_w ;
  wire [5:0] \u0.u_issue.u_pipe_ctrl.csr_result_exception_e1_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.csr_result_value_e1_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.csr_result_wdata_e1_i ;
  wire \u0.u_issue.u_pipe_ctrl.csr_result_write_e1_i ;
  wire [11:0] \u0.u_issue.u_pipe_ctrl.csr_waddr_wb_o ;
  wire \u0.u_issue.u_pipe_ctrl.csr_wb_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.csr_wdata_e2_q ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q ;
  reg \u0.u_issue.u_pipe_ctrl.csr_wr_e2_q ;
  reg \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q ;
  wire \u0.u_issue.u_pipe_ctrl.csr_write_wb_o ;
  reg [9:0] \u0.u_issue.u_pipe_ctrl.ctrl_e1_q ;
  reg [9:0] \u0.u_issue.u_pipe_ctrl.ctrl_e2_q ;
  reg [9:0] \u0.u_issue.u_pipe_ctrl.ctrl_wb_q ;
  wire \u0.u_issue.u_pipe_ctrl.div_complete_i ;
  wire \u0.u_issue.u_pipe_ctrl.div_e1_w ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.div_result_i ;
  reg [5:0] \u0.u_issue.u_pipe_ctrl.exception_e1_q ;
  reg [5:0] \u0.u_issue.u_pipe_ctrl.exception_e2_q ;
  wire [5:0] \u0.u_issue.u_pipe_ctrl.exception_e2_r ;
  wire [5:0] \u0.u_issue.u_pipe_ctrl.exception_wb_o ;
  reg [5:0] \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  wire \u0.u_issue.u_pipe_ctrl.issue_accept_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_branch_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_branch_taken_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.issue_branch_target_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_csr_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_div_i ;
  wire [5:0] \u0.u_issue.u_pipe_ctrl.issue_exception_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_lsu_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_mul_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.issue_opcode_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.issue_operand_ra_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.issue_operand_rb_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.issue_pc_i ;
  wire [4:0] \u0.u_issue.u_pipe_ctrl.issue_rd_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_rd_valid_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_stall_i ;
  wire \u0.u_issue.u_pipe_ctrl.issue_valid_i ;
  wire \u0.u_issue.u_pipe_ctrl.load_e1_o ;
  wire \u0.u_issue.u_pipe_ctrl.load_e2_o ;
  wire \u0.u_issue.u_pipe_ctrl.mem_complete_i ;
  wire [5:0] \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.mem_result_e2_i ;
  wire \u0.u_issue.u_pipe_ctrl.mul_e1_o ;
  wire \u0.u_issue.u_pipe_ctrl.mul_e2_o ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.mul_result_e2_i ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.opcode_e1_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.opcode_e1_q ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.opcode_e2_q ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.opcode_wb_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.opcode_wb_q ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.pc_e1_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.pc_e1_q ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.pc_e2_q ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.pc_wb_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  wire [4:0] \u0.u_issue.u_pipe_ctrl.rd_e1_o ;
  wire [4:0] \u0.u_issue.u_pipe_ctrl.rd_e2_o ;
  wire [4:0] \u0.u_issue.u_pipe_ctrl.rd_wb_o ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.result_e2_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.result_e2_q ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.result_e2_r ;
  wire [31:0] \u0.u_issue.u_pipe_ctrl.result_wb_o ;
  reg [31:0] \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  wire \u0.u_issue.u_pipe_ctrl.rst_i ;
  wire \u0.u_issue.u_pipe_ctrl.squash_e1_e2_i ;
  wire \u0.u_issue.u_pipe_ctrl.squash_e1_e2_o ;
  reg \u0.u_issue.u_pipe_ctrl.squash_e1_e2_q ;
  wire \u0.u_issue.u_pipe_ctrl.squash_e1_e2_w ;
  wire \u0.u_issue.u_pipe_ctrl.squash_wb_i ;
  wire \u0.u_issue.u_pipe_ctrl.stall_o ;
  wire \u0.u_issue.u_pipe_ctrl.store_e1_o ;
  wire \u0.u_issue.u_pipe_ctrl.take_interrupt_i ;
  reg \u0.u_issue.u_pipe_ctrl.valid_e1_q ;
  reg \u0.u_issue.u_pipe_ctrl.valid_e2_q ;
  wire \u0.u_issue.u_pipe_ctrl.valid_e2_w ;
  wire \u0.u_issue.u_pipe_ctrl.valid_wb_o ;
  reg \u0.u_issue.u_pipe_ctrl.valid_wb_q ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.ra0_value_r ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.rb0_value_r ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r10_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r11_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r12_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r13_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r14_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r15_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r16_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r17_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r18_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r19_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r1_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r20_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r21_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r22_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r23_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r24_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r25_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r26_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r27_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r28_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r29_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r2_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r30_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r31_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r3_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r4_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r5_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r6_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r7_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r8_q ;
  reg [31:0] \u0.u_issue.u_regfile.REGFILE.reg_r9_q ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x0_zero_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x10_a0_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x11_a1_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x12_a2_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x13_a3_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x14_a4_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x15_a5_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x16_a6_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x17_a7_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x18_s2_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x19_s3_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x1_ra_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x20_s4_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x21_s5_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x22_s6_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x23_s7_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x24_s8_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x25_s9_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x26_s10_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x27_s11_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x28_t3_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x29_t4_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x2_sp_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x30_t5_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x31_t6_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x3_gp_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x4_tp_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x5_t0_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x6_t1_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x7_t2_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x8_s0_w ;
  wire [31:0] \u0.u_issue.u_regfile.REGFILE.x9_s1_w ;
  wire \u0.u_issue.u_regfile.clk_i ;
  wire [4:0] \u0.u_issue.u_regfile.ra0_i ;
  wire [31:0] \u0.u_issue.u_regfile.ra0_value_o ;
  wire [4:0] \u0.u_issue.u_regfile.rb0_i ;
  wire [31:0] \u0.u_issue.u_regfile.rb0_value_o ;
  wire [4:0] \u0.u_issue.u_regfile.rd0_i ;
  wire [31:0] \u0.u_issue.u_regfile.rd0_value_i ;
  wire \u0.u_issue.u_regfile.rst_i ;
  wire \u0.u_issue.writeback_div_valid_i ;
  wire [31:0] \u0.u_issue.writeback_div_value_i ;
  wire [31:0] \u0.u_issue.writeback_exec_value_i ;
  wire [5:0] \u0.u_issue.writeback_mem_exception_i ;
  wire \u0.u_issue.writeback_mem_valid_i ;
  wire [31:0] \u0.u_issue.writeback_mem_value_i ;
  wire [31:0] \u0.u_issue.writeback_mul_value_i ;
  wire [1:0] \u0.u_lsu.addr_lsb_r ;
  wire \u0.u_lsu.clk_i ;
  wire \u0.u_lsu.complete_err_e2_w ;
  wire \u0.u_lsu.complete_ok_e2_w ;
  wire \u0.u_lsu.dcache_flush_w ;
  wire \u0.u_lsu.dcache_invalidate_w ;
  wire \u0.u_lsu.dcache_writeback_w ;
  wire \u0.u_lsu.delay_lsu_e2_w ;
  wire \u0.u_lsu.fault_load_align_w ;
  wire \u0.u_lsu.fault_load_bus_w ;
  wire \u0.u_lsu.fault_load_page_w ;
  wire \u0.u_lsu.fault_store_align_w ;
  wire \u0.u_lsu.fault_store_bus_w ;
  wire \u0.u_lsu.fault_store_page_w ;
  wire \u0.u_lsu.issue_lsu_e1_w ;
  wire \u0.u_lsu.load_byte_r ;
  wire \u0.u_lsu.load_half_r ;
  wire \u0.u_lsu.load_inst_w ;
  wire \u0.u_lsu.load_signed_inst_w ;
  wire \u0.u_lsu.load_signed_r ;
  wire \u0.u_lsu.mem_accept_i ;
  wire \u0.u_lsu.mem_ack_i ;
  wire [31:0] \u0.u_lsu.mem_addr_o ;
  reg [31:0] \u0.u_lsu.mem_addr_q ;
  wire [31:0] \u0.u_lsu.mem_addr_r ;
  wire \u0.u_lsu.mem_cacheable_o ;
  wire \u0.u_lsu.mem_cacheable_q ;
  wire [31:0] \u0.u_lsu.mem_data_r ;
  wire [31:0] \u0.u_lsu.mem_data_rd_i ;
  wire [31:0] \u0.u_lsu.mem_data_wr_o ;
  reg [31:0] \u0.u_lsu.mem_data_wr_q ;
  wire \u0.u_lsu.mem_error_i ;
  wire \u0.u_lsu.mem_flush_o ;
  reg \u0.u_lsu.mem_flush_q ;
  wire \u0.u_lsu.mem_invalidate_o ;
  reg \u0.u_lsu.mem_invalidate_q ;
  wire \u0.u_lsu.mem_load_fault_i ;
  reg \u0.u_lsu.mem_load_q ;
  reg \u0.u_lsu.mem_ls_q ;
  wire \u0.u_lsu.mem_rd_o ;
  reg \u0.u_lsu.mem_rd_q ;
  wire \u0.u_lsu.mem_rd_r ;
  wire [10:0] \u0.u_lsu.mem_req_tag_o ;
  wire [10:0] \u0.u_lsu.mem_resp_tag_i ;
  wire \u0.u_lsu.mem_store_fault_i ;
  reg \u0.u_lsu.mem_unaligned_e1_q ;
  reg \u0.u_lsu.mem_unaligned_e2_q ;
  wire \u0.u_lsu.mem_unaligned_r ;
  wire [3:0] \u0.u_lsu.mem_wr_o ;
  reg [3:0] \u0.u_lsu.mem_wr_q ;
  wire [3:0] \u0.u_lsu.mem_wr_r ;
  wire \u0.u_lsu.mem_writeback_o ;
  reg \u0.u_lsu.mem_writeback_q ;
  reg \u0.u_lsu.mem_xb_q ;
  reg \u0.u_lsu.mem_xh_q ;
  wire \u0.u_lsu.opcode_invalid_i ;
  wire [31:0] \u0.u_lsu.opcode_opcode_i ;
  wire [31:0] \u0.u_lsu.opcode_pc_i ;
  wire [4:0] \u0.u_lsu.opcode_ra_idx_i ;
  wire [31:0] \u0.u_lsu.opcode_ra_operand_i ;
  wire [4:0] \u0.u_lsu.opcode_rb_idx_i ;
  wire [31:0] \u0.u_lsu.opcode_rb_operand_i ;
  wire [4:0] \u0.u_lsu.opcode_rd_idx_i ;
  wire \u0.u_lsu.opcode_valid_i ;
  reg \u0.u_lsu.pending_lsu_e2_q ;
  wire \u0.u_lsu.req_lb_w ;
  wire \u0.u_lsu.req_lh_w ;
  wire \u0.u_lsu.req_sb_w ;
  wire \u0.u_lsu.req_sh_lh_w ;
  wire \u0.u_lsu.req_sh_w ;
  wire \u0.u_lsu.req_sw_lw_w ;
  wire [31:0] \u0.u_lsu.resp_addr_w ;
  wire \u0.u_lsu.resp_byte_w ;
  wire \u0.u_lsu.resp_half_w ;
  wire \u0.u_lsu.resp_load_w ;
  wire \u0.u_lsu.resp_signed_w ;
  wire \u0.u_lsu.rst_i ;
  wire \u0.u_lsu.stall_o ;
  wire \u0.u_lsu.u_lsu_request.accept_o ;
  wire \u0.u_lsu.u_lsu_request.clk_i ;
  reg [1:0] \u0.u_lsu.u_lsu_request.count_q ;
  wire [35:0] \u0.u_lsu.u_lsu_request.data_in_i ;
  wire [35:0] \u0.u_lsu.u_lsu_request.data_out_o ;
  wire \u0.u_lsu.u_lsu_request.pop_i ;
  wire \u0.u_lsu.u_lsu_request.push_i ;
  reg [35:0] \u0.u_lsu.u_lsu_request.ram_q[0] ;
  reg [35:0] \u0.u_lsu.u_lsu_request.ram_q[1] ;
  reg \u0.u_lsu.u_lsu_request.rd_ptr_q ;
  wire \u0.u_lsu.u_lsu_request.rst_i ;
  wire \u0.u_lsu.u_lsu_request.valid_o ;
  reg \u0.u_lsu.u_lsu_request.wr_ptr_q ;
  wire [31:0] \u0.u_lsu.wb_result_r ;
  wire [5:0] \u0.u_lsu.writeback_exception_o ;
  wire \u0.u_lsu.writeback_valid_o ;
  wire [31:0] \u0.u_lsu.writeback_value_o ;
  wire \u0.u_mmu.clk_i ;
  wire \u0.u_mmu.fetch_in_accept_o ;
  wire \u0.u_mmu.fetch_in_error_o ;
  wire \u0.u_mmu.fetch_in_fault_o ;
  wire \u0.u_mmu.fetch_in_flush_i ;
  wire [31:0] \u0.u_mmu.fetch_in_inst_o ;
  wire \u0.u_mmu.fetch_in_invalidate_i ;
  wire [31:0] \u0.u_mmu.fetch_in_pc_i ;
  wire \u0.u_mmu.fetch_in_rd_i ;
  wire \u0.u_mmu.fetch_in_valid_o ;
  wire \u0.u_mmu.fetch_out_accept_i ;
  wire \u0.u_mmu.fetch_out_error_i ;
  wire \u0.u_mmu.fetch_out_flush_o ;
  wire [31:0] \u0.u_mmu.fetch_out_inst_i ;
  wire \u0.u_mmu.fetch_out_invalidate_o ;
  wire [31:0] \u0.u_mmu.fetch_out_pc_o ;
  wire \u0.u_mmu.fetch_out_rd_o ;
  wire \u0.u_mmu.fetch_out_valid_i ;
  wire \u0.u_mmu.lsu_in_accept_o ;
  wire \u0.u_mmu.lsu_in_ack_o ;
  wire [31:0] \u0.u_mmu.lsu_in_addr_i ;
  wire \u0.u_mmu.lsu_in_cacheable_i ;
  wire [31:0] \u0.u_mmu.lsu_in_data_rd_o ;
  wire [31:0] \u0.u_mmu.lsu_in_data_wr_i ;
  wire \u0.u_mmu.lsu_in_error_o ;
  wire \u0.u_mmu.lsu_in_flush_i ;
  wire \u0.u_mmu.lsu_in_invalidate_i ;
  wire \u0.u_mmu.lsu_in_load_fault_o ;
  wire \u0.u_mmu.lsu_in_rd_i ;
  wire [10:0] \u0.u_mmu.lsu_in_req_tag_i ;
  wire [10:0] \u0.u_mmu.lsu_in_resp_tag_o ;
  wire \u0.u_mmu.lsu_in_store_fault_o ;
  wire [3:0] \u0.u_mmu.lsu_in_wr_i ;
  wire \u0.u_mmu.lsu_in_writeback_i ;
  wire \u0.u_mmu.lsu_out_accept_i ;
  wire \u0.u_mmu.lsu_out_ack_i ;
  wire [31:0] \u0.u_mmu.lsu_out_addr_o ;
  wire \u0.u_mmu.lsu_out_cacheable_o ;
  wire [31:0] \u0.u_mmu.lsu_out_data_rd_i ;
  wire [31:0] \u0.u_mmu.lsu_out_data_wr_o ;
  wire \u0.u_mmu.lsu_out_error_i ;
  wire \u0.u_mmu.lsu_out_flush_o ;
  wire \u0.u_mmu.lsu_out_invalidate_o ;
  wire \u0.u_mmu.lsu_out_rd_o ;
  wire [10:0] \u0.u_mmu.lsu_out_req_tag_o ;
  wire [10:0] \u0.u_mmu.lsu_out_resp_tag_i ;
  wire [3:0] \u0.u_mmu.lsu_out_wr_o ;
  wire \u0.u_mmu.lsu_out_writeback_o ;
  wire \u0.u_mmu.mxr_i ;
  wire \u0.u_mmu.rst_i ;
  wire [31:0] \u0.u_mmu.satp_i ;
  wire \u0.u_mmu.sum_i ;
  wire \u0.u_mul.clk_i ;
  wire \u0.u_mul.hold_i ;
  reg \u0.u_mul.mulhi_sel_e1_q ;
  wire \u0.u_mul.mult_inst_w ;
  wire [63:0] \u0.u_mul.mult_result_w ;
  wire \u0.u_mul.opcode_invalid_i ;
  wire [31:0] \u0.u_mul.opcode_opcode_i ;
  wire [31:0] \u0.u_mul.opcode_pc_i ;
  wire [4:0] \u0.u_mul.opcode_ra_idx_i ;
  wire [31:0] \u0.u_mul.opcode_ra_operand_i ;
  wire [4:0] \u0.u_mul.opcode_rb_idx_i ;
  wire [31:0] \u0.u_mul.opcode_rb_operand_i ;
  wire [4:0] \u0.u_mul.opcode_rd_idx_i ;
  wire \u0.u_mul.opcode_valid_i ;
  reg [32:0] \u0.u_mul.operand_a_e1_q ;
  wire [32:0] \u0.u_mul.operand_a_r ;
  reg [32:0] \u0.u_mul.operand_b_e1_q ;
  wire [32:0] \u0.u_mul.operand_b_r ;
  reg [31:0] \u0.u_mul.result_e2_q ;
  wire [31:0] \u0.u_mul.result_r ;
  wire \u0.u_mul.rst_i ;
  wire [31:0] \u0.u_mul.writeback_value_o ;
  wire \u0.writeback_div_valid_w ;
  wire [31:0] \u0.writeback_div_value_w ;
  wire [31:0] \u0.writeback_exec_value_w ;
  wire [5:0] \u0.writeback_mem_exception_w ;
  wire \u0.writeback_mem_valid_w ;
  wire [31:0] \u0.writeback_mem_value_w ;
  wire [31:0] \u0.writeback_mul_value_w ;
  wire wr_d_addr;
  wire wr_d_data_wr;
  wire wr_d_rd;
  wire wr_i_rd;
  wire wri_rd;
  assign _0000_ = 1'h0 == 1'h0;
  assign _0001_ = 1'h1 == 1'h0;
  assign _0002_ = _1197_ == 1'h0;
  assign _0003_ = 1'h0 == 1'h1;
  assign _0004_ = 1'h1 == 1'h1;
  assign _0005_ = _1197_ == 1'h1;
  always @(posedge clk_i)
    \fifo_d_addr.r0  <= _0006_;
  always @(posedge clk_i)
    \fifo_d_addr.r1  <= _0007_;
  assign _0008_ = \fifo_d_addr.wr  ? \fifo_d_addr.r0  : \fifo_d_addr.r1 ;
  assign _0007_ = rst_i ? 32'h00000000 : _0008_;
  assign _0009_ = \fifo_d_addr.wr  ? 32'h00000000 : \fifo_d_addr.r0 ;
  assign _0006_ = rst_i ? 32'h00000000 : _0009_;
  always @(posedge clk_i)
    \fifo_d_data_wr.r0  <= _0010_;
  always @(posedge clk_i)
    \fifo_d_data_wr.r1  <= _0011_;
  assign _0012_ = \u0.u_lsu.mem_wr_o [0] ? \fifo_d_data_wr.r0  : \fifo_d_data_wr.r1 ;
  assign _0011_ = rst_i ? 32'h00000000 : _0012_;
  assign _0013_ = \u0.u_lsu.mem_wr_o [0] ? { 31'h00000000, \u0.u_lsu.mem_data_wr_q [0] } : \fifo_d_data_wr.r0 ;
  assign _0010_ = rst_i ? 32'h00000000 : _0013_;
  always @(posedge clk_i)
    \fifo_d_rd.r0  <= _0014_;
  always @(posedge clk_i)
    \fifo_d_rd.r1  <= _0015_;
  assign _0016_ = \fifo_d_rd.in  ? \fifo_d_rd.r0  : \fifo_d_rd.r1 ;
  assign _0015_ = rst_i ? 1'h0 : _0016_;
  assign _0017_ = \fifo_d_rd.in  ? \fifo_d_rd.in  : \fifo_d_rd.r0 ;
  assign _0014_ = rst_i ? 1'h0 : _0017_;
  always @(posedge clk_i)
    \fifo_d_wr.r0  <= _0018_;
  always @(posedge clk_i)
    \fifo_d_wr.r1  <= _0019_;
  assign _0020_ = \u0.u_lsu.mem_wr_o [0] ? \fifo_d_wr.r0  : \fifo_d_wr.r1 ;
  assign _0019_ = rst_i ? 4'h0 : _0020_;
  assign _0021_ = \u0.u_lsu.mem_wr_o [0] ? { 3'h0, \u0.u_lsu.mem_wr_o [0] } : \fifo_d_wr.r0 ;
  assign _0018_ = rst_i ? 4'h0 : _0021_;
  always @(posedge clk_i)
    \fifo_i_pc.r0  <= _0022_;
  always @(posedge clk_i)
    \fifo_i_pc.r1  <= _0023_;
  assign _0024_ = \fifo_i_pc.wr  ? \fifo_i_pc.r0  : \fifo_i_pc.r1 ;
  assign _0023_ = rst_i ? 32'h00000000 : _0024_;
  assign _0025_ = \fifo_i_pc.wr  ? 32'h00000000 : \fifo_i_pc.r0 ;
  assign _0022_ = rst_i ? 32'h00000000 : _0025_;
  always @(posedge clk_i)
    \fifo_i_rd.r0  <= _0026_;
  always @(posedge clk_i)
    \fifo_i_rd.r1  <= _0027_;
  assign _0028_ = \fifo_i_rd.in  ? \fifo_i_rd.r0  : \fifo_i_rd.r1 ;
  assign _0027_ = rst_i ? 1'h0 : _0028_;
  assign _0029_ = \fifo_i_rd.in  ? \fifo_i_rd.in  : \fifo_i_rd.r0 ;
  assign _0026_ = rst_i ? 1'h0 : _0029_;
  assign _0038_ = 5'h18 + { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] };
  assign _0039_ = \u0.u_csr.opcode_opcode_i  & 15'h707f;
  assign _0040_ = \u0.u_csr.opcode_opcode_i  & 32'hfe007fff;
  assign _0041_ = \u0.u_csr.opcode_opcode_i  & 32'hffffffff;
  assign _0042_ = \u0.u_csr.opcode_opcode_i  & 32'hdfffffff;
  assign _0043_ = \u0.u_csr.csr_rdata_w  & _0064_;
  assign _0044_ = _0089_ & _0065_;
  assign _0045_ = _0039_ == 13'h1073;
  assign _0046_ = _0039_ == 14'h2073;
  assign _0047_ = _0039_ == 14'h3073;
  assign _0048_ = _0039_ == 15'h5073;
  assign _0049_ = _0039_ == 15'h6073;
  assign _0050_ = _0039_ == 15'h7073;
  assign _0051_ = _0040_ == 29'h12000073;
  assign _0052_ = _0039_ == 13'h100f;
  assign _0053_ = \u0.u_csr.opcode_opcode_i [31:20] == 9'h180;
  assign _0054_ = _0041_ == 7'h73;
  assign _0055_ = _0042_ == 29'h10200073;
  assign _0056_ = _0041_ == 21'h100073;
  assign \u0.u_csr.csrrw_w  = \u0.u_csr.opcode_valid_i  && _0045_;
  assign \u0.u_csr.csrrs_w  = \u0.u_csr.opcode_valid_i  && _0046_;
  assign \u0.u_csr.csrrc_w  = \u0.u_csr.opcode_valid_i  && _0047_;
  assign \u0.u_csr.csrrwi_w  = \u0.u_csr.opcode_valid_i  && _0048_;
  assign \u0.u_csr.csrrsi_w  = \u0.u_csr.opcode_valid_i  && _0049_;
  assign \u0.u_csr.csrrci_w  = \u0.u_csr.opcode_valid_i  && _0050_;
  assign \u0.u_csr.sfence_w  = \u0.u_csr.opcode_valid_i  && _0051_;
  assign \u0.u_csr.ifence_w  = \u0.u_csr.opcode_valid_i  && _0052_;
  assign _0057_ = \u0.u_csr.opcode_valid_i  && _0059_;
  assign _0058_ = _0057_ && \u0.u_csr.csr_write_r ;
  assign \u0.u_csr.satp_update_w  = _0058_ && _0053_;
  assign _0060_ = \u0.u_csr.set_r  && \u0.u_csr.clr_r ;
  assign _0059_ = \u0.u_csr.set_r  || \u0.u_csr.clr_r ;
  assign _0061_ = \u0.u_csr.satp_update_w  || \u0.u_csr.ifence_w ;
  assign _0062_ = _0061_ || \u0.u_csr.sfence_w ;
  assign _0063_ = | \u0.u_csr.opcode_opcode_i [19:15];
  assign _0064_ = ~ \u0.u_csr.data_r ;
  assign _0065_ = ~ \u0.u_csr.interrupt_inhibit_i ;
  assign _0066_ = \u0.u_csr.csrrw_w  | \u0.u_csr.csrrs_w ;
  assign _0067_ = _0066_ | \u0.u_csr.csrrwi_w ;
  assign \u0.u_csr.set_r  = _0067_ | \u0.u_csr.csrrsi_w ;
  assign _0068_ = \u0.u_csr.csrrw_w  | \u0.u_csr.csrrc_w ;
  assign _0069_ = _0068_ | \u0.u_csr.csrrwi_w ;
  assign \u0.u_csr.clr_r  = _0069_ | \u0.u_csr.csrrci_w ;
  assign _0070_ = _0063_ | \u0.u_csr.csrrw_w ;
  assign \u0.u_csr.csr_write_r  = _0070_ | \u0.u_csr.csrrwi_w ;
  assign _0071_ = \u0.u_csr.csrrwi_w  | \u0.u_csr.csrrsi_w ;
  assign _0072_ = _0071_ | \u0.u_csr.csrrci_w ;
  assign _0073_ = \u0.u_csr.csr_rdata_w  | \u0.u_csr.data_r ;
  always @(posedge clk_i)
    \u0.u_csr.branch_q  <= _0030_;
  always @(posedge clk_i)
    \u0.u_csr.branch_target_q  <= _0031_;
  always @(posedge clk_i)
    \u0.u_csr.reset_q  <= _0036_;
  always @(posedge clk_i)
    \u0.u_csr.take_interrupt_q  <= _0037_;
  always @(posedge clk_i)
    \u0.u_csr.rd_valid_e1_q  <= _0035_;
  always @(posedge clk_i)
    \u0.u_csr.rd_result_e1_q  <= _0034_;
  always @(posedge clk_i)
    \u0.u_csr.csr_wdata_e1_q  <= _0032_;
  always @(posedge clk_i)
    \u0.u_csr.exception_e1_q  <= _0033_;
  assign _0074_ = \u0.u_csr.reset_q  ? 1'h1 : \u0.u_csr.csr_branch_w ;
  assign _0030_ = rst_i ? 1'h0 : _0074_;
  assign _0075_ = \u0.u_csr.reset_q  ? reset_vector_i : \u0.u_csr.csr_target_w ;
  assign _0031_ = rst_i ? 32'h00000000 : _0075_;
  assign _0036_ = rst_i ? 1'h1 : 1'h0;
  assign _0037_ = rst_i ? 1'h0 : _0044_;
  assign _0076_ = _0062_ ? 6'h31 : 6'h00;
  assign _0077_ = \u0.u_csr.opcode_invalid_i  ? 6'h12 : _0076_;
  assign _0078_ = _0056_ ? 6'h13 : _0077_;
  assign _0079_ = _0055_ ? 6'h30 : _0078_;
  assign _0080_ = _0054_ ? _0038_ : _0079_;
  assign _0081_ = \u0.u_csr.opcode_valid_i  ? _0080_ : 6'h00;
  assign _0033_ = rst_i ? 6'h00 : _0081_;
  assign _0082_ = \u0.u_csr.opcode_invalid_i  ? \u0.u_csr.opcode_opcode_i  : \u0.u_csr.csr_rdata_w ;
  assign _0083_ = \u0.u_csr.opcode_valid_i  ? _0082_ : 32'h00000000;
  assign _0034_ = rst_i ? 32'h00000000 : _0083_;
  assign _0084_ = \u0.u_csr.opcode_valid_i  ? _0059_ : 1'h0;
  assign _0035_ = rst_i ? 1'h0 : _0084_;
  assign _0085_ = \u0.u_csr.clr_r  ? _0043_ : \u0.u_csr.csr_wdata_e1_q ;
  assign _0086_ = \u0.u_csr.set_r  ? _0073_ : _0085_;
  assign _0087_ = _0060_ ? \u0.u_csr.data_r  : _0086_;
  assign _0088_ = \u0.u_csr.opcode_valid_i  ? _0087_ : 32'h00000000;
  assign _0032_ = rst_i ? 32'h00000000 : _0088_;
  assign _0089_ = | \u0.u_csr.interrupt_w ;
  assign \u0.u_csr.data_r  = _0072_ ? { 27'h0000000, \u0.u_csr.opcode_opcode_i [19:15] } : \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_csr.u_csrfile.csr_waddr_i  = \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q  ? \u0.u_issue.u_pipe_ctrl.opcode_wb_q [31:20] : 12'h000;
  assign \u0.u_csr.u_csrfile.csr_mcycle_r  = \u0.u_csr.u_csrfile.csr_mcycle_q  + 1'h1;
  assign _0161_ = \u0.u_issue.u_pipe_ctrl.pc_wb_q  + 3'h4;
  assign \u0.u_csr.u_csrfile.irq_pending_r  = \u0.u_csr.u_csrfile.csr_mip_q  & \u0.u_csr.u_csrfile.csr_mie_q ;
  assign _0162_ = \u0.u_csr.u_csrfile.csr_mscratch_q  & 32'hffffffff;
  assign _0163_ = \u0.u_csr.u_csrfile.csr_mepc_q  & 32'hffffffff;
  assign _0164_ = \u0.u_csr.u_csrfile.csr_mtvec_q  & 32'hffffffff;
  assign _0165_ = \u0.u_csr.u_csrfile.csr_mcause_q  & 32'h8000000f;
  assign _0166_ = \u0.u_csr.u_csrfile.csr_mtval_q  & 32'hffffffff;
  assign _0167_ = \u0.u_csr.u_csrfile.csr_sr_q  & 32'hffffffff;
  assign _0168_ = \u0.u_csr.u_csrfile.csr_mip_q  & 12'haaa;
  assign _0169_ = \u0.u_csr.u_csrfile.csr_mie_q  & 12'haaa;
  assign _0170_ = \u0.u_issue.u_pipe_ctrl.exception_wb_q  & 6'h30;
  assign _0171_ = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  & 32'hffffffff;
  assign _0172_ = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  & 32'h8000000f;
  assign _0173_ = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  & 12'haaa;
  assign _0174_ = \u0.u_csr.u_csrfile.csr_sr_q  & 32'hfffbfecc;
  assign _0175_ = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  & 19'h40133;
  assign _0176_ = \u0.u_csr.u_csrfile.csr_mip_q  & 32'hfffffddd;
  assign _0177_ = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  & 10'h222;
  assign _0178_ = \u0.u_csr.u_csrfile.csr_mie_q  & 32'hfffffddd;
  assign _0179_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h344;
  assign _0180_ = \u0.u_csr.opcode_opcode_i [31:20] == 9'h144;
  assign _0181_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h344;
  assign _0182_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 9'h144;
  assign \u0.u_csr.u_csrfile.is_exception_w  = _0170_ == 5'h10;
  assign _0183_ = _0170_ == 6'h20;
  assign _0184_ = \u0.u_csr.u_csrfile.irq_priv_q  == 2'h3;
  assign _0185_ = { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] } == 1'h1;
  assign _0186_ = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 6'h30;
  assign _0187_ = { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] } == 2'h3;
  assign _0188_ = \u0.u_csr.u_csrfile.csr_mcycle_q  == \u0.u_csr.u_csrfile.csr_mtimecmp_q ;
  assign _0189_ = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 6'h20;
  assign _0190_ = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 6'h31;
  assign _0191_ = \u0.u_csr.opcode_valid_i  && _0179_;
  assign _0192_ = \u0.u_csr.opcode_valid_i  && _0180_;
  assign _0193_ = $signed(32'h00000001) && _0188_;
  assign _0194_ = _0191_ || _0192_;
  assign _0195_ = _0181_ || _0182_;
  assign _0196_ = _0195_ || _0231_;
  assign _0197_ = _0191_ | _0192_;
  assign \u0.u_csr.u_csrfile.buffer_mip_w  = _0197_ | \u0.u_csr.u_csrfile.csr_mip_upd_q ;
  assign _0198_ = _0174_ | _0175_;
  assign _0199_ = _0176_ | _0177_;
  assign _0200_ = _0178_ | _0177_;
  assign \u0.u_csr.u_csrfile.csr_mip_r  = _0109_ | { \u0.u_csr.u_csrfile.csr_mip_next_q [31:12], \u0.u_csr.u_csrfile.csr_mip_next_r [11], \u0.u_csr.u_csrfile.csr_mip_next_q [10:8], \u0.u_csr.u_csrfile.csr_mip_next_r [7], \u0.u_csr.u_csrfile.csr_mip_next_q [6:0] };
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mepc_q  <= _0092_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mcause_q  <= _0090_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_sr_q  <= _0102_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mtvec_q  <= _0101_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mip_q  <= _0095_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mie_q  <= _0093_;
  reg \u0.u_csr.u_csrfile.csr_mpriv_q_reg[0] ;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mpriv_q_reg[0]  <= 1'h1;
  assign \u0.u_csr.u_csrfile.csr_mpriv_q [0] = \u0.u_csr.u_csrfile.csr_mpriv_q_reg[0] ;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mcycle_q  <= _0091_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mscratch_q  <= _0097_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mtval_q  <= _0100_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mtimecmp_q  <= _0099_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mtime_ie_q  <= _0098_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mip_next_q  <= _0094_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.csr_mip_upd_q  <= _0096_;
  always @(posedge clk_i)
    \u0.u_csr.u_csrfile.irq_priv_q  <= _0103_;
  assign _0150_ = _0190_ ? _0161_ : 32'h00000000;
  assign _0149_ = _0190_ ? 1'h1 : 1'h0;
  assign _0135_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mtvec_q  : _0150_;
  assign _0134_ = \u0.u_csr.u_csrfile.is_exception_w  ? 1'h1 : _0149_;
  assign _0123_ = _0187_ ? \u0.u_csr.u_csrfile.csr_mepc_q  : 32'h00000000;
  assign _0112_ = _0186_ ? _0123_ : _0135_;
  assign _0111_ = _0186_ ? 1'h1 : _0134_;
  assign \u0.u_csr.csr_target_w  = _0189_ ? _0233_ : _0112_;
  assign \u0.u_csr.csr_branch_w  = _0189_ ? 1'h1 : _0111_;
  assign _0094_ = rst_i ? 32'h00000000 : _0232_;
  assign _0098_ = rst_i ? 1'h0 : \u0.u_csr.u_csrfile.csr_mtime_ie_r ;
  assign _0099_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mtimecmp_r ;
  assign _0097_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mscratch_r ;
  assign _0091_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mcycle_r ;
  assign _0093_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mie_r ;
  assign _0095_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mip_r ;
  assign _0101_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mtvec_r ;
  assign _0100_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mtval_r ;
  assign _0090_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mcause_r ;
  assign _0102_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_sr_r ;
  assign _0092_ = rst_i ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mepc_r ;
  assign \u0.u_csr.u_csrfile.csr_mtime_ie_r  = _0193_ ? 1'h0 : _0110_;
  assign \u0.u_csr.u_csrfile.csr_mip_next_r [7] = _0193_ ? \u0.u_csr.u_csrfile.csr_mtime_ie_q  : _0138_;
  assign _0138_ = 1'h0 ? 1'h1 : \u0.u_csr.u_csrfile.csr_mip_next_q [7];
  assign \u0.u_csr.u_csrfile.csr_mip_next_r [11] = intr_i ? 1'h1 : \u0.u_csr.u_csrfile.csr_mip_next_q [11];
  assign _0144_ = _0201_ ? _0171_ : \u0.u_csr.u_csrfile.csr_mscratch_q ;
  assign _0201_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h340;
  assign _0145_ = _0202_ ? 1'h1 : \u0.u_csr.u_csrfile.csr_mtime_ie_q ;
  assign _0202_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 11'h7c0;
  assign _0146_ = _0202_ ? _0171_ : \u0.u_csr.u_csrfile.csr_mtimecmp_q ;
  function [31:0] _1468_;
    input [31:0] a;
    input [63:0] b;
    input [1:0] s;
    casez (s) // synopsys parallel_case
      2'b?1:
        _1468_ = b[31:0];
      2'b1?:
        _1468_ = b[63:32];
      default:
        _1468_ = a;
    endcase
  endfunction
  assign _0142_ = _1468_(\u0.u_csr.u_csrfile.csr_mie_q , { _0173_, _0200_ }, { _0204_, _0203_ });
  assign _0203_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 9'h104;
  assign _0204_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h304;
  function [31:0] _1471_;
    input [31:0] a;
    input [63:0] b;
    input [1:0] s;
    casez (s) // synopsys parallel_case
      2'b?1:
        _1471_ = b[31:0];
      2'b1?:
        _1471_ = b[63:32];
      default:
        _1471_ = a;
    endcase
  endfunction
  assign _0143_ = _1471_(\u0.u_csr.u_csrfile.csr_mip_q , { _0173_, _0199_ }, { _0181_, _0182_ });
  assign _0147_ = _0205_ ? _0171_ : \u0.u_csr.u_csrfile.csr_mtvec_q ;
  assign _0205_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h305;
  function [31:0] _1474_;
    input [31:0] a;
    input [63:0] b;
    input [1:0] s;
    casez (s) // synopsys parallel_case
      2'b?1:
        _1474_ = b[31:0];
      2'b1?:
        _1474_ = b[63:32];
      default:
        _1474_ = a;
    endcase
  endfunction
  assign _0108_ = _1474_(\u0.u_csr.u_csrfile.csr_sr_q , { _0171_, _0198_ }, { _0207_, _0206_ });
  assign _0206_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 9'h100;
  assign _0207_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h300;
  assign _0156_ = _0208_ ? _0171_ : \u0.u_csr.u_csrfile.csr_mtval_q ;
  assign _0208_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h343;
  assign _0159_ = _0209_ ? _0172_ : \u0.u_csr.u_csrfile.csr_mcause_q ;
  assign _0209_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h342;
  assign _0152_ = _0210_ ? _0171_ : \u0.u_csr.u_csrfile.csr_mepc_q ;
  assign _0210_ = \u0.u_csr.u_csrfile.csr_waddr_i  == 10'h341;
  assign _0107_[31:13] = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_sr_q [31:13] : _0108_[31:13];
  assign _0107_[10:8] = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_sr_q [10:8] : _0108_[10:8];
  assign _0107_[6:4] = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_sr_q [6:4] : _0108_[6:4];
  assign _0107_[2:0] = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_sr_q [2:0] : _0108_[2:0];
  assign _0155_ = \u0.u_csr.u_csrfile.is_exception_w  ? { 28'h0000000, \u0.u_issue.u_pipe_ctrl.exception_wb_q [3:0] } : _0159_;
  assign _0139_ = \u0.u_csr.u_csrfile.is_exception_w  ? _0153_ : _0156_;
  assign _0137_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_issue.u_pipe_ctrl.pc_wb_q  : _0152_;
  assign _0107_[3] = \u0.u_csr.u_csrfile.is_exception_w  ? 1'h0 : _0108_[3];
  assign _0107_[12:11] = \u0.u_csr.u_csrfile.is_exception_w  ? { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] } : _0108_[12:11];
  assign _0107_[7] = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_sr_q [3] : _0108_[7];
  assign _0129_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mtime_ie_q  : _0145_;
  assign _0130_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mtimecmp_q  : _0146_;
  assign _0128_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mscratch_q  : _0144_;
  assign _0126_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mie_q  : _0142_;
  assign _0127_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mip_q  : _0143_;
  assign _0132_ = \u0.u_csr.u_csrfile.is_exception_w  ? \u0.u_csr.u_csrfile.csr_mtvec_q  : _0147_;
  function [31:0] _1499_;
    input [31:0] a;
    input [63:0] b;
    input [1:0] s;
    casez (s) // synopsys parallel_case
      2'b?1:
        _1499_ = b[31:0];
      2'b1?:
        _1499_ = b[63:32];
      default:
        _1499_ = a;
    endcase
  endfunction
  assign _0153_ = _1499_(32'h00000000, { \u0.u_issue.u_pipe_ctrl.pc_wb_q , \u0.u_issue.u_pipe_ctrl.result_wb_q  }, { _0214_, _0212_ });
  assign _0212_ = | _0211_;
  assign _0211_[0] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h12;
  assign _0211_[1] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h14;
  assign _0211_[2] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h15;
  assign _0211_[3] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h16;
  assign _0211_[4] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h17;
  assign _0211_[5] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h1d;
  assign _0211_[6] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h1f;
  assign _0214_ = | _0213_;
  assign _0213_[0] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h10;
  assign _0213_[1] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h11;
  assign _0213_[2] = \u0.u_issue.u_pipe_ctrl.exception_wb_q  == 5'h1c;
  assign _0157_[31:13] = _0186_ ? \u0.u_csr.u_csrfile.csr_sr_q [31:13] : _0107_[31:13];
  assign _0157_[10:9] = _0186_ ? \u0.u_csr.u_csrfile.csr_sr_q [10:9] : _0107_[10:9];
  assign _0157_[6] = _0186_ ? \u0.u_csr.u_csrfile.csr_sr_q [6] : _0107_[6];
  assign _0157_[4] = _0186_ ? \u0.u_csr.u_csrfile.csr_sr_q [4] : _0107_[4];
  assign _0157_[2] = _0186_ ? \u0.u_csr.u_csrfile.csr_sr_q [2] : _0107_[2];
  assign _0157_[0] = _0186_ ? \u0.u_csr.u_csrfile.csr_sr_q [0] : _0107_[0];
  assign _0105_[0] = _0187_ ? 1'h1 : \u0.u_csr.u_csrfile.csr_sr_q [7];
  assign _0160_ = _0187_ ? \u0.u_csr.u_csrfile.csr_sr_q [7] : \u0.u_csr.u_csrfile.csr_sr_q [3];
  assign _0105_[1] = _0187_ ? \u0.u_csr.u_csrfile.csr_sr_q [8] : 1'h0;
  assign _0104_ = _0187_ ? \u0.u_csr.u_csrfile.csr_sr_q [5] : 1'h1;
  assign _0158_ = _0187_ ? \u0.u_csr.u_csrfile.csr_sr_q [1] : \u0.u_csr.u_csrfile.csr_sr_q [5];
  assign _0157_[12:11] = _0186_ ? _0106_ : _0107_[12:11];
  assign _0157_[8:7] = _0186_ ? _0105_ : _0107_[8:7];
  assign _0157_[5] = _0186_ ? _0104_ : _0107_[5];
  assign _0157_[3] = _0186_ ? _0160_ : _0107_[3];
  assign _0157_[1] = _0186_ ? _0158_ : _0107_[1];
  assign _0118_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mtime_ie_q  : _0129_;
  assign _0119_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mtimecmp_q  : _0130_;
  assign _0117_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mscratch_q  : _0128_;
  assign _0115_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mie_q  : _0126_;
  assign _0116_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mip_q  : _0127_;
  assign _0121_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mtvec_q  : _0132_;
  assign _0106_ = _0187_ ? 2'h0 : \u0.u_csr.u_csrfile.csr_sr_q [12:11];
  assign _0131_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mtval_q  : _0139_;
  assign _0151_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mcause_q  : _0155_;
  assign _0125_ = _0186_ ? \u0.u_csr.u_csrfile.csr_mepc_q  : _0137_;
  assign \u0.u_csr.u_csrfile.csr_sr_r [31:13] = _0183_ ? \u0.u_csr.u_csrfile.csr_sr_q [31:13] : _0157_[31:13];
  assign \u0.u_csr.u_csrfile.csr_sr_r [10:9] = _0183_ ? \u0.u_csr.u_csrfile.csr_sr_q [10:9] : _0157_[10:9];
  assign \u0.u_csr.u_csrfile.csr_sr_r [6] = _0183_ ? \u0.u_csr.u_csrfile.csr_sr_q [6] : _0157_[6];
  assign \u0.u_csr.u_csrfile.csr_sr_r [4] = _0183_ ? \u0.u_csr.u_csrfile.csr_sr_q [4] : _0157_[4];
  assign \u0.u_csr.u_csrfile.csr_sr_r [2] = _0183_ ? \u0.u_csr.u_csrfile.csr_sr_q [2] : _0157_[2];
  assign \u0.u_csr.u_csrfile.csr_sr_r [0] = _0183_ ? \u0.u_csr.u_csrfile.csr_sr_q [0] : _0157_[0];
  assign _0141_ = \u0.u_csr.interrupt_w [11] ? 32'h8000000b : \u0.u_csr.u_csrfile.csr_mcause_q ;
  assign _0136_ = \u0.u_csr.interrupt_w [7] ? 32'h80000007 : _0141_;
  assign _0124_ = \u0.u_csr.interrupt_w [3] ? 32'h80000003 : _0136_;
  assign _0113_ = _0184_ ? _0124_ : \u0.u_csr.u_csrfile.csr_mcause_q ;
  assign _0120_ = _0184_ ? 32'h00000000 : \u0.u_csr.u_csrfile.csr_mtval_q ;
  assign _0114_ = _0184_ ? \u0.u_issue.u_pipe_ctrl.pc_wb_q  : \u0.u_csr.u_csrfile.csr_mepc_q ;
  assign _0133_ = _0184_ ? 1'h0 : \u0.u_csr.u_csrfile.csr_sr_q [3];
  assign _0154_ = _0184_ ? { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] } : \u0.u_csr.u_csrfile.csr_sr_q [12:11];
  assign _0148_[0] = _0184_ ? \u0.u_csr.u_csrfile.csr_sr_q [3] : \u0.u_csr.u_csrfile.csr_sr_q [7];
  assign _0148_[1] = _0184_ ? \u0.u_csr.u_csrfile.csr_sr_q [8] : _0185_;
  assign _0140_ = _0184_ ? \u0.u_csr.u_csrfile.csr_sr_q [5] : \u0.u_csr.u_csrfile.csr_sr_q [1];
  assign _0122_ = _0184_ ? \u0.u_csr.u_csrfile.csr_sr_q [1] : 1'h0;
  assign \u0.u_csr.u_csrfile.csr_sr_r [12:11] = _0183_ ? _0154_ : _0157_[12:11];
  assign \u0.u_csr.u_csrfile.csr_sr_r [8:7] = _0183_ ? _0148_ : _0157_[8:7];
  assign \u0.u_csr.u_csrfile.csr_sr_r [5] = _0183_ ? _0140_ : _0157_[5];
  assign \u0.u_csr.u_csrfile.csr_sr_r [3] = _0183_ ? _0133_ : _0157_[3];
  assign \u0.u_csr.u_csrfile.csr_sr_r [1] = _0183_ ? _0122_ : _0157_[1];
  assign \u0.u_csr.u_csrfile.csr_mtval_r  = _0183_ ? _0120_ : _0131_;
  assign \u0.u_csr.u_csrfile.csr_mcause_r  = _0183_ ? _0113_ : _0151_;
  assign \u0.u_csr.u_csrfile.csr_mepc_r  = _0183_ ? _0114_ : _0125_;
  assign _0110_ = _0183_ ? \u0.u_csr.u_csrfile.csr_mtime_ie_q  : _0118_;
  assign \u0.u_csr.u_csrfile.csr_mtimecmp_r  = _0183_ ? \u0.u_csr.u_csrfile.csr_mtimecmp_q  : _0119_;
  assign \u0.u_csr.u_csrfile.csr_mscratch_r  = _0183_ ? \u0.u_csr.u_csrfile.csr_mscratch_q  : _0117_;
  assign \u0.u_csr.u_csrfile.csr_mie_r  = _0183_ ? \u0.u_csr.u_csrfile.csr_mie_q  : _0115_;
  assign _0109_ = _0183_ ? \u0.u_csr.u_csrfile.csr_mip_q  : _0116_;
  assign \u0.u_csr.u_csrfile.csr_mtvec_r  = _0183_ ? \u0.u_csr.u_csrfile.csr_mtvec_q  : _0121_;
  function [31:0] _1570_;
    input [31:0] a;
    input [383:0] b;
    input [11:0] s;
    casez (s) // synopsys parallel_case
      12'b???????????1:
        _1570_ = b[31:0];
      12'b??????????1?:
        _1570_ = b[63:32];
      12'b?????????1??:
        _1570_ = b[95:64];
      12'b????????1???:
        _1570_ = b[127:96];
      12'b???????1????:
        _1570_ = b[159:128];
      12'b??????1?????:
        _1570_ = b[191:160];
      12'b?????1??????:
        _1570_ = b[223:192];
      12'b????1???????:
        _1570_ = b[255:224];
      12'b???1????????:
        _1570_ = b[287:256];
      12'b??1?????????:
        _1570_ = b[319:288];
      12'b?1??????????:
        _1570_ = b[351:320];
      12'b1???????????:
        _1570_ = b[383:352];
      default:
        _1570_ = a;
    endcase
  endfunction
  assign \u0.u_csr.csr_rdata_w  = _1570_(32'h00000000, { _0162_, _0163_, _0164_, _0165_, _0166_, _0167_, _0168_, _0169_, \u0.u_csr.u_csrfile.csr_mcycle_q , cpu_id_i, 32'h40001100, \u0.u_csr.u_csrfile.csr_mtimecmp_q  }, { _0226_, _0225_, _0224_, _0223_, _0222_, _0221_, _0179_, _0220_, _0219_, _0217_, _0216_, _0215_ });
  assign _0215_ = \u0.u_csr.opcode_opcode_i [31:20] == 11'h7c0;
  assign _0216_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h301;
  assign _0217_ = \u0.u_csr.opcode_opcode_i [31:20] == 12'hf14;
  assign _0219_ = | _0218_;
  assign _0218_[0] = \u0.u_csr.opcode_opcode_i [31:20] == 12'hc00;
  assign _0218_[1] = \u0.u_csr.opcode_opcode_i [31:20] == 12'hc01;
  assign _0220_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h304;
  assign _0221_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h300;
  assign _0222_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h343;
  assign _0223_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h342;
  assign _0224_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h305;
  assign _0225_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h341;
  assign _0226_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h340;
  assign _0227_ = _0196_ ? 1'h0 : \u0.u_csr.u_csrfile.csr_mip_upd_q ;
  assign _0228_ = _0194_ ? 1'h1 : _0227_;
  assign _0096_ = rst_i ? 1'h0 : _0228_;
  assign _0229_ = _0230_ ? 2'h3 : \u0.u_csr.u_csrfile.irq_priv_q ;
  assign _0103_ = rst_i ? 2'h3 : _0229_;
  assign _0230_ = | \u0.u_csr.interrupt_w ;
  assign _0231_ = | \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.u_csr.interrupt_w  = \u0.u_csr.u_csrfile.csr_sr_q [3] ? \u0.u_csr.u_csrfile.irq_pending_r  : 32'h00000000;
  assign _0232_ = \u0.u_csr.u_csrfile.buffer_mip_w  ? { \u0.u_csr.u_csrfile.csr_mip_next_q [31:12], \u0.u_csr.u_csrfile.csr_mip_next_r [11], \u0.u_csr.u_csrfile.csr_mip_next_q [10:8], \u0.u_csr.u_csrfile.csr_mip_next_r [7], \u0.u_csr.u_csrfile.csr_mip_next_q [6:0] } : 32'h00000000;
  assign _0233_ = _0184_ ? \u0.u_csr.u_csrfile.csr_mtvec_q  : 32'h00000000;
  assign \u0.u_decode.genblk1.u_dec.fetch_fault_i  = \u0.u_decode.fetch_in_fault_page_i  | \u0.u_decode.fetch_in_fault_fetch_i ;
  assign \u0.u_csr.opcode_opcode_i  = \u0.u_decode.genblk1.u_dec.fetch_fault_i  ? 32'h00000000 : \u0.u_decode.fetch_in_instr_i ;
  assign _0234_ = \u0.u_csr.opcode_opcode_i  & 32'hffffffff;
  assign _0235_ = \u0.u_csr.opcode_opcode_i  & 32'hdfffffff;
  assign _0236_ = \u0.u_csr.opcode_opcode_i  & 15'h707f;
  assign _0237_ = \u0.u_csr.opcode_opcode_i  & 32'hffff8fff;
  assign _0238_ = \u0.u_csr.opcode_opcode_i  & 32'hfe007fff;
  assign _0239_ = \u0.u_csr.opcode_opcode_i  & 32'hfe00707f;
  assign _0240_ = \u0.u_csr.opcode_opcode_i  & 7'h7f;
  assign _0241_ = \u0.u_csr.opcode_opcode_i  & 32'hfc00707f;
  assign _0242_ = _0234_ == 7'h73;
  assign _0243_ = _0234_ == 21'h100073;
  assign _0244_ = _0235_ == 29'h10200073;
  assign _0245_ = _0236_ == 13'h1073;
  assign _0246_ = _0236_ == 14'h2073;
  assign _0247_ = _0236_ == 14'h3073;
  assign _0248_ = _0236_ == 15'h5073;
  assign _0249_ = _0236_ == 15'h6073;
  assign _0250_ = _0236_ == 15'h7073;
  assign _0251_ = _0237_ == 29'h10500073;
  assign _0252_ = _0236_ == 4'hf;
  assign _0253_ = _0236_ == 13'h100f;
  assign _0254_ = _0238_ == 29'h12000073;
  assign _0255_ = _0239_ == 26'h2000033;
  assign _0256_ = _0239_ == 26'h2001033;
  assign _0257_ = _0239_ == 26'h2002033;
  assign _0258_ = _0239_ == 26'h2003033;
  assign _0259_ = _0239_ == 26'h2004033;
  assign _0260_ = _0239_ == 26'h2005033;
  assign _0261_ = _0239_ == 26'h2006033;
  assign _0262_ = _0239_ == 26'h2007033;
  assign _0263_ = _0236_ == 7'h67;
  assign _0264_ = _0240_ == 7'h6f;
  assign _0265_ = _0240_ == 6'h37;
  assign _0266_ = _0240_ == 5'h17;
  assign _0267_ = _0236_ == 5'h13;
  assign _0268_ = _0241_ == 13'h1013;
  assign _0269_ = _0236_ == 14'h2013;
  assign _0270_ = _0236_ == 14'h3013;
  assign _0271_ = _0236_ == 15'h4013;
  assign _0272_ = _0241_ == 15'h5013;
  assign _0273_ = _0241_ == 31'h40005013;
  assign _0274_ = _0236_ == 15'h6013;
  assign _0275_ = _0236_ == 15'h7013;
  assign _0276_ = _0239_ == 6'h33;
  assign _0277_ = _0239_ == 31'h40000033;
  assign _0278_ = _0239_ == 13'h1033;
  assign _0279_ = _0239_ == 14'h2033;
  assign _0280_ = _0239_ == 14'h3033;
  assign _0281_ = _0239_ == 15'h4033;
  assign _0282_ = _0239_ == 15'h5033;
  assign _0283_ = _0239_ == 31'h40005033;
  assign _0284_ = _0239_ == 15'h6033;
  assign _0285_ = _0239_ == 15'h7033;
  assign _0286_ = _0236_ == 2'h3;
  assign _0287_ = _0236_ == 13'h1003;
  assign _0288_ = _0236_ == 14'h2003;
  assign _0289_ = _0236_ == 15'h4003;
  assign _0290_ = _0236_ == 15'h5003;
  assign _0291_ = _0236_ == 15'h6003;
  assign _0292_ = _0236_ == 6'h23;
  assign _0293_ = _0236_ == 13'h1023;
  assign _0294_ = _0236_ == 14'h2023;
  assign _0295_ = _0236_ == 7'h63;
  assign _0296_ = _0236_ == 13'h1063;
  assign _0297_ = _0236_ == 15'h4063;
  assign _0298_ = _0236_ == 15'h5063;
  assign _0299_ = _0236_ == 15'h6063;
  assign _0300_ = _0236_ == 15'h7063;
  assign _0301_ = 1'h1 && _0255_;
  assign _0302_ = 1'h1 && _0256_;
  assign _0303_ = 1'h1 && _0257_;
  assign _0304_ = 1'h1 && _0258_;
  assign _0305_ = 1'h1 && _0259_;
  assign _0306_ = 1'h1 && _0260_;
  assign _0307_ = 1'h1 && _0261_;
  assign _0308_ = 1'h1 && _0262_;
  assign \u0.u_decode.genblk1.u_dec.mul_o  = 1'h1 && _0383_;
  assign \u0.u_decode.genblk1.u_dec.div_o  = 1'h1 && _0386_;
  assign \u0.u_decode.genblk1.u_dec.invalid_w  = \u0.u_decode.genblk1.u_dec.valid_i  && _0438_;
  assign _0309_ = _0263_ || _0264_;
  assign _0310_ = _0309_ || _0265_;
  assign _0311_ = _0310_ || _0266_;
  assign _0312_ = _0311_ || _0267_;
  assign _0313_ = _0312_ || _0268_;
  assign _0314_ = _0313_ || _0269_;
  assign _0315_ = _0314_ || _0270_;
  assign _0316_ = _0315_ || _0271_;
  assign _0317_ = _0316_ || _0272_;
  assign _0318_ = _0317_ || _0273_;
  assign _0319_ = _0318_ || _0274_;
  assign _0320_ = _0319_ || _0275_;
  assign _0321_ = _0320_ || _0276_;
  assign _0322_ = _0321_ || _0277_;
  assign _0323_ = _0322_ || _0278_;
  assign _0324_ = _0323_ || _0279_;
  assign _0325_ = _0324_ || _0280_;
  assign _0326_ = _0325_ || _0281_;
  assign _0327_ = _0326_ || _0282_;
  assign _0328_ = _0327_ || _0283_;
  assign _0329_ = _0328_ || _0284_;
  assign _0330_ = _0329_ || _0285_;
  assign _0331_ = _0330_ || _0286_;
  assign _0332_ = _0331_ || _0287_;
  assign _0333_ = _0332_ || _0288_;
  assign _0334_ = _0333_ || _0289_;
  assign _0335_ = _0334_ || _0290_;
  assign _0336_ = _0335_ || _0291_;
  assign _0337_ = _0336_ || _0255_;
  assign _0338_ = _0337_ || _0256_;
  assign _0339_ = _0338_ || _0257_;
  assign _0340_ = _0339_ || _0258_;
  assign _0341_ = _0340_ || _0259_;
  assign _0342_ = _0341_ || _0260_;
  assign _0343_ = _0342_ || _0261_;
  assign _0344_ = _0343_ || _0262_;
  assign _0345_ = _0344_ || _0245_;
  assign _0346_ = _0345_ || _0246_;
  assign _0347_ = _0346_ || _0247_;
  assign _0348_ = _0347_ || _0248_;
  assign _0349_ = _0348_ || _0249_;
  assign \u0.u_decode.genblk1.u_dec.rd_valid_o  = _0349_ || _0250_;
  assign _0350_ = _0275_ || _0267_;
  assign _0351_ = _0350_ || _0269_;
  assign _0352_ = _0351_ || _0270_;
  assign _0353_ = _0352_ || _0274_;
  assign _0354_ = _0353_ || _0271_;
  assign _0355_ = _0354_ || _0268_;
  assign _0356_ = _0355_ || _0272_;
  assign _0357_ = _0356_ || _0273_;
  assign _0358_ = _0357_ || _0265_;
  assign _0359_ = _0358_ || _0266_;
  assign _0360_ = _0359_ || _0276_;
  assign _0361_ = _0360_ || _0277_;
  assign _0362_ = _0361_ || _0279_;
  assign _0363_ = _0362_ || _0280_;
  assign _0364_ = _0363_ || _0281_;
  assign _0365_ = _0364_ || _0284_;
  assign _0366_ = _0365_ || _0285_;
  assign _0367_ = _0366_ || _0278_;
  assign _0368_ = _0367_ || _0282_;
  assign \u0.u_decode.genblk1.u_dec.exec_o  = _0368_ || _0283_;
  assign _0369_ = _0286_ || _0287_;
  assign _0370_ = _0369_ || _0288_;
  assign _0371_ = _0370_ || _0289_;
  assign _0372_ = _0371_ || _0290_;
  assign _0373_ = _0372_ || _0291_;
  assign _0374_ = _0373_ || _0292_;
  assign _0375_ = _0374_ || _0293_;
  assign \u0.u_decode.genblk1.u_dec.lsu_o  = _0375_ || _0294_;
  assign _0376_ = _0309_ || _0295_;
  assign _0377_ = _0376_ || _0296_;
  assign _0378_ = _0377_ || _0297_;
  assign _0379_ = _0378_ || _0298_;
  assign _0380_ = _0379_ || _0299_;
  assign \u0.u_decode.genblk1.u_dec.branch_o  = _0380_ || _0300_;
  assign _0381_ = _0255_ || _0256_;
  assign _0382_ = _0381_ || _0257_;
  assign _0383_ = _0382_ || _0258_;
  assign _0384_ = _0259_ || _0260_;
  assign _0385_ = _0384_ || _0261_;
  assign _0386_ = _0385_ || _0262_;
  assign _0387_ = _0242_ || _0243_;
  assign _0388_ = _0387_ || _0244_;
  assign _0389_ = _0388_ || _0245_;
  assign _0390_ = _0389_ || _0246_;
  assign _0391_ = _0390_ || _0247_;
  assign _0392_ = _0391_ || _0248_;
  assign _0393_ = _0392_ || _0249_;
  assign _0394_ = _0393_ || _0250_;
  assign _0395_ = _0394_ || _0251_;
  assign _0396_ = _0395_ || _0252_;
  assign _0397_ = _0396_ || _0253_;
  assign _0398_ = _0397_ || _0254_;
  assign _0399_ = _0398_ || \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign \u0.u_decode.genblk1.u_dec.csr_o  = _0399_ || \u0.u_decode.genblk1.u_dec.fetch_fault_i ;
  assign _0400_ = \u0.u_decode.genblk1.u_dec.exec_o  || _0264_;
  assign _0401_ = _0400_ || _0263_;
  assign _0402_ = _0401_ || _0295_;
  assign _0403_ = _0402_ || _0296_;
  assign _0404_ = _0403_ || _0297_;
  assign _0405_ = _0404_ || _0298_;
  assign _0406_ = _0405_ || _0299_;
  assign _0407_ = _0406_ || _0300_;
  assign _0408_ = _0407_ || _0286_;
  assign _0409_ = _0408_ || _0287_;
  assign _0410_ = _0409_ || _0288_;
  assign _0411_ = _0410_ || _0289_;
  assign _0412_ = _0411_ || _0290_;
  assign _0413_ = _0412_ || _0291_;
  assign _0414_ = _0413_ || _0292_;
  assign _0415_ = _0414_ || _0293_;
  assign _0416_ = _0415_ || _0294_;
  assign _0417_ = _0416_ || _0242_;
  assign _0418_ = _0417_ || _0243_;
  assign _0419_ = _0418_ || _0244_;
  assign _0420_ = _0419_ || _0245_;
  assign _0421_ = _0420_ || _0246_;
  assign _0422_ = _0421_ || _0247_;
  assign _0423_ = _0422_ || _0248_;
  assign _0424_ = _0423_ || _0249_;
  assign _0425_ = _0424_ || _0250_;
  assign _0426_ = _0425_ || _0251_;
  assign _0427_ = _0426_ || _0252_;
  assign _0428_ = _0427_ || _0253_;
  assign _0429_ = _0428_ || _0254_;
  assign _0430_ = _0429_ || _0301_;
  assign _0431_ = _0430_ || _0302_;
  assign _0432_ = _0431_ || _0303_;
  assign _0433_ = _0432_ || _0304_;
  assign _0434_ = _0433_ || _0305_;
  assign _0435_ = _0434_ || _0306_;
  assign _0436_ = _0435_ || _0307_;
  assign _0437_ = _0436_ || _0308_;
  assign _0438_ = ~ _0437_;
  assign \u0.u_div.div_complete_w  = _0459_ & \u0.u_div.div_busy_q ;
  assign _0448_ = \u0.u_csr.opcode_opcode_i  & 32'hfe00707f;
  assign \u0.u_div.div_start_w  = \u0.u_div.opcode_valid_i  & \u0.u_div.div_rem_inst_w ;
  assign _0449_ = _0448_ == 26'h2004033;
  assign _0450_ = _0448_ == 26'h2006033;
  assign _0451_ = _0448_ == 26'h2005033;
  assign _0452_ = _0448_ == 26'h2007033;
  assign _0453_ = \u0.u_div.divisor_q  <= \u0.u_div.dividend_q ;
  assign _0454_ = \u0.u_div.signed_operation_w  && \u0.u_csr.opcode_ra_operand_i [31];
  assign _0455_ = \u0.u_div.signed_operation_w  && \u0.u_div.opcode_rb_operand_i [31];
  assign _0456_ = _0449_ && _0462_;
  assign _0457_ = _0456_ && _0490_;
  assign _0458_ = _0450_ && \u0.u_csr.opcode_ra_operand_i [31];
  assign _0459_ = ! _0489_;
  assign _0460_ = _0457_ || _0458_;
  assign \u0.u_div.div_operation_w  = _0449_ || _0451_;
  assign _0461_ = \u0.u_div.div_operation_w  || _0450_;
  assign \u0.u_div.div_rem_inst_w  = _0461_ || _0452_;
  assign \u0.u_div.signed_operation_w  = _0449_ || _0450_;
  assign _0462_ = \u0.u_csr.opcode_ra_operand_i [31] != \u0.u_div.opcode_rb_operand_i [31];
  assign _0463_ = - \u0.u_csr.opcode_ra_operand_i ;
  assign _0464_ = - \u0.u_div.opcode_rb_operand_i ;
  assign _0465_ = - \u0.u_div.quotient_q ;
  assign _0466_ = - \u0.u_div.dividend_q ;
  assign _0467_ = \u0.u_div.quotient_q  | \u0.u_div.q_mask_q ;
  always @(posedge clk_i)
    \u0.u_div.wb_result_q  <= _0447_;
  always @(posedge clk_i)
    \u0.u_div.valid_q  <= _0446_;
  always @(posedge clk_i)
    \u0.u_div.dividend_q  <= _0441_;
  always @(posedge clk_i)
    \u0.u_div.divisor_q  <= _0442_;
  always @(posedge clk_i)
    \u0.u_div.quotient_q  <= _0445_;
  always @(posedge clk_i)
    \u0.u_div.q_mask_q  <= _0444_;
  always @(posedge clk_i)
    \u0.u_div.div_inst_q  <= _0440_;
  always @(posedge clk_i)
    \u0.u_div.div_busy_q  <= _0439_;
  always @(posedge clk_i)
    \u0.u_div.invert_res_q  <= _0443_;
  assign _0468_ = \u0.u_div.div_complete_w  ? \u0.u_div.div_result_r  : \u0.u_div.wb_result_q ;
  assign _0447_ = rst_i ? 32'h00000000 : _0468_;
  assign _0446_ = rst_i ? 1'h0 : \u0.u_div.div_complete_w ;
  assign \u0.u_div.div_result_r  = \u0.u_div.div_inst_q  ? _0492_ : _0493_;
  assign _0469_ = \u0.u_div.div_start_w  ? _0460_ : \u0.u_div.invert_res_q ;
  assign _0443_ = rst_i ? 1'h0 : _0469_;
  assign _0470_ = \u0.u_div.div_complete_w  ? 1'h0 : \u0.u_div.div_busy_q ;
  assign _0471_ = \u0.u_div.div_start_w  ? 1'h1 : _0470_;
  assign _0439_ = rst_i ? 1'h0 : _0471_;
  assign _0472_ = \u0.u_div.div_start_w  ? \u0.u_div.div_operation_w  : \u0.u_div.div_inst_q ;
  assign _0440_ = rst_i ? 1'h0 : _0472_;
  assign _0473_ = \u0.u_div.div_busy_q  ? { 1'h0, \u0.u_div.q_mask_q [31:1] } : \u0.u_div.q_mask_q ;
  assign _0474_ = \u0.u_div.div_complete_w  ? \u0.u_div.q_mask_q  : _0473_;
  assign _0475_ = \u0.u_div.div_start_w  ? 32'h80000000 : _0474_;
  assign _0444_ = rst_i ? 32'h00000000 : _0475_;
  assign _0476_ = _0453_ ? _0467_ : \u0.u_div.quotient_q ;
  assign _0477_ = \u0.u_div.div_busy_q  ? _0476_ : \u0.u_div.quotient_q ;
  assign _0478_ = \u0.u_div.div_complete_w  ? \u0.u_div.quotient_q  : _0477_;
  assign _0479_ = \u0.u_div.div_start_w  ? 32'h00000000 : _0478_;
  assign _0445_ = rst_i ? 32'h00000000 : _0479_;
  assign _0480_ = \u0.u_div.div_busy_q  ? { 1'h0, \u0.u_div.divisor_q [62:1] } : \u0.u_div.divisor_q ;
  assign _0481_ = \u0.u_div.div_complete_w  ? \u0.u_div.divisor_q  : _0480_;
  assign _0482_ = _0455_ ? { _0464_, 31'h00000000 } : { \u0.u_div.opcode_rb_operand_i , 31'h00000000 };
  assign _0483_ = \u0.u_div.div_start_w  ? _0482_ : _0481_;
  assign _0442_ = rst_i ? 63'h0000000000000000 : _0483_;
  assign _0484_ = _0453_ ? _0491_ : \u0.u_div.dividend_q ;
  assign _0485_ = \u0.u_div.div_busy_q  ? _0484_ : \u0.u_div.dividend_q ;
  assign _0486_ = \u0.u_div.div_complete_w  ? \u0.u_div.dividend_q  : _0485_;
  assign _0487_ = _0454_ ? _0463_ : \u0.u_csr.opcode_ra_operand_i ;
  assign _0488_ = \u0.u_div.div_start_w  ? _0487_ : _0486_;
  assign _0441_ = rst_i ? 32'h00000000 : _0488_;
  assign _0489_ = | \u0.u_div.q_mask_q ;
  assign _0490_ = | \u0.u_div.opcode_rb_operand_i ;
  assign _0491_ = \u0.u_div.dividend_q  - \u0.u_div.divisor_q [31:0];
  assign _0492_ = \u0.u_div.invert_res_q  ? _0465_ : \u0.u_div.quotient_q ;
  assign _0493_ = \u0.u_div.invert_res_q  ? _0466_ : \u0.u_div.dividend_q ;
  assign _0574_ = \u0.u_exec.opcode_pc_i  + { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [7], \u0.u_csr.opcode_opcode_i [30:25], \u0.u_csr.opcode_opcode_i [11:8], 1'h0 };
  assign _0575_ = \u0.u_exec.opcode_pc_i  + { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [19:12], \u0.u_csr.opcode_opcode_i [20], \u0.u_csr.opcode_opcode_i [30:21], 1'h0 };
  assign _0576_ = \u0.u_csr.opcode_ra_operand_i  + { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] };
  assign _0577_ = \u0.u_csr.opcode_opcode_i  & 32'hfe00707f;
  assign _0578_ = \u0.u_csr.opcode_opcode_i  & 15'h707f;
  assign _0579_ = \u0.u_csr.opcode_opcode_i  & 32'hfc00707f;
  assign _0580_ = \u0.u_csr.opcode_opcode_i  & 7'h7f;
  assign _0581_ = _0577_ == 6'h33;
  assign _0582_ = _0577_ == 15'h7033;
  assign _0583_ = _0577_ == 15'h6033;
  assign _0584_ = _0577_ == 13'h1033;
  assign _0585_ = _0577_ == 31'h40005033;
  assign _0586_ = _0577_ == 15'h5033;
  assign _0587_ = _0577_ == 31'h40000033;
  assign _0588_ = _0577_ == 15'h4033;
  assign _0589_ = _0577_ == 14'h2033;
  assign _0590_ = _0577_ == 14'h3033;
  assign _0591_ = _0578_ == 5'h13;
  assign _0592_ = _0578_ == 15'h7013;
  assign _0593_ = _0578_ == 14'h2013;
  assign _0594_ = _0578_ == 14'h3013;
  assign _0595_ = _0578_ == 15'h6013;
  assign _0596_ = _0578_ == 15'h4013;
  assign _0597_ = _0579_ == 13'h1013;
  assign _0598_ = _0579_ == 15'h5013;
  assign _0599_ = _0579_ == 31'h40005013;
  assign _0600_ = _0580_ == 6'h37;
  assign _0601_ = _0580_ == 5'h17;
  assign _0602_ = _0580_ == 7'h6f;
  assign _0603_ = _0578_ == 7'h67;
  assign _0604_ = _0578_ == 7'h63;
  assign _0605_ = \u0.u_csr.opcode_ra_operand_i  == \u0.u_div.opcode_rb_operand_i ;
  assign _0606_ = _0578_ == 13'h1063;
  assign _0607_ = _0578_ == 15'h4063;
  assign _0608_ = _0578_ == 15'h5063;
  assign _0609_ = _0578_ == 15'h6063;
  assign _0610_ = _0578_ == 15'h7063;
  assign _0611_ = \u0.u_csr.opcode_ra_operand_i  >= \u0.u_div.opcode_rb_operand_i ;
  assign _0612_ = \u0.u_exec.branch_r  && \u0.u_div.opcode_valid_i ;
  assign \u0.u_exec.branch_d_request_o  = _0612_ && \u0.u_exec.branch_taken_r ;
  assign _0613_ = _0602_ || _0603_;
  assign _0614_ = \u0.u_csr.opcode_ra_operand_i  < \u0.u_div.opcode_rb_operand_i ;
  assign _0615_ = \u0.u_csr.opcode_ra_operand_i [31] != \u0.u_div.opcode_rb_operand_i [31];
  assign _0616_ = \u0.u_csr.opcode_ra_operand_i  != \u0.u_div.opcode_rb_operand_i ;
  assign _0617_ = _0565_ | _0605_;
  always @(posedge clk_i)
    \u0.u_exec.result_q  <= _0494_;
  assign _0570_ = _0610_ ? _0611_ : 1'h0;
  assign _0569_ = _0610_ ? 1'h1 : 1'h0;
  assign _0564_ = _0609_ ? _0614_ : _0570_;
  assign _0563_ = _0609_ ? 1'h1 : _0569_;
  assign _0618_ = _0615_ ? \u0.u_div.opcode_rb_operand_i [31] : _0626_[31];
  assign _0619_ = _0608_ ? _0618_ : 1'hx;
  assign _0620_ = _0607_ ? 1'hx : _0619_;
  assign _0621_ = _0606_ ? 1'hx : _0620_;
  assign _0622_ = _0604_ ? 1'hx : _0621_;
  assign _0623_ = _0603_ ? 1'hx : _0622_;
  assign _0565_ = _0602_ ? 1'hx : _0623_;
  assign _0558_ = _0608_ ? _0617_ : _0564_;
  assign _0557_ = _0608_ ? 1'h1 : _0563_;
  assign _0559_ = _0615_ ? \u0.u_csr.opcode_ra_operand_i [31] : _0625_[31];
  assign _0553_ = _0607_ ? _0559_ : _0558_;
  assign _0552_ = _0607_ ? 1'h1 : _0557_;
  assign _0548_ = _0606_ ? _0616_ : _0553_;
  assign _0547_ = _0606_ ? 1'h1 : _0552_;
  assign _0543_ = _0604_ ? _0605_ : _0548_;
  assign _0542_ = _0604_ ? 1'h1 : _0547_;
  assign _0538_[31:1] = _0603_ ? _0576_[31:1] : _0574_[31:1];
  assign _0538_[0] = _0603_ ? 1'h0 : _0574_[0];
  assign _0537_ = _0603_ ? 1'h1 : _0543_;
  assign _0536_ = _0603_ ? 1'h1 : _0542_;
  assign \u0.u_exec.branch_target_r  = _0602_ ? _0575_ : _0538_;
  assign \u0.u_exec.branch_taken_r  = _0602_ ? 1'h1 : _0537_;
  assign \u0.u_exec.branch_r  = _0602_ ? 1'h1 : _0536_;
  assign _0624_ = \u0.u_exec.hold_i  ? \u0.u_exec.result_q  : \u0.u_exec.alu_p_w ;
  assign _0494_ = rst_i ? 32'h00000000 : _0624_;
  assign _0531_ = _0613_ ? 3'h4 : 3'h0;
  assign _0532_ = _0613_ ? \u0.u_exec.opcode_pc_i  : 32'h00000000;
  assign _0530_ = _0601_ ? { \u0.u_csr.opcode_opcode_i [31:12], 12'h000 } : { 29'h00000000, _0531_ };
  assign _0529_ = _0601_ ? \u0.u_exec.opcode_pc_i  : _0532_;
  assign _0528_ = _0601_ ? 3'h4 : _0531_;
  assign _0526_ = _0600_ ? { \u0.u_csr.opcode_opcode_i [31:12], 12'h000 } : _0529_;
  assign _0527_ = _0600_ ? 32'h00000000 : _0530_;
  assign _0525_ = _0600_ ? 3'h0 : _0528_;
  assign _0524_ = _0599_ ? { 27'h0000000, \u0.u_csr.opcode_opcode_i [24:20] } : _0527_;
  assign _0523_ = _0599_ ? \u0.u_csr.opcode_ra_operand_i  : _0526_;
  assign _0522_ = _0599_ ? 3'h3 : _0525_;
  assign _0521_ = _0598_ ? { 27'h0000000, \u0.u_csr.opcode_opcode_i [24:20] } : _0524_;
  assign _0520_ = _0598_ ? \u0.u_csr.opcode_ra_operand_i  : _0523_;
  assign _0519_ = _0598_ ? 3'h2 : _0522_;
  assign _0518_ = _0597_ ? { 27'h0000000, \u0.u_csr.opcode_opcode_i [24:20] } : _0521_;
  assign _0517_ = _0597_ ? \u0.u_csr.opcode_ra_operand_i  : _0520_;
  assign _0516_ = _0597_ ? 3'h1 : _0519_;
  assign _0515_ = _0596_ ? { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] } : _0518_;
  assign _0514_ = _0596_ ? \u0.u_csr.opcode_ra_operand_i  : _0517_;
  assign _0513_ = _0596_ ? 4'h9 : { 1'h0, _0516_ };
  assign _0512_ = _0595_ ? { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] } : _0515_;
  assign _0511_ = _0595_ ? \u0.u_csr.opcode_ra_operand_i  : _0514_;
  assign _0510_ = _0595_ ? 4'h8 : _0513_;
  assign _0509_ = _0594_ ? { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] } : _0512_;
  assign _0508_ = _0594_ ? \u0.u_csr.opcode_ra_operand_i  : _0511_;
  assign _0507_ = _0594_ ? 4'ha : _0510_;
  assign _0506_ = _0593_ ? { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] } : _0509_;
  assign _0505_ = _0593_ ? \u0.u_csr.opcode_ra_operand_i  : _0508_;
  assign _0504_ = _0593_ ? 4'hb : _0507_;
  assign _0503_ = _0592_ ? { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] } : _0506_;
  assign _0502_ = _0592_ ? \u0.u_csr.opcode_ra_operand_i  : _0505_;
  assign _0501_ = _0592_ ? 4'h7 : _0504_;
  assign _0500_ = _0591_ ? { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] } : _0503_;
  assign _0499_ = _0591_ ? \u0.u_csr.opcode_ra_operand_i  : _0502_;
  assign _0498_ = _0591_ ? 4'h4 : _0501_;
  assign _0497_ = _0590_ ? \u0.u_div.opcode_rb_operand_i  : _0500_;
  assign _0496_ = _0590_ ? \u0.u_csr.opcode_ra_operand_i  : _0499_;
  assign _0495_ = _0590_ ? 4'ha : _0498_;
  assign _0573_ = _0589_ ? \u0.u_div.opcode_rb_operand_i  : _0497_;
  assign _0572_ = _0589_ ? \u0.u_csr.opcode_ra_operand_i  : _0496_;
  assign _0571_ = _0589_ ? 4'hb : _0495_;
  assign _0568_ = _0588_ ? \u0.u_div.opcode_rb_operand_i  : _0573_;
  assign _0567_ = _0588_ ? \u0.u_csr.opcode_ra_operand_i  : _0572_;
  assign _0566_ = _0588_ ? 4'h9 : _0571_;
  assign _0562_ = _0587_ ? \u0.u_div.opcode_rb_operand_i  : _0568_;
  assign _0561_ = _0587_ ? \u0.u_csr.opcode_ra_operand_i  : _0567_;
  assign _0560_ = _0587_ ? 4'h6 : _0566_;
  assign _0556_ = _0586_ ? \u0.u_div.opcode_rb_operand_i  : _0562_;
  assign _0555_ = _0586_ ? \u0.u_csr.opcode_ra_operand_i  : _0561_;
  assign _0554_ = _0586_ ? 4'h2 : _0560_;
  assign _0551_ = _0585_ ? \u0.u_div.opcode_rb_operand_i  : _0556_;
  assign _0550_ = _0585_ ? \u0.u_csr.opcode_ra_operand_i  : _0555_;
  assign _0549_ = _0585_ ? 4'h3 : _0554_;
  assign _0546_ = _0584_ ? \u0.u_div.opcode_rb_operand_i  : _0551_;
  assign _0545_ = _0584_ ? \u0.u_csr.opcode_ra_operand_i  : _0550_;
  assign _0544_ = _0584_ ? 4'h1 : _0549_;
  assign _0541_ = _0583_ ? \u0.u_div.opcode_rb_operand_i  : _0546_;
  assign _0540_ = _0583_ ? \u0.u_csr.opcode_ra_operand_i  : _0545_;
  assign _0539_ = _0583_ ? 4'h8 : _0544_;
  assign _0535_ = _0582_ ? \u0.u_div.opcode_rb_operand_i  : _0541_;
  assign _0534_ = _0582_ ? \u0.u_csr.opcode_ra_operand_i  : _0540_;
  assign _0533_ = _0582_ ? 4'h7 : _0539_;
  assign \u0.u_exec.alu_input_b_r  = _0581_ ? \u0.u_div.opcode_rb_operand_i  : _0535_;
  assign \u0.u_exec.alu_input_a_r  = _0581_ ? \u0.u_csr.opcode_ra_operand_i  : _0534_;
  assign \u0.u_exec.alu_func_r  = _0581_ ? 4'h4 : _0533_;
  assign _0625_ = \u0.u_csr.opcode_ra_operand_i  - \u0.u_div.opcode_rb_operand_i ;
  assign _0626_ = \u0.u_div.opcode_rb_operand_i  - \u0.u_csr.opcode_ra_operand_i ;
  assign _0639_ = \u0.u_exec.alu_input_a_r  + \u0.u_exec.alu_input_b_r ;
  assign _0640_ = \u0.u_exec.alu_input_a_r  & \u0.u_exec.alu_input_b_r ;
  assign _0642_ = \u0.u_exec.alu_func_r  == 2'h3;
  assign _0643_ = \u0.u_exec.alu_input_a_r [31] && _0642_;
  assign _0644_ = \u0.u_exec.alu_input_a_r  < \u0.u_exec.alu_input_b_r ;
  assign _0645_ = \u0.u_exec.alu_input_a_r [31] != \u0.u_exec.alu_input_b_r [31];
  assign _0646_ = \u0.u_exec.alu_input_a_r  | \u0.u_exec.alu_input_b_r ;
  assign _0638_ = _0645_ ? _0657_[0] : _0658_[0];
  assign _0647_ = \u0.u_exec.alu_func_r  == 4'hb;
  assign _0637_ = \u0.u_exec.alu_input_b_r [4] ? { _0636_, _0635_[31:16] } : _0635_;
  assign _0648_[0] = \u0.u_exec.alu_func_r  == 2'h2;
  assign _0635_ = \u0.u_exec.alu_input_b_r [3] ? { _0636_[15:8], _0634_[31:8] } : _0634_;
  assign _0634_ = \u0.u_exec.alu_input_b_r [2] ? { _0636_[15:12], _0633_[31:4] } : _0633_;
  assign _0649_ = | { _0648_[0], _0642_ };
  assign _0633_ = \u0.u_exec.alu_input_b_r [1] ? { _0636_[15:14], _0632_[31:2] } : _0632_;
  assign _0632_ = \u0.u_exec.alu_input_b_r [0] ? { _0636_[15], \u0.u_exec.alu_input_a_r [31:1] } : \u0.u_exec.alu_input_a_r ;
  assign _0636_ = _0643_ ? 16'hffff : 16'h0000;
  assign _0627_ = \u0.u_exec.alu_input_b_r [4] ? { _0631_[15:0], 16'h0000 } : _0631_;
  assign _0650_ = \u0.u_exec.alu_func_r  == 1'h1;
  assign _0631_ = \u0.u_exec.alu_input_b_r [3] ? { _0630_[23:0], 8'h00 } : _0630_;
  assign _0630_ = \u0.u_exec.alu_input_b_r [2] ? { _0629_[27:0], 4'h0 } : _0629_;
  assign _0629_ = \u0.u_exec.alu_input_b_r [1] ? { _0628_[29:0], 2'h0 } : _0628_;
  assign _0628_ = \u0.u_exec.alu_input_b_r [0] ? { \u0.u_exec.alu_input_a_r [30:0], 1'h0 } : \u0.u_exec.alu_input_a_r ;
  function [31:0] _2044_;
    input [31:0] a;
    input [287:0] b;
    input [8:0] s;
    casez (s) // synopsys parallel_case
      9'b????????1:
        _2044_ = b[31:0];
      9'b???????1?:
        _2044_ = b[63:32];
      9'b??????1??:
        _2044_ = b[95:64];
      9'b?????1???:
        _2044_ = b[127:96];
      9'b????1????:
        _2044_ = b[159:128];
      9'b???1?????:
        _2044_ = b[191:160];
      9'b??1??????:
        _2044_ = b[223:192];
      9'b?1???????:
        _2044_ = b[255:224];
      9'b1????????:
        _2044_ = b[287:256];
      default:
        _2044_ = a;
    endcase
  endfunction
  assign \u0.u_exec.alu_p_w  = _2044_(\u0.u_exec.alu_input_a_r , { _0627_, _0637_, _0639_, \u0.u_exec.u_alu.sub_res_w , _0640_, _0646_, _0659_, 31'h00000000, _0641_[0], 31'h00000000, _0638_ }, { _0650_, _0649_, _0656_, _0655_, _0654_, _0653_, _0652_, _0651_, _0647_ });
  assign _0651_ = \u0.u_exec.alu_func_r  == 4'ha;
  assign _0652_ = \u0.u_exec.alu_func_r  == 4'h9;
  assign _0653_ = \u0.u_exec.alu_func_r  == 4'h8;
  assign _0654_ = \u0.u_exec.alu_func_r  == 3'h7;
  assign _0655_ = \u0.u_exec.alu_func_r  == 3'h6;
  assign _0656_ = \u0.u_exec.alu_func_r  == 3'h4;
  assign \u0.u_exec.u_alu.sub_res_w  = \u0.u_exec.alu_input_a_r  - \u0.u_exec.alu_input_b_r ;
  assign _0641_[0] = _0644_ ? 1'h1 : 1'h0;
  assign _0657_[0] = \u0.u_exec.alu_input_a_r [31] ? 1'h1 : 1'h0;
  assign _0658_[0] = \u0.u_exec.u_alu.sub_res_w [31] ? 1'h1 : 1'h0;
  assign _0659_ = \u0.u_exec.alu_input_a_r  ^ \u0.u_exec.alu_input_b_r ;
  assign _0669_ = { \u0.u_fetch.pc_f_q [31:2], 2'h0 } + 3'h4;
  assign _0670_ = \u0.u_fetch.active_q  & \u0.u_fetch.fetch_accept_i ;
  assign \fifo_i_rd.in  = _0670_ & _0676_;
  assign \u0.u_decode.genblk1.u_dec.valid_i  = _0680_ & _0678_;
  assign _0671_ = \fifo_i_rd.in  && mem_i_accept_i;
  assign _0672_ = \u0.u_fetch.branch_q  && _0681_;
  assign \u0.u_fetch.icache_busy_w  = \u0.u_fetch.icache_fetch_q  && _0677_;
  assign _0673_ = \u0.u_decode.genblk1.u_dec.valid_i  && _0674_;
  assign _0674_ = ! \u0.u_fetch.fetch_accept_i ;
  assign _0675_ = ! mem_i_accept_i;
  assign _0676_ = ! \u0.u_fetch.icache_busy_w ;
  assign _0677_ = ! mem_i_valid_i;
  assign _0678_ = ! \u0.u_fetch.fetch_resp_drop_w ;
  assign _0679_ = _0674_ || \u0.u_fetch.icache_busy_w ;
  assign \u0.u_fetch.stall_w  = _0679_ || _0675_;
  assign _0680_ = mem_i_valid_i || \u0.u_fetch.skid_valid_q ;
  assign _0681_ = ~ \u0.u_fetch.stall_w ;
  assign \u0.u_fetch.fetch_resp_drop_w  = \u0.u_fetch.branch_q  | \u0.u_fetch.branch_d_q ;
  always @(posedge clk_i)
    \u0.u_fetch.skid_buffer_q  <= _0667_;
  always @(posedge clk_i)
    \u0.u_fetch.skid_valid_q  <= _0668_;
  always @(posedge clk_i)
    \u0.u_fetch.pc_d_q  <= _0665_;
  always @(posedge clk_i)
    \u0.u_fetch.branch_d_q  <= _0661_;
  always @(posedge clk_i)
    \u0.u_fetch.pc_f_q  <= _0666_;
  always @(posedge clk_i)
    \u0.u_fetch.icache_fetch_q  <= _0664_;
  always @(posedge clk_i)
    \u0.u_fetch.active_q  <= _0660_;
  always @(posedge clk_i)
    \u0.u_fetch.branch_q  <= _0663_;
  always @(posedge clk_i)
    \u0.u_fetch.branch_pc_q  <= _0662_;
  assign _0682_ = _0673_ ? 1'h1 : 1'h0;
  assign _0668_ = rst_i ? 1'h0 : _0682_;
  assign _0683_ = _0673_ ? { \u0.u_decode.fetch_in_fault_page_i , \u0.u_decode.fetch_in_fault_fetch_i , \u0.u_exec.opcode_pc_i , \u0.u_decode.fetch_in_instr_i  } : 66'h00000000000000000;
  assign _0667_ = rst_i ? 66'h00000000000000000 : _0683_;
  assign _0684_ = _0671_ ? \u0.u_fetch.pc_f_q  : \u0.u_fetch.pc_d_q ;
  assign _0665_ = rst_i ? 32'h00000000 : _0684_;
  assign _0685_ = \u0.u_fetch.stall_w  ? \u0.u_fetch.branch_d_q  : 1'h0;
  assign _0686_ = _0672_ ? 1'h1 : _0685_;
  assign _0661_ = rst_i ? 1'h0 : _0686_;
  assign _0687_ = \u0.u_fetch.stall_w  ? \u0.u_fetch.pc_f_q  : _0669_;
  assign _0688_ = _0672_ ? \u0.u_fetch.branch_pc_q  : _0687_;
  assign _0666_ = rst_i ? 32'h00000000 : _0688_;
  assign _0689_ = mem_i_valid_i ? 1'h0 : \u0.u_fetch.icache_fetch_q ;
  assign _0690_ = _0671_ ? 1'h1 : _0689_;
  assign _0664_ = rst_i ? 1'h0 : _0690_;
  assign _0691_ = _0672_ ? 1'h1 : \u0.u_fetch.active_q ;
  assign _0660_ = rst_i ? 1'h0 : _0691_;
  assign _0692_ = _0671_ ? 32'h00000000 : \u0.u_fetch.branch_pc_q ;
  assign _0693_ = \u0.u_fetch.branch_request_i  ? \u0.u_fetch.branch_pc_i  : _0692_;
  assign _0662_ = rst_i ? 32'h00000000 : _0693_;
  assign _0694_ = _0671_ ? 1'h0 : \u0.u_fetch.branch_q ;
  assign _0695_ = \u0.u_fetch.branch_request_i  ? 1'h1 : _0694_;
  assign _0663_ = rst_i ? 1'h0 : _0695_;
  assign \u0.u_exec.opcode_pc_i  = \u0.u_fetch.skid_valid_q  ? \u0.u_fetch.skid_buffer_q [63:32] : { \u0.u_fetch.pc_d_q [31:2], 2'h0 };
  assign \u0.u_decode.fetch_in_instr_i  = \u0.u_fetch.skid_valid_q  ? \u0.u_fetch.skid_buffer_q [31:0] : mem_i_inst_i;
  assign \u0.u_decode.fetch_in_fault_fetch_i  = \u0.u_fetch.skid_valid_q  ? \u0.u_fetch.skid_buffer_q [64] : mem_i_error_i;
  assign \u0.u_decode.fetch_in_fault_page_i  = \u0.u_fetch.skid_valid_q  ? \u0.u_fetch.skid_buffer_q [65] : 1'h0;
  assign _0707_ = 1'h0 & _0732_;
  assign _0708_ = \u0.u_decode.genblk1.u_dec.valid_i  & _0733_;
  assign \u0.u_issue.opcode_valid_w  = _0708_ & _0734_;
  assign \u0.u_csr.opcode_valid_i  = \u0.u_div.opcode_valid_i  & _0735_;
  assign _0710_ = \u0.u_issue.pipe_rd_wb_w  == \u0.u_csr.opcode_opcode_i [19:15];
  assign _0711_ = \u0.u_issue.pipe_rd_wb_w  == \u0.u_csr.opcode_opcode_i [24:20];
  assign _0712_ = \u0.u_issue.pipe_rd_e2_w  == \u0.u_csr.opcode_opcode_i [19:15];
  assign _0713_ = \u0.u_issue.pipe_rd_e2_w  == \u0.u_csr.opcode_opcode_i [24:20];
  assign _0714_ = \u0.u_issue.pipe_rd_e1_w  == \u0.u_csr.opcode_opcode_i [19:15];
  assign _0715_ = \u0.u_issue.pipe_rd_e1_w  == \u0.u_csr.opcode_opcode_i [24:20];
  assign _0716_ = ! \u0.u_csr.opcode_opcode_i [19:15];
  assign _0717_ = ! \u0.u_csr.opcode_opcode_i [24:20];
  assign _0718_ = \u0.u_div.opcode_valid_i  && \u0.u_decode.genblk1.u_dec.div_o ;
  assign _0719_ = \u0.u_csr.opcode_valid_i  && \u0.u_decode.genblk1.u_dec.csr_o ;
  assign _0720_ = _0724_ && _0726_;
  assign _0721_ = \u0.u_issue.opcode_valid_w  && _0722_;
  assign \u0.u_csr.opcode_invalid_i  = \u0.u_div.opcode_valid_i  && \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign _0722_ = ! _0731_;
  assign _0723_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [1] || \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [5];
  assign _0724_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [1] || \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [2];
  assign _0725_ = \u0.u_decode.genblk1.u_dec.mul_o  || \u0.u_decode.genblk1.u_dec.div_o ;
  assign _0726_ = _0725_ || \u0.u_decode.genblk1.u_dec.csr_o ;
  assign _0727_ = \u0.u_issue.lsu_stall_i  || \u0.u_exec.hold_i ;
  assign _0728_ = _0727_ || \u0.u_issue.div_pending_q ;
  assign _0729_ = _0728_ || \u0.u_issue.csr_pending_q ;
  assign _0730_ = _0743_ || _0744_;
  assign _0731_ = _0730_ || _0745_;
  assign \u0.u_csr.interrupt_inhibit_i  = \u0.u_issue.csr_pending_q  || \u0.u_decode.genblk1.u_dec.csr_o ;
  assign _0732_ = ~ _0746_;
  assign _0733_ = ~ \u0.u_issue.pipe_squash_e1_e2_w ;
  assign _0734_ = ~ \u0.u_csr.branch_q ;
  assign _0735_ = ~ \u0.u_csr.take_interrupt_q ;
  assign _0736_ = _0707_ | _0746_;
  assign \u0.u_fetch.branch_request_i  = \u0.u_csr.branch_q  | \u0.u_exec.branch_d_request_o ;
  always @(posedge clk_i)
    \u0.u_issue.csr_pending_q  <= _0696_;
  always @(posedge clk_i)
    \u0.u_issue.div_pending_q  <= _0697_;
  assign \u0.u_div.opcode_rb_operand_i  = _0717_ ? 32'h00000000 : _0706_;
  assign \u0.u_csr.opcode_ra_operand_i  = _0716_ ? 32'h00000000 : _0705_;
  assign _0706_ = _0715_ ? \u0.u_exec.result_q  : _0702_;
  assign _0705_ = _0714_ ? \u0.u_exec.result_q  : _0701_;
  assign _0702_ = _0713_ ? \u0.u_issue.pipe_result_e2_w  : _0699_;
  assign _0701_ = _0712_ ? \u0.u_issue.pipe_result_e2_w  : _0698_;
  assign _0699_ = _0711_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.issue_rb_value_w ;
  assign _0698_ = _0710_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.issue_ra_value_w ;
  assign _0703_ = _0721_ ? 1'h1 : 1'h0;
  assign \u0.u_div.opcode_valid_i  = _0729_ ? 1'h0 : _0703_;
  assign _0704_ = _0720_ ? 32'hffffffff : _0700_;
  assign _0700_ = _0723_ ? _0736_ : 32'h00000000;
  assign _0737_ = \u0.u_issue.pipe_csr_wb_w  ? 1'h0 : \u0.u_issue.csr_pending_q ;
  assign _0738_ = _0719_ ? 1'h1 : _0737_;
  assign _0739_ = \u0.u_issue.pipe_squash_e1_e2_w  ? 1'h0 : _0738_;
  assign _0696_ = rst_i ? 1'h0 : _0739_;
  assign _0740_ = \u0.u_div.valid_q  ? 1'h0 : \u0.u_issue.div_pending_q ;
  assign _0741_ = _0718_ ? 1'h1 : _0740_;
  assign _0742_ = \u0.u_issue.pipe_squash_e1_e2_w  ? 1'h0 : _0741_;
  assign _0697_ = rst_i ? 1'h0 : _0742_;
  wire [31:0] _2828_ = _0704_;
  assign _0743_ = _2828_[\u0.u_csr.opcode_opcode_i [19:15] +: 1];
  wire [31:0] _2829_ = _0704_;
  assign _0744_ = _2829_[\u0.u_csr.opcode_opcode_i [24:20] +: 1];
  wire [31:0] _2830_ = _0704_;
  assign _0745_ = _2830_[\u0.u_csr.opcode_opcode_i [11:7] +: 1];
  assign _0746_ = 1'h1 << \u0.u_issue.pipe_rd_e1_w ;
  assign \u0.u_fetch.branch_pc_i  = \u0.u_csr.branch_q  ? \u0.u_csr.branch_target_q  : \u0.u_exec.branch_target_r ;
  assign \u0.u_issue.issue_fault_w  = \u0.u_decode.fetch_in_fault_fetch_i  ? 5'h11 : _0709_[4:0];
  assign _0709_[4:0] = \u0.u_decode.fetch_in_fault_page_i  ? 5'h1c : 5'h00;
  assign \u0.u_fetch.fetch_accept_i  = \u0.u_issue.opcode_valid_w  ? \u0.u_csr.opcode_valid_i  : 1'h1;
  assign _0770_ = \u0.u_decode.genblk1.u_dec.lsu_o  & \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign _0771_ = _0770_ & _0801_;
  assign _0772_ = \u0.u_decode.genblk1.u_dec.lsu_o  & _0802_;
  assign _0773_ = _0772_ & _0801_;
  assign _0774_ = \u0.u_decode.genblk1.u_dec.csr_o  & _0801_;
  assign _0775_ = \u0.u_decode.genblk1.u_dec.div_o  & _0801_;
  assign _0776_ = \u0.u_decode.genblk1.u_dec.mul_o  & _0801_;
  assign _0777_ = \u0.u_decode.genblk1.u_dec.branch_o  & _0801_;
  assign _0778_ = \u0.u_decode.genblk1.u_dec.rd_valid_o  & _0801_;
  assign \u0.u_issue.pipe_rd_e1_w  = { \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [7], \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [7], \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [7], \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [7], \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [7] } & \u0.u_issue.u_pipe_ctrl.opcode_e1_q [11:7];
  assign \u0.u_issue.u_pipe_ctrl.valid_e2_w  = \u0.u_issue.u_pipe_ctrl.valid_e2_q  & _0803_;
  assign \u0.u_issue.pipe_rd_e2_w  = { _0788_, _0788_, _0788_, _0788_, _0788_ } & \u0.u_issue.u_pipe_ctrl.opcode_e2_q [11:7];
  assign _0779_ = _0810_ & _0806_;
  assign _0780_ = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q  & 10'h37f;
  assign \u0.u_issue.u_pipe_ctrl.valid_wb_o  = \u0.u_issue.u_pipe_ctrl.valid_wb_q  & _0803_;
  assign \u0.u_issue.pipe_csr_wb_w  = \u0.u_issue.u_pipe_ctrl.ctrl_wb_q [3] & _0803_;
  assign \u0.u_issue.pipe_rd_wb_w  = { _0795_, _0795_, _0795_, _0795_, _0795_ } & \u0.u_issue.u_pipe_ctrl.opcode_wb_q [11:7];
  assign \u0.u_issue.u_pipe_ctrl.branch_misaligned_w  = \u0.u_exec.branch_d_request_o  && _0798_;
  assign _0782_ = \u0.u_div.opcode_valid_i  && \u0.u_div.opcode_valid_i ;
  assign _0783_ = _0782_ && _0799_;
  assign _0784_ = $signed(32'h00000001) && \u0.u_issue.u_pipe_ctrl.valid_e2_w ;
  assign _0785_ = _0784_ && _0797_;
  assign _0786_ = _0784_ && \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [5];
  assign _0787_ = \u0.u_issue.u_pipe_ctrl.valid_e2_w  && \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [7];
  assign _0788_ = _0787_ && _0804_;
  assign _0789_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [4] && _0805_;
  assign _0790_ = \u0.u_issue.u_pipe_ctrl.valid_e2_q  && _0797_;
  assign _0791_ = _0790_ && \u0.u_issue.u_pipe_ctrl.mem_complete_i ;
  assign _0792_ = \u0.u_issue.u_pipe_ctrl.valid_e2_w  && _0797_;
  assign _0793_ = \u0.u_issue.u_pipe_ctrl.valid_e2_w  && \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [5];
  assign _0794_ = \u0.u_issue.u_pipe_ctrl.valid_wb_o  && \u0.u_issue.u_pipe_ctrl.ctrl_wb_q [7];
  assign _0795_ = _0794_ && _0804_;
  assign _0796_ = \u0.u_issue.pipe_squash_e1_e2_w  || 1'h0;
  assign _0797_ = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [1] || \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [2];
  assign \u0.u_exec.hold_i  = _0789_ || _0779_;
  assign _0798_ = | \u0.u_exec.branch_target_r [1:0];
  assign _0799_ = ~ _0796_;
  assign _0800_ = ~ _0809_;
  assign _0801_ = ~ \u0.u_csr.take_interrupt_q ;
  assign _0802_ = ~ \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign _0803_ = ~ \u0.u_exec.hold_i ;
  assign _0804_ = ~ \u0.u_exec.hold_i ;
  assign _0805_ = ~ \u0.u_div.valid_q ;
  assign _0806_ = ~ \u0.u_issue.u_pipe_ctrl.mem_complete_i ;
  assign _0807_ = \u0.u_decode.genblk1.u_dec.lsu_o  | \u0.u_decode.genblk1.u_dec.csr_o ;
  assign _0808_ = _0807_ | \u0.u_decode.genblk1.u_dec.div_o ;
  assign _0809_ = _0808_ | \u0.u_decode.genblk1.u_dec.mul_o ;
  assign _0810_ = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [1] | \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [2];
  assign \u0.u_issue.pipe_squash_e1_e2_w  = \u0.u_issue.u_pipe_ctrl.squash_e1_e2_w  | \u0.u_issue.u_pipe_ctrl.squash_e1_e2_q ;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.valid_wb_q  <= _0768_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.ctrl_wb_q  <= _0753_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q  <= _0750_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  <= _0748_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.result_wb_q  <= _0764_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.pc_wb_q  <= _0762_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.opcode_wb_q  <= _0759_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.exception_wb_q  <= _0756_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.squash_e1_e2_q  <= _0765_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.result_e2_q  <= _0763_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.valid_e2_q  <= _0767_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.ctrl_e2_q  <= _0752_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.csr_wr_e2_q  <= _0749_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.csr_wdata_e2_q  <= _0747_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.pc_e2_q  <= _0761_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.opcode_e2_q  <= _0758_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.exception_e2_q  <= _0755_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.exception_e1_q  <= _0754_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.valid_e1_q  <= _0766_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.ctrl_e1_q  <= _0751_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.pc_e1_q  <= _0760_;
  always @(posedge clk_i)
    \u0.u_issue.u_pipe_ctrl.opcode_e1_q  <= _0757_;
  assign _0811_ = 1'h0 ? 6'h00 : \u0.u_issue.u_pipe_ctrl.exception_e2_r ;
  assign _0812_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.exception_wb_q  : _0811_;
  assign _0756_ = rst_i ? 6'h00 : _0812_;
  assign _0813_ = 1'h0 ? 32'h00000000 : \u0.u_issue.u_pipe_ctrl.opcode_e2_q ;
  assign _0814_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.opcode_wb_q  : _0813_;
  assign _0759_ = rst_i ? 32'h00000000 : _0814_;
  assign _0815_ = 1'h0 ? 32'h00000000 : \u0.u_issue.u_pipe_ctrl.pc_e2_q ;
  assign _0816_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.pc_wb_q  : _0815_;
  assign _0762_ = rst_i ? 32'h00000000 : _0816_;
  assign _0817_ = _0793_ ? \u0.u_mul.result_e2_q  : \u0.u_issue.u_pipe_ctrl.result_e2_q ;
  assign _0818_ = _0792_ ? \u0.u_issue.u_pipe_ctrl.mem_result_e2_i  : _0817_;
  assign _0819_ = 1'h0 ? 32'h00000000 : _0818_;
  assign _0820_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : _0819_;
  assign _0764_ = rst_i ? 32'h00000000 : _0820_;
  assign _0821_ = 1'h0 ? 32'h00000000 : \u0.u_issue.u_pipe_ctrl.csr_wdata_e2_q ;
  assign _0822_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q  : _0821_;
  assign _0748_ = rst_i ? 32'h00000000 : _0822_;
  assign _0823_ = 1'h0 ? 1'h0 : \u0.u_issue.u_pipe_ctrl.csr_wr_e2_q ;
  assign _0824_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q  : _0823_;
  assign _0750_ = rst_i ? 1'h0 : _0824_;
  assign _0825_ = \u0.u_issue.u_pipe_ctrl.squash_e1_e2_w  ? _0780_ : \u0.u_issue.u_pipe_ctrl.ctrl_e2_q ;
  assign _0826_ = 1'h0 ? 10'h000 : _0825_;
  assign _0827_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_wb_q  : _0826_;
  assign _0753_ = rst_i ? 10'h000 : _0827_;
  assign _0828_ = _0830_ ? 1'h0 : \u0.u_issue.u_pipe_ctrl.valid_e2_q ;
  assign _0830_ = | _0829_;
  assign _0829_[0] = \u0.u_issue.u_pipe_ctrl.exception_e2_r  == 5'h14;
  assign _0829_[1] = \u0.u_issue.u_pipe_ctrl.exception_e2_r  == 5'h15;
  assign _0829_[2] = \u0.u_issue.u_pipe_ctrl.exception_e2_r  == 5'h16;
  assign _0829_[3] = \u0.u_issue.u_pipe_ctrl.exception_e2_r  == 5'h17;
  assign _0829_[4] = \u0.u_issue.u_pipe_ctrl.exception_e2_r  == 5'h1d;
  assign _0829_[5] = \u0.u_issue.u_pipe_ctrl.exception_e2_r  == 5'h1f;
  assign _0831_ = 1'h0 ? 1'h0 : _0828_;
  assign _0832_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.valid_wb_q  : _0831_;
  assign _0768_ = rst_i ? 1'h0 : _0832_;
  assign _0833_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.squash_e1_e2_q  : \u0.u_issue.u_pipe_ctrl.squash_e1_e2_w ;
  assign _0765_ = rst_i ? 1'h0 : _0833_;
  assign \u0.u_issue.u_pipe_ctrl.exception_e2_r  = _0791_ ? { 1'h0, \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i [4:0] } : \u0.u_issue.u_pipe_ctrl.exception_e2_q ;
  assign _0769_ = _0786_ ? \u0.u_mul.result_e2_q  : \u0.u_issue.u_pipe_ctrl.result_e2_q ;
  assign \u0.u_issue.pipe_result_e2_w  = _0785_ ? \u0.u_issue.u_pipe_ctrl.mem_result_e2_i  : _0769_;
  assign _0834_ = _0835_ ? \u0.u_issue.u_pipe_ctrl.exception_e1_q  : \u0.u_csr.exception_e1_q ;
  assign _0836_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [8] ? 6'h20 : _0834_;
  assign _0837_ = _0796_ ? 6'h00 : _0836_;
  assign _0838_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.exception_e2_q  : _0837_;
  assign _0755_ = rst_i ? 6'h00 : _0838_;
  assign _0839_ = _0796_ ? 32'h00000000 : \u0.u_issue.u_pipe_ctrl.opcode_e1_q ;
  assign _0840_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.opcode_e2_q  : _0839_;
  assign _0758_ = rst_i ? 32'h00000000 : _0840_;
  assign _0841_ = _0796_ ? 32'h00000000 : \u0.u_issue.u_pipe_ctrl.pc_e1_q ;
  assign _0842_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.pc_e2_q  : _0841_;
  assign _0761_ = rst_i ? 32'h00000000 : _0842_;
  assign _0843_ = _0796_ ? 32'h00000000 : \u0.u_csr.csr_wdata_e1_q ;
  assign _0844_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.csr_wdata_e2_q  : _0843_;
  assign _0747_ = rst_i ? 32'h00000000 : _0844_;
  assign _0845_ = _0796_ ? 1'h0 : \u0.u_csr.rd_valid_e1_q ;
  assign _0846_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.csr_wr_e2_q  : _0845_;
  assign _0749_ = rst_i ? 1'h0 : _0846_;
  assign _0847_ = _0796_ ? 10'h000 : \u0.u_issue.u_pipe_ctrl.ctrl_e1_q ;
  assign _0848_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e2_q  : _0847_;
  assign _0752_ = rst_i ? 10'h000 : _0848_;
  assign _0849_ = _0835_ ? 1'h0 : \u0.u_issue.u_pipe_ctrl.valid_e1_q ;
  assign _0850_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [8] ? \u0.u_issue.u_pipe_ctrl.valid_e1_q  : _0849_;
  assign _0851_ = _0796_ ? 1'h0 : _0850_;
  assign _0852_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.valid_e2_q  : _0851_;
  assign _0767_ = rst_i ? 1'h0 : _0852_;
  assign _0853_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [3] ? \u0.u_csr.rd_result_e1_q  : \u0.u_exec.result_q ;
  assign _0854_ = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [4] ? \u0.u_div.wb_result_q  : _0853_;
  assign _0855_ = _0796_ ? 32'h00000000 : _0854_;
  assign _0856_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.result_e2_q  : _0855_;
  assign _0763_ = rst_i ? 32'h00000000 : _0856_;
  assign _0857_ = _0783_ ? 1'h1 : 1'h0;
  assign _0858_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [9] : _0857_;
  assign _0751_[9] = rst_i ? 1'h0 : _0858_;
  assign _0859_ = _0783_ ? _0778_ : 1'h0;
  assign _0860_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [7] : _0859_;
  assign _0751_[7] = rst_i ? 1'h0 : _0860_;
  assign _0861_ = _0783_ ? _0777_ : 1'h0;
  assign _0862_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [6] : _0861_;
  assign _0751_[6] = rst_i ? 1'h0 : _0862_;
  assign _0863_ = _0783_ ? _0776_ : 1'h0;
  assign _0864_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [5] : _0863_;
  assign _0751_[5] = rst_i ? 1'h0 : _0864_;
  assign _0865_ = _0783_ ? _0775_ : 1'h0;
  assign _0866_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [4] : _0865_;
  assign _0751_[4] = rst_i ? 1'h0 : _0866_;
  assign _0867_ = _0783_ ? _0774_ : 1'h0;
  assign _0868_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [3] : _0867_;
  assign _0751_[3] = rst_i ? 1'h0 : _0868_;
  assign _0869_ = _0783_ ? _0773_ : 1'h0;
  assign _0870_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [2] : _0869_;
  assign _0751_[2] = rst_i ? 1'h0 : _0870_;
  assign _0871_ = _0783_ ? _0771_ : 1'h0;
  assign _0872_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [1] : _0871_;
  assign _0751_[1] = rst_i ? 1'h0 : _0872_;
  assign _0873_ = _0783_ ? _0800_ : 1'h0;
  assign _0874_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [0] : _0873_;
  assign _0751_[0] = rst_i ? 1'h0 : _0874_;
  assign _0875_ = _0783_ ? \u0.u_csr.take_interrupt_q  : 1'h0;
  assign _0876_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [8] : _0875_;
  assign _0751_[8] = rst_i ? 1'h0 : _0876_;
  assign _0877_ = _0783_ ? \u0.u_csr.opcode_opcode_i  : 32'h00000000;
  assign _0878_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.opcode_e1_q  : _0877_;
  assign _0757_ = rst_i ? 32'h00000000 : _0878_;
  assign _0879_ = _0783_ ? \u0.u_exec.opcode_pc_i  : 32'h00000000;
  assign _0880_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.pc_e1_q  : _0879_;
  assign _0760_ = rst_i ? 32'h00000000 : _0880_;
  assign _0881_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.valid_e1_q  : _0857_;
  assign _0766_ = rst_i ? 1'h0 : _0881_;
  assign _0882_ = _0783_ ? _0885_ : 6'h00;
  assign _0883_ = \u0.u_exec.hold_i  ? \u0.u_issue.u_pipe_ctrl.exception_e1_q  : _0882_;
  assign _0754_ = rst_i ? 6'h00 : _0883_;
  assign _0884_ = | { 1'h0, \u0.u_issue.issue_fault_w  };
  assign _0835_ = | \u0.u_issue.u_pipe_ctrl.exception_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.squash_e1_e2_w  = | \u0.u_issue.u_pipe_ctrl.exception_e2_r ;
  assign _0885_ = _0884_ ? { 1'h0, \u0.u_issue.issue_fault_w  } : { 1'h0, _0781_[4:0] };
  assign _0781_[4:0] = \u0.u_issue.u_pipe_ctrl.branch_misaligned_w  ? 5'h10 : 5'h00;
  assign _0917_ = \u0.u_issue.pipe_rd_wb_w  == 1'h1;
  assign _0918_ = \u0.u_issue.pipe_rd_wb_w  == 2'h2;
  assign _0919_ = \u0.u_issue.pipe_rd_wb_w  == 2'h3;
  assign _0920_ = \u0.u_issue.pipe_rd_wb_w  == 3'h4;
  assign _0921_ = \u0.u_issue.pipe_rd_wb_w  == 3'h5;
  assign _0922_ = \u0.u_issue.pipe_rd_wb_w  == 3'h6;
  assign _0923_ = \u0.u_issue.pipe_rd_wb_w  == 3'h7;
  assign _0924_ = \u0.u_issue.pipe_rd_wb_w  == 4'h8;
  assign _0925_ = \u0.u_issue.pipe_rd_wb_w  == 4'h9;
  assign _0926_ = \u0.u_issue.pipe_rd_wb_w  == 4'ha;
  assign _0927_ = \u0.u_issue.pipe_rd_wb_w  == 4'hb;
  assign _0928_ = \u0.u_issue.pipe_rd_wb_w  == 4'hc;
  assign _0929_ = \u0.u_issue.pipe_rd_wb_w  == 4'hd;
  assign _0930_ = \u0.u_issue.pipe_rd_wb_w  == 4'he;
  assign _0931_ = \u0.u_issue.pipe_rd_wb_w  == 4'hf;
  assign _0932_ = \u0.u_issue.pipe_rd_wb_w  == 5'h10;
  assign _0933_ = \u0.u_issue.pipe_rd_wb_w  == 5'h11;
  assign _0934_ = \u0.u_issue.pipe_rd_wb_w  == 5'h12;
  assign _0935_ = \u0.u_issue.pipe_rd_wb_w  == 5'h13;
  assign _0936_ = \u0.u_issue.pipe_rd_wb_w  == 5'h14;
  assign _0937_ = \u0.u_issue.pipe_rd_wb_w  == 5'h15;
  assign _0938_ = \u0.u_issue.pipe_rd_wb_w  == 5'h16;
  assign _0939_ = \u0.u_issue.pipe_rd_wb_w  == 5'h17;
  assign _0940_ = \u0.u_issue.pipe_rd_wb_w  == 5'h18;
  assign _0941_ = \u0.u_issue.pipe_rd_wb_w  == 5'h19;
  assign _0942_ = \u0.u_issue.pipe_rd_wb_w  == 5'h1a;
  assign _0943_ = \u0.u_issue.pipe_rd_wb_w  == 5'h1b;
  assign _0944_ = \u0.u_issue.pipe_rd_wb_w  == 5'h1c;
  assign _0945_ = \u0.u_issue.pipe_rd_wb_w  == 5'h1d;
  assign _0946_ = \u0.u_issue.pipe_rd_wb_w  == 5'h1e;
  assign _0947_ = \u0.u_issue.pipe_rd_wb_w  == 5'h1f;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r1_q  <= _0896_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r2_q  <= _0907_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r3_q  <= _0910_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r4_q  <= _0911_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r5_q  <= _0912_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r6_q  <= _0913_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r7_q  <= _0914_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r8_q  <= _0915_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r9_q  <= _0916_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r10_q  <= _0886_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r11_q  <= _0887_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r12_q  <= _0888_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r13_q  <= _0889_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r14_q  <= _0890_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r15_q  <= _0891_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r16_q  <= _0892_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r17_q  <= _0893_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r18_q  <= _0894_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r19_q  <= _0895_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r20_q  <= _0897_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r21_q  <= _0898_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r22_q  <= _0899_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r23_q  <= _0900_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r24_q  <= _0901_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r25_q  <= _0902_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r26_q  <= _0903_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r27_q  <= _0904_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r28_q  <= _0905_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r29_q  <= _0906_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r30_q  <= _0908_;
  always @(posedge clk_i)
    \u0.u_issue.u_regfile.REGFILE.reg_r31_q  <= _0909_;
  function [31:0] _2423_;
    input [31:0] a;
    input [991:0] b;
    input [30:0] s;
    casez (s) // synopsys parallel_case
      31'b??????????????????????????????1:
        _2423_ = b[31:0];
      31'b?????????????????????????????1?:
        _2423_ = b[63:32];
      31'b????????????????????????????1??:
        _2423_ = b[95:64];
      31'b???????????????????????????1???:
        _2423_ = b[127:96];
      31'b??????????????????????????1????:
        _2423_ = b[159:128];
      31'b?????????????????????????1?????:
        _2423_ = b[191:160];
      31'b????????????????????????1??????:
        _2423_ = b[223:192];
      31'b???????????????????????1???????:
        _2423_ = b[255:224];
      31'b??????????????????????1????????:
        _2423_ = b[287:256];
      31'b?????????????????????1?????????:
        _2423_ = b[319:288];
      31'b????????????????????1??????????:
        _2423_ = b[351:320];
      31'b???????????????????1???????????:
        _2423_ = b[383:352];
      31'b??????????????????1????????????:
        _2423_ = b[415:384];
      31'b?????????????????1?????????????:
        _2423_ = b[447:416];
      31'b????????????????1??????????????:
        _2423_ = b[479:448];
      31'b???????????????1???????????????:
        _2423_ = b[511:480];
      31'b??????????????1????????????????:
        _2423_ = b[543:512];
      31'b?????????????1?????????????????:
        _2423_ = b[575:544];
      31'b????????????1??????????????????:
        _2423_ = b[607:576];
      31'b???????????1???????????????????:
        _2423_ = b[639:608];
      31'b??????????1????????????????????:
        _2423_ = b[671:640];
      31'b?????????1?????????????????????:
        _2423_ = b[703:672];
      31'b????????1??????????????????????:
        _2423_ = b[735:704];
      31'b???????1???????????????????????:
        _2423_ = b[767:736];
      31'b??????1????????????????????????:
        _2423_ = b[799:768];
      31'b?????1?????????????????????????:
        _2423_ = b[831:800];
      31'b????1??????????????????????????:
        _2423_ = b[863:832];
      31'b???1???????????????????????????:
        _2423_ = b[895:864];
      31'b??1????????????????????????????:
        _2423_ = b[927:896];
      31'b?1?????????????????????????????:
        _2423_ = b[959:928];
      31'b1??????????????????????????????:
        _2423_ = b[991:960];
      default:
        _2423_ = a;
    endcase
  endfunction
  assign \u0.u_issue.issue_rb_value_w  = _2423_(32'h00000000, { \u0.u_issue.u_regfile.REGFILE.reg_r1_q , \u0.u_issue.u_regfile.REGFILE.reg_r2_q , \u0.u_issue.u_regfile.REGFILE.reg_r3_q , \u0.u_issue.u_regfile.REGFILE.reg_r4_q , \u0.u_issue.u_regfile.REGFILE.reg_r5_q , \u0.u_issue.u_regfile.REGFILE.reg_r6_q , \u0.u_issue.u_regfile.REGFILE.reg_r7_q , \u0.u_issue.u_regfile.REGFILE.reg_r8_q , \u0.u_issue.u_regfile.REGFILE.reg_r9_q , \u0.u_issue.u_regfile.REGFILE.reg_r10_q , \u0.u_issue.u_regfile.REGFILE.reg_r11_q , \u0.u_issue.u_regfile.REGFILE.reg_r12_q , \u0.u_issue.u_regfile.REGFILE.reg_r13_q , \u0.u_issue.u_regfile.REGFILE.reg_r14_q , \u0.u_issue.u_regfile.REGFILE.reg_r15_q , \u0.u_issue.u_regfile.REGFILE.reg_r16_q , \u0.u_issue.u_regfile.REGFILE.reg_r17_q , \u0.u_issue.u_regfile.REGFILE.reg_r18_q , \u0.u_issue.u_regfile.REGFILE.reg_r19_q , \u0.u_issue.u_regfile.REGFILE.reg_r20_q , \u0.u_issue.u_regfile.REGFILE.reg_r21_q , \u0.u_issue.u_regfile.REGFILE.reg_r22_q , \u0.u_issue.u_regfile.REGFILE.reg_r23_q , \u0.u_issue.u_regfile.REGFILE.reg_r24_q , \u0.u_issue.u_regfile.REGFILE.reg_r25_q , \u0.u_issue.u_regfile.REGFILE.reg_r26_q , \u0.u_issue.u_regfile.REGFILE.reg_r27_q , \u0.u_issue.u_regfile.REGFILE.reg_r28_q , \u0.u_issue.u_regfile.REGFILE.reg_r29_q , \u0.u_issue.u_regfile.REGFILE.reg_r30_q , \u0.u_issue.u_regfile.REGFILE.reg_r31_q  }, { _0978_, _0977_, _0976_, _0975_, _0974_, _0973_, _0972_, _0971_, _0970_, _0969_, _0968_, _0967_, _0966_, _0965_, _0964_, _0963_, _0962_, _0961_, _0960_, _0959_, _0958_, _0957_, _0956_, _0955_, _0954_, _0953_, _0952_, _0951_, _0950_, _0949_, _0948_ });
  assign _0948_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h1f;
  assign _0949_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h1e;
  assign _0950_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h1d;
  assign _0951_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h1c;
  assign _0952_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h1b;
  assign _0953_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h1a;
  assign _0954_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h19;
  assign _0955_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h18;
  assign _0956_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h17;
  assign _0957_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h16;
  assign _0958_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h15;
  assign _0959_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h14;
  assign _0960_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h13;
  assign _0961_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h12;
  assign _0962_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h11;
  assign _0963_ = \u0.u_csr.opcode_opcode_i [24:20] == 5'h10;
  assign _0964_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'hf;
  assign _0965_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'he;
  assign _0966_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'hd;
  assign _0967_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'hc;
  assign _0968_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'hb;
  assign _0969_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'ha;
  assign _0970_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'h9;
  assign _0971_ = \u0.u_csr.opcode_opcode_i [24:20] == 4'h8;
  assign _0972_ = \u0.u_csr.opcode_opcode_i [24:20] == 3'h7;
  assign _0973_ = \u0.u_csr.opcode_opcode_i [24:20] == 3'h6;
  assign _0974_ = \u0.u_csr.opcode_opcode_i [24:20] == 3'h5;
  assign _0975_ = \u0.u_csr.opcode_opcode_i [24:20] == 3'h4;
  assign _0976_ = \u0.u_csr.opcode_opcode_i [24:20] == 2'h3;
  assign _0977_ = \u0.u_csr.opcode_opcode_i [24:20] == 2'h2;
  assign _0978_ = \u0.u_csr.opcode_opcode_i [24:20] == 1'h1;
  function [31:0] _2455_;
    input [31:0] a;
    input [991:0] b;
    input [30:0] s;
    casez (s) // synopsys parallel_case
      31'b??????????????????????????????1:
        _2455_ = b[31:0];
      31'b?????????????????????????????1?:
        _2455_ = b[63:32];
      31'b????????????????????????????1??:
        _2455_ = b[95:64];
      31'b???????????????????????????1???:
        _2455_ = b[127:96];
      31'b??????????????????????????1????:
        _2455_ = b[159:128];
      31'b?????????????????????????1?????:
        _2455_ = b[191:160];
      31'b????????????????????????1??????:
        _2455_ = b[223:192];
      31'b???????????????????????1???????:
        _2455_ = b[255:224];
      31'b??????????????????????1????????:
        _2455_ = b[287:256];
      31'b?????????????????????1?????????:
        _2455_ = b[319:288];
      31'b????????????????????1??????????:
        _2455_ = b[351:320];
      31'b???????????????????1???????????:
        _2455_ = b[383:352];
      31'b??????????????????1????????????:
        _2455_ = b[415:384];
      31'b?????????????????1?????????????:
        _2455_ = b[447:416];
      31'b????????????????1??????????????:
        _2455_ = b[479:448];
      31'b???????????????1???????????????:
        _2455_ = b[511:480];
      31'b??????????????1????????????????:
        _2455_ = b[543:512];
      31'b?????????????1?????????????????:
        _2455_ = b[575:544];
      31'b????????????1??????????????????:
        _2455_ = b[607:576];
      31'b???????????1???????????????????:
        _2455_ = b[639:608];
      31'b??????????1????????????????????:
        _2455_ = b[671:640];
      31'b?????????1?????????????????????:
        _2455_ = b[703:672];
      31'b????????1??????????????????????:
        _2455_ = b[735:704];
      31'b???????1???????????????????????:
        _2455_ = b[767:736];
      31'b??????1????????????????????????:
        _2455_ = b[799:768];
      31'b?????1?????????????????????????:
        _2455_ = b[831:800];
      31'b????1??????????????????????????:
        _2455_ = b[863:832];
      31'b???1???????????????????????????:
        _2455_ = b[895:864];
      31'b??1????????????????????????????:
        _2455_ = b[927:896];
      31'b?1?????????????????????????????:
        _2455_ = b[959:928];
      31'b1??????????????????????????????:
        _2455_ = b[991:960];
      default:
        _2455_ = a;
    endcase
  endfunction
  assign \u0.u_issue.issue_ra_value_w  = _2455_(32'h00000000, { \u0.u_issue.u_regfile.REGFILE.reg_r1_q , \u0.u_issue.u_regfile.REGFILE.reg_r2_q , \u0.u_issue.u_regfile.REGFILE.reg_r3_q , \u0.u_issue.u_regfile.REGFILE.reg_r4_q , \u0.u_issue.u_regfile.REGFILE.reg_r5_q , \u0.u_issue.u_regfile.REGFILE.reg_r6_q , \u0.u_issue.u_regfile.REGFILE.reg_r7_q , \u0.u_issue.u_regfile.REGFILE.reg_r8_q , \u0.u_issue.u_regfile.REGFILE.reg_r9_q , \u0.u_issue.u_regfile.REGFILE.reg_r10_q , \u0.u_issue.u_regfile.REGFILE.reg_r11_q , \u0.u_issue.u_regfile.REGFILE.reg_r12_q , \u0.u_issue.u_regfile.REGFILE.reg_r13_q , \u0.u_issue.u_regfile.REGFILE.reg_r14_q , \u0.u_issue.u_regfile.REGFILE.reg_r15_q , \u0.u_issue.u_regfile.REGFILE.reg_r16_q , \u0.u_issue.u_regfile.REGFILE.reg_r17_q , \u0.u_issue.u_regfile.REGFILE.reg_r18_q , \u0.u_issue.u_regfile.REGFILE.reg_r19_q , \u0.u_issue.u_regfile.REGFILE.reg_r20_q , \u0.u_issue.u_regfile.REGFILE.reg_r21_q , \u0.u_issue.u_regfile.REGFILE.reg_r22_q , \u0.u_issue.u_regfile.REGFILE.reg_r23_q , \u0.u_issue.u_regfile.REGFILE.reg_r24_q , \u0.u_issue.u_regfile.REGFILE.reg_r25_q , \u0.u_issue.u_regfile.REGFILE.reg_r26_q , \u0.u_issue.u_regfile.REGFILE.reg_r27_q , \u0.u_issue.u_regfile.REGFILE.reg_r28_q , \u0.u_issue.u_regfile.REGFILE.reg_r29_q , \u0.u_issue.u_regfile.REGFILE.reg_r30_q , \u0.u_issue.u_regfile.REGFILE.reg_r31_q  }, { _1009_, _1008_, _1007_, _1006_, _1005_, _1004_, _1003_, _1002_, _1001_, _1000_, _0999_, _0998_, _0997_, _0996_, _0995_, _0994_, _0993_, _0992_, _0991_, _0990_, _0989_, _0988_, _0987_, _0986_, _0985_, _0984_, _0983_, _0982_, _0981_, _0980_, _0979_ });
  assign _0979_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h1f;
  assign _0980_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h1e;
  assign _0981_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h1d;
  assign _0982_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h1c;
  assign _0983_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h1b;
  assign _0984_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h1a;
  assign _0985_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h19;
  assign _0986_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h18;
  assign _0987_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h17;
  assign _0988_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h16;
  assign _0989_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h15;
  assign _0990_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h14;
  assign _0991_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h13;
  assign _0992_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h12;
  assign _0993_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h11;
  assign _0994_ = \u0.u_csr.opcode_opcode_i [19:15] == 5'h10;
  assign _0995_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'hf;
  assign _0996_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'he;
  assign _0997_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'hd;
  assign _0998_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'hc;
  assign _0999_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'hb;
  assign _1000_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'ha;
  assign _1001_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'h9;
  assign _1002_ = \u0.u_csr.opcode_opcode_i [19:15] == 4'h8;
  assign _1003_ = \u0.u_csr.opcode_opcode_i [19:15] == 3'h7;
  assign _1004_ = \u0.u_csr.opcode_opcode_i [19:15] == 3'h6;
  assign _1005_ = \u0.u_csr.opcode_opcode_i [19:15] == 3'h5;
  assign _1006_ = \u0.u_csr.opcode_opcode_i [19:15] == 3'h4;
  assign _1007_ = \u0.u_csr.opcode_opcode_i [19:15] == 2'h3;
  assign _1008_ = \u0.u_csr.opcode_opcode_i [19:15] == 2'h2;
  assign _1009_ = \u0.u_csr.opcode_opcode_i [19:15] == 1'h1;
  assign _1010_ = _0947_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r31_q ;
  assign _0909_ = rst_i ? 32'h00000000 : _1010_;
  assign _1011_ = _0946_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r30_q ;
  assign _0908_ = rst_i ? 32'h00000000 : _1011_;
  assign _1012_ = _0945_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r29_q ;
  assign _0906_ = rst_i ? 32'h00000000 : _1012_;
  assign _1013_ = _0944_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r28_q ;
  assign _0905_ = rst_i ? 32'h00000000 : _1013_;
  assign _1014_ = _0943_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r27_q ;
  assign _0904_ = rst_i ? 32'h00000000 : _1014_;
  assign _1015_ = _0942_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r26_q ;
  assign _0903_ = rst_i ? 32'h00000000 : _1015_;
  assign _1016_ = _0941_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r25_q ;
  assign _0902_ = rst_i ? 32'h00000000 : _1016_;
  assign _1017_ = _0940_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r24_q ;
  assign _0901_ = rst_i ? 32'h00000000 : _1017_;
  assign _1018_ = _0939_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r23_q ;
  assign _0900_ = rst_i ? 32'h00000000 : _1018_;
  assign _1019_ = _0938_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r22_q ;
  assign _0899_ = rst_i ? 32'h00000000 : _1019_;
  assign _1020_ = _0937_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r21_q ;
  assign _0898_ = rst_i ? 32'h00000000 : _1020_;
  assign _1021_ = _0936_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r20_q ;
  assign _0897_ = rst_i ? 32'h00000000 : _1021_;
  assign _1022_ = _0935_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r19_q ;
  assign _0895_ = rst_i ? 32'h00000000 : _1022_;
  assign _1023_ = _0934_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r18_q ;
  assign _0894_ = rst_i ? 32'h00000000 : _1023_;
  assign _1024_ = _0933_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r17_q ;
  assign _0893_ = rst_i ? 32'h00000000 : _1024_;
  assign _1025_ = _0932_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r16_q ;
  assign _0892_ = rst_i ? 32'h00000000 : _1025_;
  assign _1026_ = _0931_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r15_q ;
  assign _0891_ = rst_i ? 32'h00000000 : _1026_;
  assign _1027_ = _0930_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r14_q ;
  assign _0890_ = rst_i ? 32'h00000000 : _1027_;
  assign _1028_ = _0929_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r13_q ;
  assign _0889_ = rst_i ? 32'h00000000 : _1028_;
  assign _1029_ = _0928_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r12_q ;
  assign _0888_ = rst_i ? 32'h00000000 : _1029_;
  assign _1030_ = _0927_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r11_q ;
  assign _0887_ = rst_i ? 32'h00000000 : _1030_;
  assign _1031_ = _0926_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r10_q ;
  assign _0886_ = rst_i ? 32'h00000000 : _1031_;
  assign _1032_ = _0925_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r9_q ;
  assign _0916_ = rst_i ? 32'h00000000 : _1032_;
  assign _1033_ = _0924_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r8_q ;
  assign _0915_ = rst_i ? 32'h00000000 : _1033_;
  assign _1034_ = _0923_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r7_q ;
  assign _0914_ = rst_i ? 32'h00000000 : _1034_;
  assign _1035_ = _0922_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r6_q ;
  assign _0913_ = rst_i ? 32'h00000000 : _1035_;
  assign _1036_ = _0921_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r5_q ;
  assign _0912_ = rst_i ? 32'h00000000 : _1036_;
  assign _1037_ = _0920_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r4_q ;
  assign _0911_ = rst_i ? 32'h00000000 : _1037_;
  assign _1038_ = _0919_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r3_q ;
  assign _0910_ = rst_i ? 32'h00000000 : _1038_;
  assign _1039_ = _0918_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r2_q ;
  assign _0907_ = rst_i ? 32'h00000000 : _1039_;
  assign _1040_ = _0917_ ? \u0.u_issue.u_pipe_ctrl.result_wb_q  : \u0.u_issue.u_regfile.REGFILE.reg_r1_q ;
  assign _0896_ = rst_i ? 32'h00000000 : _1040_;
  assign _1072_ = \u0.u_csr.opcode_ra_operand_i  + { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] };
  assign _1073_ = \u0.u_csr.opcode_ra_operand_i  + { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:25], \u0.u_csr.opcode_opcode_i [11:7] };
  assign \u0.u_lsu.complete_ok_e2_w  = mem_d_ack_i & _1136_;
  assign \u0.u_lsu.complete_err_e2_w  = mem_d_ack_i & mem_d_error_i;
  assign _1074_ = \u0.u_lsu.mem_unaligned_e1_q  & _1137_;
  assign _1075_ = \u0.u_csr.opcode_opcode_i  & 15'h707f;
  assign _1076_ = \u0.u_csr.opcode_valid_i  & \u0.u_lsu.dcache_invalidate_w ;
  assign _1077_ = \u0.u_csr.opcode_valid_i  & \u0.u_lsu.dcache_writeback_w ;
  assign _1078_ = \u0.u_csr.opcode_valid_i  & \u0.u_lsu.dcache_flush_w ;
  assign \fifo_d_rd.in  = \u0.u_lsu.mem_rd_q  & _1137_;
  assign \u0.u_lsu.mem_wr_o  = \u0.u_lsu.mem_wr_q  & _1138_;
  assign \u0.u_lsu.fault_load_align_w  = \u0.u_lsu.mem_unaligned_e2_q  & \u0.u_lsu.u_lsu_request.data_out_o [0];
  assign \u0.u_lsu.fault_store_align_w  = \u0.u_lsu.mem_unaligned_e2_q  & _1139_;
  assign _1085_ = _1075_ == 2'h3;
  assign _1086_ = _1075_ == 13'h1003;
  assign _1087_ = _1075_ == 14'h2003;
  assign _1088_ = _1075_ == 15'h4003;
  assign _1089_ = _1075_ == 15'h5003;
  assign _1090_ = _1075_ == 15'h6003;
  assign \u0.u_lsu.req_sb_w  = _1075_ == 6'h23;
  assign \u0.u_lsu.req_sh_w  = _1075_ == 13'h1023;
  assign _1091_ = _1075_ == 14'h2023;
  assign _1092_ = _1075_ == 13'h1073;
  assign _1093_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h3a0;
  assign _1094_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h3a1;
  assign _1095_ = \u0.u_csr.opcode_opcode_i [31:20] == 10'h3a2;
  assign \u0.u_lsu.issue_lsu_e1_w  = _1118_ && mem_d_accept_i;
  assign \u0.u_lsu.delay_lsu_e2_w  = \u0.u_lsu.pending_lsu_e2_q  && _1112_;
  assign _1096_ = \u0.u_csr.opcode_valid_i  && _1092_;
  assign _1097_ = \u0.u_csr.opcode_valid_i  && \u0.u_lsu.load_inst_w ;
  assign _1098_ = \u0.u_csr.opcode_valid_i  && \u0.u_lsu.req_sw_lw_w ;
  assign _1099_ = \u0.u_csr.opcode_valid_i  && \u0.u_lsu.req_sh_lh_w ;
  assign \u0.u_lsu.mem_rd_r  = _1097_ && _1113_;
  assign _1100_ = \u0.u_csr.opcode_valid_i  && _1091_;
  assign _1101_ = _1100_ && _1113_;
  assign _1102_ = \u0.u_csr.opcode_valid_i  && \u0.u_lsu.req_sh_w ;
  assign _1103_ = _1102_ && _1113_;
  assign _1104_ = \u0.u_csr.opcode_valid_i  && \u0.u_lsu.req_sb_w ;
  assign \u0.u_lsu.dcache_flush_w  = _1092_ && _1093_;
  assign \u0.u_lsu.dcache_writeback_w  = _1092_ && _1094_;
  assign \u0.u_lsu.dcache_invalidate_w  = _1092_ && _1095_;
  assign _1105_ = _1127_ && \u0.u_lsu.delay_lsu_e2_w ;
  assign _1106_ = _1131_ && _1114_;
  assign _1107_ = \u0.u_lsu.mem_unaligned_e1_q  && _1137_;
  assign _1108_ = mem_d_ack_i && mem_d_error_i;
  assign _1109_ = mem_d_ack_i && \u0.u_lsu.u_lsu_request.data_out_o [0];
  assign _1110_ = \u0.u_lsu.u_lsu_request.data_out_o [3] && _1065_[7];
  assign _1111_ = \u0.u_lsu.u_lsu_request.data_out_o [3] && _1070_[15];
  assign \u0.u_lsu.fault_load_bus_w  = mem_d_error_i && \u0.u_lsu.u_lsu_request.data_out_o [0];
  assign \u0.u_lsu.fault_store_bus_w  = mem_d_error_i && _1139_;
  assign \u0.u_lsu.fault_load_page_w  = mem_d_error_i && 1'h0;
  assign \u0.u_lsu.fault_store_page_w  = mem_d_error_i && 1'h0;
  assign _1112_ = ! \u0.u_lsu.complete_ok_e2_w ;
  assign _1113_ = ! \u0.u_lsu.mem_unaligned_r ;
  assign _1114_ = ! mem_d_accept_i;
  assign _1115_ = \fifo_d_rd.in  || _1194_;
  assign _1116_ = _1115_ || \u0.u_lsu.mem_writeback_q ;
  assign _1117_ = _1116_ || \u0.u_lsu.mem_invalidate_q ;
  assign _1118_ = _1117_ || \u0.u_lsu.mem_flush_q ;
  assign _1119_ = \u0.u_lsu.complete_ok_e2_w  || \u0.u_lsu.complete_err_e2_w ;
  assign _1120_ = _1085_ || _1086_;
  assign \u0.u_lsu.load_signed_inst_w  = _1120_ || _1087_;
  assign _1121_ = \u0.u_lsu.load_signed_inst_w  || _1088_;
  assign _1122_ = _1121_ || _1089_;
  assign \u0.u_lsu.load_inst_w  = _1122_ || _1090_;
  assign \u0.u_lsu.req_lb_w  = _1085_ || _1088_;
  assign \u0.u_lsu.req_lh_w  = _1086_ || _1089_;
  assign _1123_ = _1091_ || _1087_;
  assign \u0.u_lsu.req_sw_lw_w  = _1123_ || _1090_;
  assign _1124_ = \u0.u_lsu.req_sh_w  || _1086_;
  assign \u0.u_lsu.req_sh_lh_w  = _1124_ || _1089_;
  assign _1125_ = \u0.u_lsu.complete_err_e2_w  || \u0.u_lsu.mem_unaligned_e2_q ;
  assign _1126_ = \u0.u_lsu.mem_rd_q  || _1195_;
  assign _1127_ = _1126_ || \u0.u_lsu.mem_unaligned_e1_q ;
  assign _1128_ = \u0.u_lsu.mem_writeback_q  || \u0.u_lsu.mem_invalidate_q ;
  assign _1129_ = _1128_ || \u0.u_lsu.mem_flush_q ;
  assign _1130_ = _1129_ || \fifo_d_rd.in ;
  assign _1131_ = _1130_ || _1135_;
  assign _1132_ = _1106_ || \u0.u_lsu.delay_lsu_e2_w ;
  assign \u0.u_issue.lsu_stall_i  = _1132_ || \u0.u_lsu.mem_unaligned_e1_q ;
  assign \u0.u_lsu.u_lsu_request.push_i  = \u0.u_lsu.issue_lsu_e1_w  || _1107_;
  assign \u0.u_lsu.u_lsu_request.pop_i  = mem_d_ack_i || \u0.u_lsu.mem_unaligned_e2_q ;
  assign _1133_ = _1108_ || \u0.u_lsu.mem_unaligned_e2_q ;
  assign _1134_ = | \u0.u_lsu.mem_addr_r [1:0];
  assign _1135_ = | \u0.u_lsu.mem_wr_o ;
  assign _1136_ = ~ mem_d_error_i;
  assign _1137_ = ~ \u0.u_lsu.delay_lsu_e2_w ;
  assign _1138_ = ~ { \u0.u_lsu.delay_lsu_e2_w , \u0.u_lsu.delay_lsu_e2_w , \u0.u_lsu.delay_lsu_e2_w , \u0.u_lsu.delay_lsu_e2_w  };
  assign _1139_ = ~ \u0.u_lsu.u_lsu_request.data_out_o [0];
  assign _1140_ = \u0.u_lsu.req_lb_w  | \u0.u_lsu.req_sb_w ;
  assign _1141_ = \u0.u_lsu.req_lh_w  | \u0.u_lsu.req_sh_w ;
  assign \u0.u_issue.u_pipe_ctrl.mem_complete_i  = mem_d_ack_i | \u0.u_lsu.mem_unaligned_e2_q ;
  always @(posedge clk_i)
    \u0.u_lsu.mem_addr_q  <= _1041_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_data_wr_q  <= _1042_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_rd_q  <= _1047_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_wr_q  <= _1050_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_invalidate_q  <= _1044_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_writeback_q  <= _1051_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_flush_q  <= _1043_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_unaligned_e1_q  <= _1048_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_load_q  <= _1045_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_xb_q  <= _1052_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_xh_q  <= _1053_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_ls_q  <= _1046_;
  always @(posedge clk_i)
    \u0.u_lsu.mem_unaligned_e2_q  <= _1049_;
  always @(posedge clk_i)
    \u0.u_lsu.pending_lsu_e2_q  <= _1054_;
  assign _1071_ = _1111_ ? { 16'hffff, _1070_[15:0] } : _1070_;
  assign _1079_[15:0] = \u0.u_lsu.u_lsu_request.data_out_o [5] ? mem_d_data_rd_i[31:16] : mem_d_data_rd_i[15:0];
  assign _1142_ = \u0.u_lsu.u_lsu_request.data_out_o [2] ? { 16'h0000, _1079_[15:0] } : 32'hxxxxxxxx;
  assign _1143_ = \u0.u_lsu.u_lsu_request.data_out_o [1] ? 32'hxxxxxxxx : _1142_;
  assign _1144_ = _1109_ ? _1143_ : 32'hxxxxxxxx;
  assign _1070_ = _1133_ ? 32'hxxxxxxxx : _1144_;
  assign _1069_ = \u0.u_lsu.u_lsu_request.data_out_o [2] ? _1071_ : mem_d_data_rd_i;
  assign _1068_ = _1110_ ? { 24'hffffff, _1065_[7:0] } : _1065_;
  function [31:0] _2663_;
    input [31:0] a;
    input [127:0] b;
    input [3:0] s;
    casez (s) // synopsys parallel_case
      4'b???1:
        _2663_ = b[31:0];
      4'b??1?:
        _2663_ = b[63:32];
      4'b?1??:
        _2663_ = b[95:64];
      4'b1???:
        _2663_ = b[127:96];
      default:
        _2663_ = a;
    endcase
  endfunction
  assign _1145_ = _2663_(32'hxxxxxxxx, { 24'h000000, mem_d_data_rd_i[31:24], 24'h000000, mem_d_data_rd_i[23:16], 24'h000000, mem_d_data_rd_i[15:8], 24'h000000, mem_d_data_rd_i[7:0] }, { _1149_, _1148_, _1147_, _1146_ });
  assign _1146_ = ! \u0.u_lsu.u_lsu_request.data_out_o [5:4];
  assign _1147_ = \u0.u_lsu.u_lsu_request.data_out_o [5:4] == 1'h1;
  assign _1148_ = \u0.u_lsu.u_lsu_request.data_out_o [5:4] == 2'h2;
  assign _1149_ = \u0.u_lsu.u_lsu_request.data_out_o [5:4] == 2'h3;
  assign _1150_ = \u0.u_lsu.u_lsu_request.data_out_o [1] ? _1145_ : 32'hxxxxxxxx;
  assign _1151_ = _1109_ ? _1150_ : 32'hxxxxxxxx;
  assign _1065_ = _1133_ ? 32'hxxxxxxxx : _1151_;
  assign _1062_ = \u0.u_lsu.u_lsu_request.data_out_o [1] ? _1068_ : _1069_;
  assign _1059_ = _1109_ ? _1062_ : 32'h00000000;
  assign \u0.u_issue.u_pipe_ctrl.mem_result_e2_i  = _1133_ ? \u0.u_lsu.u_lsu_request.data_out_o [35:4] : _1059_;
  assign _1152_ = _1106_ ? \u0.u_lsu.mem_ls_q  : \u0.u_lsu.load_signed_inst_w ;
  assign _1153_ = _1105_ ? \u0.u_lsu.mem_ls_q  : _1152_;
  assign _1154_ = _1125_ ? 1'h0 : _1153_;
  assign _1046_ = rst_i ? 1'h0 : _1154_;
  assign _1155_ = _1106_ ? \u0.u_lsu.mem_xh_q  : _1141_;
  assign _1156_ = _1105_ ? \u0.u_lsu.mem_xh_q  : _1155_;
  assign _1157_ = _1125_ ? 1'h0 : _1156_;
  assign _1053_ = rst_i ? 1'h0 : _1157_;
  assign _1158_ = _1106_ ? \u0.u_lsu.mem_xb_q  : _1140_;
  assign _1159_ = _1105_ ? \u0.u_lsu.mem_xb_q  : _1158_;
  assign _1160_ = _1125_ ? 1'h0 : _1159_;
  assign _1052_ = rst_i ? 1'h0 : _1160_;
  assign _1161_ = _1106_ ? \u0.u_lsu.mem_load_q  : _1097_;
  assign _1162_ = _1105_ ? \u0.u_lsu.mem_load_q  : _1161_;
  assign _1163_ = _1125_ ? 1'h0 : _1162_;
  assign _1045_ = rst_i ? 1'h0 : _1163_;
  assign _1164_ = _1106_ ? \u0.u_lsu.mem_unaligned_e1_q  : \u0.u_lsu.mem_unaligned_r ;
  assign _1165_ = _1105_ ? \u0.u_lsu.mem_unaligned_e1_q  : _1164_;
  assign _1166_ = _1125_ ? 1'h0 : _1165_;
  assign _1048_ = rst_i ? 1'h0 : _1166_;
  assign _1167_ = _1106_ ? \u0.u_lsu.mem_flush_q  : _1078_;
  assign _1168_ = _1105_ ? \u0.u_lsu.mem_flush_q  : _1167_;
  assign _1169_ = _1125_ ? 1'h0 : _1168_;
  assign _1043_ = rst_i ? 1'h0 : _1169_;
  assign _1170_ = _1106_ ? \u0.u_lsu.mem_writeback_q  : _1077_;
  assign _1171_ = _1105_ ? \u0.u_lsu.mem_writeback_q  : _1170_;
  assign _1172_ = _1125_ ? 1'h0 : _1171_;
  assign _1051_ = rst_i ? 1'h0 : _1172_;
  assign _1173_ = _1106_ ? \u0.u_lsu.mem_invalidate_q  : _1076_;
  assign _1174_ = _1105_ ? \u0.u_lsu.mem_invalidate_q  : _1173_;
  assign _1175_ = _1125_ ? 1'h0 : _1174_;
  assign _1044_ = rst_i ? 1'h0 : _1175_;
  assign _1176_ = _1106_ ? \u0.u_lsu.mem_wr_q  : \u0.u_lsu.mem_wr_r ;
  assign _1177_ = _1105_ ? \u0.u_lsu.mem_wr_q  : _1176_;
  assign _1178_ = _1125_ ? 4'h0 : _1177_;
  assign _1050_ = rst_i ? 4'h0 : _1178_;
  assign _1179_ = _1106_ ? \u0.u_lsu.mem_rd_q  : \u0.u_lsu.mem_rd_r ;
  assign _1180_ = _1105_ ? \u0.u_lsu.mem_rd_q  : _1179_;
  assign _1181_ = _1125_ ? 1'h0 : _1180_;
  assign _1047_ = rst_i ? 1'h0 : _1181_;
  assign _1182_ = _1106_ ? \u0.u_lsu.mem_data_wr_q  : \u0.u_lsu.mem_data_r ;
  assign _1183_ = _1105_ ? \u0.u_lsu.mem_data_wr_q  : _1182_;
  assign _1184_ = _1125_ ? 32'h00000000 : _1183_;
  assign _1042_ = rst_i ? 32'h00000000 : _1184_;
  assign _1185_ = _1106_ ? \u0.u_lsu.mem_addr_q  : \u0.u_lsu.mem_addr_r ;
  assign _1186_ = _1105_ ? \u0.u_lsu.mem_addr_q  : _1185_;
  assign _1187_ = _1125_ ? 32'h00000000 : _1186_;
  assign _1041_ = rst_i ? 32'h00000000 : _1187_;
  function [3:0] _2722_;
    input [3:0] a;
    input [15:0] b;
    input [3:0] s;
    casez (s) // synopsys parallel_case
      4'b???1:
        _2722_ = b[3:0];
      4'b??1?:
        _2722_ = b[7:4];
      4'b?1??:
        _2722_ = b[11:8];
      4'b1???:
        _2722_ = b[15:12];
      default:
        _2722_ = a;
    endcase
  endfunction
  assign _1067_ = _2722_(4'hx, 16'h8421, { _1191_, _1190_, _1189_, _1188_ });
  assign _1188_ = ! \u0.u_lsu.mem_addr_r [1:0];
  assign _1189_ = \u0.u_lsu.mem_addr_r [1:0] == 1'h1;
  assign _1190_ = \u0.u_lsu.mem_addr_r [1:0] == 2'h2;
  assign _1191_ = \u0.u_lsu.mem_addr_r [1:0] == 2'h3;
  function [31:0] _2727_;
    input [31:0] a;
    input [127:0] b;
    input [3:0] s;
    casez (s) // synopsys parallel_case
      4'b???1:
        _2727_ = b[31:0];
      4'b??1?:
        _2727_ = b[63:32];
      4'b?1??:
        _2727_ = b[95:64];
      4'b1???:
        _2727_ = b[127:96];
      default:
        _2727_ = a;
    endcase
  endfunction
  assign _1066_ = _2727_(32'hxxxxxxxx, { \u0.u_div.opcode_rb_operand_i [7:0], 32'h00000000, \u0.u_div.opcode_rb_operand_i [7:0], 32'h00000000, \u0.u_div.opcode_rb_operand_i [7:0], 32'h00000000, \u0.u_div.opcode_rb_operand_i [7:0] }, { _1191_, _1190_, _1189_, _1188_ });
  assign _1064_ = _1104_ ? _1067_ : 4'h0;
  assign _1063_ = _1104_ ? _1066_ : 32'h00000000;
  assign _1061_ = _1190_ ? 4'hc : 4'h3;
  assign _1060_ = _1190_ ? { \u0.u_div.opcode_rb_operand_i [15:0], 16'h0000 } : { 16'h0000, \u0.u_div.opcode_rb_operand_i [15:0] };
  assign _1058_ = _1103_ ? _1061_ : _1064_;
  assign _1056_ = _1103_ ? _1060_ : _1063_;
  assign \u0.u_lsu.mem_wr_r  = _1101_ ? 4'hf : _1058_;
  assign \u0.u_lsu.mem_data_r  = _1101_ ? \u0.u_div.opcode_rb_operand_i  : _1056_;
  assign _1057_ = _1099_ ? \u0.u_lsu.mem_addr_r [0] : 1'h0;
  assign \u0.u_lsu.mem_unaligned_r  = _1098_ ? _1134_ : _1057_;
  assign _1055_ = _1097_ ? _1072_ : _1073_;
  assign \u0.u_lsu.mem_addr_r  = _1096_ ? \u0.u_csr.opcode_ra_operand_i  : _1055_;
  assign _1049_ = rst_i ? 1'h0 : _1074_;
  assign _1192_ = _1119_ ? 1'h0 : \u0.u_lsu.pending_lsu_e2_q ;
  assign _1193_ = \u0.u_lsu.issue_lsu_e1_w  ? 1'h1 : _1192_;
  assign _1054_ = rst_i ? 1'h0 : _1193_;
  assign _1194_ = | \u0.u_lsu.mem_wr_o ;
  assign _1195_ = | \u0.u_lsu.mem_wr_q ;
  assign \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i [4:0] = \u0.u_lsu.fault_load_align_w  ? 5'h14 : _1080_[4:0];
  assign _1080_[4:0] = \u0.u_lsu.fault_store_align_w  ? 5'h16 : _1081_[4:0];
  assign _1081_[4:0] = \u0.u_lsu.fault_load_page_w  ? 5'h1d : _1082_[4:0];
  assign _1082_[4:0] = \u0.u_lsu.fault_store_page_w  ? 5'h1f : _1083_[4:0];
  assign _1083_[4:0] = \u0.u_lsu.fault_load_bus_w  ? 5'h15 : _1084_[4:0];
  assign _1084_[4:0] = \u0.u_lsu.fault_store_bus_w  ? 5'h17 : 5'h00;
  assign _1203_ = \u0.u_lsu.u_lsu_request.wr_ptr_q  + 1'h1;
  assign _1204_[0] = \u0.u_lsu.u_lsu_request.rd_ptr_q  + 1'h1;
  assign _1205_[1:0] = \u0.u_lsu.u_lsu_request.count_q  + 1'h1;
  assign _1206_ = \u0.u_lsu.u_lsu_request.push_i  & \u0.u_lsu.u_lsu_request.accept_o ;
  assign _1207_ = \u0.u_lsu.u_lsu_request.pop_i  & \u0.u_lsu.u_lsu_request.valid_o ;
  assign _1208_ = _1206_ & _1210_;
  assign _1209_ = _1211_ & _1207_;
  assign \u0.u_lsu.u_lsu_request.valid_o  = | \u0.u_lsu.u_lsu_request.count_q ;
  assign \u0.u_lsu.u_lsu_request.accept_o  = \u0.u_lsu.u_lsu_request.count_q  != 2'h2;
  assign _1210_ = ~ _1207_;
  assign _1211_ = ~ _1206_;
  always @(posedge clk_i)
    \u0.u_lsu.u_lsu_request.rd_ptr_q  <= _1201_;
  always @(posedge clk_i)
    \u0.u_lsu.u_lsu_request.wr_ptr_q  <= _1202_;
  always @(posedge clk_i)
    \u0.u_lsu.u_lsu_request.count_q  <= _1200_;
  assign _1196_[35] = rst_i ? 1'h1 : 1'h0;
  assign _1212_[35] = _1206_ ? 1'h1 : 1'h0;
  assign _1199_[35] = rst_i ? 1'h0 : _1212_[35];
  assign _1213_ = _1206_ ? { \u0.u_lsu.mem_addr_q , \u0.u_lsu.mem_ls_q , \u0.u_lsu.mem_xh_q , \u0.u_lsu.mem_xb_q , \u0.u_lsu.mem_load_q  } : 36'hxxxxxxxxx;
  assign _1198_ = rst_i ? 36'hxxxxxxxxx : _1213_;
  assign _1214_ = _1206_ ? \u0.u_lsu.u_lsu_request.wr_ptr_q  : 1'hx;
  assign _1197_ = rst_i ? 1'hx : _1214_;
  assign _1215_ = _1209_ ? _1219_[1:0] : \u0.u_lsu.u_lsu_request.count_q ;
  assign _1216_ = _1208_ ? _1205_[1:0] : _1215_;
  assign _1200_ = rst_i ? 2'h0 : _1216_;
  assign _1217_ = _1206_ ? _1203_ : \u0.u_lsu.u_lsu_request.wr_ptr_q ;
  assign _1202_ = rst_i ? 1'h0 : _1217_;
  assign _1218_ = _1207_ ? _1204_[0] : \u0.u_lsu.u_lsu_request.rd_ptr_q ;
  assign _1201_ = rst_i ? 1'h0 : _1218_;
  assign _1219_[1:0] = \u0.u_lsu.u_lsu_request.count_q  - 1'h1;
  assign _1226_ = \u0.u_csr.opcode_opcode_i  & 32'hfe00707f;
  assign _1227_ = _1226_ == 26'h2002033;
  assign _1228_ = _1226_ == 26'h2001033;
  assign _1229_ = _1226_ == 26'h2000033;
  assign _1230_ = _1226_ == 26'h2003033;
  assign _1231_ = \u0.u_div.opcode_valid_i  && \u0.u_mul.mult_inst_w ;
  assign _1232_ = _1229_ || _1228_;
  assign _1233_ = _1232_ || _1227_;
  assign \u0.u_mul.mult_inst_w  = _1233_ || _1230_;
  assign \u0.u_mul.mult_result_w  = { \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q [32], \u0.u_mul.operand_a_e1_q  } * { \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q [32], \u0.u_mul.operand_b_e1_q  };
  assign _1234_ = ~ _1229_;
  always @(posedge clk_i)
    \u0.u_mul.result_e2_q  <= _1223_;
  always @(posedge clk_i)
    \u0.u_mul.operand_a_e1_q  <= _1221_;
  always @(posedge clk_i)
    \u0.u_mul.operand_b_e1_q  <= _1222_;
  always @(posedge clk_i)
    \u0.u_mul.mulhi_sel_e1_q  <= _1220_;
  assign _1235_ = \u0.u_exec.hold_i  ? \u0.u_mul.result_e2_q  : \u0.u_mul.result_r ;
  assign _1223_ = rst_i ? 32'h00000000 : _1235_;
  assign _1236_ = _1231_ ? _1234_ : 1'h0;
  assign _1237_ = \u0.u_exec.hold_i  ? \u0.u_mul.mulhi_sel_e1_q  : _1236_;
  assign _1220_ = rst_i ? 1'h0 : _1237_;
  assign _1238_ = _1231_ ? \u0.u_mul.operand_b_r  : 33'h000000000;
  assign _1239_ = \u0.u_exec.hold_i  ? \u0.u_mul.operand_b_e1_q  : _1238_;
  assign _1222_ = rst_i ? 33'h000000000 : _1239_;
  assign _1240_ = _1231_ ? \u0.u_mul.operand_a_r  : 33'h000000000;
  assign _1241_ = \u0.u_exec.hold_i  ? \u0.u_mul.operand_a_e1_q  : _1240_;
  assign _1221_ = rst_i ? 33'h000000000 : _1241_;
  assign _1225_ = _1228_ ? { \u0.u_div.opcode_rb_operand_i [31], \u0.u_div.opcode_rb_operand_i  } : { 1'h0, \u0.u_div.opcode_rb_operand_i  };
  assign \u0.u_mul.operand_b_r  = _1227_ ? { 1'h0, \u0.u_div.opcode_rb_operand_i  } : _1225_;
  assign _1224_ = _1228_ ? { \u0.u_csr.opcode_ra_operand_i [31], \u0.u_csr.opcode_ra_operand_i  } : { 1'h0, \u0.u_csr.opcode_ra_operand_i  };
  assign \u0.u_mul.operand_a_r  = _1227_ ? { \u0.u_csr.opcode_ra_operand_i [31], \u0.u_csr.opcode_ra_operand_i  } : _1224_;
  assign \u0.u_mul.result_r  = \u0.u_mul.mulhi_sel_e1_q  ? \u0.u_mul.mult_result_w [63:32] : \u0.u_mul.mult_result_w [31:0];
  assign \fifo_d_addr.wr  = \u0.u_lsu.mem_wr_o [0] || \fifo_d_rd.in ;
  assign \u0.u_lsu.u_lsu_request.data_out_o  = \u0.u_lsu.u_lsu_request.rd_ptr_q  ? \u0.u_lsu.u_lsu_request.ram_q[1]  : \u0.u_lsu.u_lsu_request.ram_q[0] ;
  assign _1242_ = _0000_ & _1196_[35];
  assign _1243_ = _0001_ & _1196_[35];
  assign _1244_ = _0002_ & _1199_[35];
  assign _1245_ = _0003_ & _1196_[35];
  assign _1246_ = _0004_ & _1196_[35];
  assign _1247_ = _0005_ & _1199_[35];
  assign _1248_ = _1242_ ? 36'h000000000 : \u0.u_lsu.u_lsu_request.ram_q[0] ;
  assign _1249_ = _1243_ ? 36'h000000000 : _1248_;
  assign _1250_ = _1244_ ? _1198_ : _1249_;
  assign _1251_ = _1245_ ? 36'h000000000 : \u0.u_lsu.u_lsu_request.ram_q[1] ;
  assign _1252_ = _1246_ ? 36'h000000000 : _1251_;
  assign _1253_ = _1247_ ? _1198_ : _1252_;
  always @(posedge clk_i)
    \u0.u_lsu.u_lsu_request.ram_q[0]  <= _1250_;
  always @(posedge clk_i)
    \u0.u_lsu.u_lsu_request.ram_q[1]  <= _1253_;
  assign _0641_[31:1] = 31'h00000000;
  assign _0648_[1] = _0642_;
  assign _0657_[31:1] = 31'h00000000;
  assign _0658_[31:1] = 31'h00000000;
  assign _0709_[5] = 1'h0;
  assign _0781_[5] = 1'h0;
  assign _1079_[31:16] = 16'h0000;
  assign _1080_[5] = 1'h0;
  assign _1081_[5] = 1'h0;
  assign _1082_[5] = 1'h0;
  assign _1083_[5] = 1'h0;
  assign _1084_[5] = 1'h0;
  assign _1196_[34:0] = { _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35], _1196_[35] };
  assign _1199_[34:0] = { _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35], _1199_[35] };
  assign _1212_[34:0] = { _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35], _1212_[35] };
  assign \fifo_d_addr.clk  = clk_i;
  assign \fifo_d_addr.in  = 32'h00000000;
  assign \fifo_d_addr.out  = \fifo_d_addr.r1 ;
  assign \fifo_d_addr.rst  = rst_i;
  assign \fifo_d_data_wr.clk  = clk_i;
  assign \fifo_d_data_wr.in  = { 31'h00000000, \u0.u_lsu.mem_data_wr_q [0] };
  assign \fifo_d_data_wr.out  = \fifo_d_data_wr.r1 ;
  assign \fifo_d_data_wr.rst  = rst_i;
  assign \fifo_d_data_wr.wr  = \u0.u_lsu.mem_wr_o [0];
  assign \fifo_d_rd.clk  = clk_i;
  assign \fifo_d_rd.out  = \fifo_d_rd.r1 ;
  assign \fifo_d_rd.rst  = rst_i;
  assign \fifo_d_rd.wr  = \fifo_d_rd.in ;
  assign \fifo_d_wr.clk  = clk_i;
  assign \fifo_d_wr.in  = { 3'h0, \u0.u_lsu.mem_wr_o [0] };
  assign \fifo_d_wr.out  = \fifo_d_wr.r1 ;
  assign \fifo_d_wr.rst  = rst_i;
  assign \fifo_d_wr.wr  = \u0.u_lsu.mem_wr_o [0];
  assign \fifo_i_pc.clk  = clk_i;
  assign \fifo_i_pc.in  = 32'h00000000;
  assign \fifo_i_pc.out  = \fifo_i_pc.r1 ;
  assign \fifo_i_pc.rst  = rst_i;
  assign \fifo_i_rd.clk  = clk_i;
  assign \fifo_i_rd.out  = \fifo_i_rd.r1 ;
  assign \fifo_i_rd.rst  = rst_i;
  assign \fifo_i_rd.wr  = \fifo_i_rd.in ;
  assign mem_d_addr_o = 1'h0;
  assign mem_d_addr_o_fifo = \fifo_d_addr.r1 ;
  assign mem_d_cacheable_o = \u0.mem_d_cacheable_o ;
  assign mem_d_data_wr_o = \u0.u_lsu.mem_data_wr_q [0];
  assign mem_d_data_wr_o_fifo = \fifo_d_data_wr.r1 ;
  assign mem_d_flush_o = \u0.u_lsu.mem_flush_q ;
  assign mem_d_invalidate_o = \u0.u_lsu.mem_invalidate_q ;
  assign mem_d_rd_o = \fifo_d_rd.in ;
  assign mem_d_rd_o_fifo = \fifo_d_rd.r1 ;
  assign mem_d_req_tag_o = 1'h0;
  assign mem_d_wr_o = \u0.u_lsu.mem_wr_o [0];
  assign mem_d_wr_o_fifo = \fifo_d_wr.r1 ;
  assign mem_d_writeback_o = \u0.u_lsu.mem_writeback_q ;
  assign mem_i_flush_o = \u0.ifence_w ;
  assign mem_i_invalidate_o = 1'h0;
  assign mem_i_pc_o = 1'h0;
  assign mem_i_pc_o_fifo = \fifo_i_pc.r1 ;
  assign mem_i_rd_o = \fifo_i_rd.in ;
  assign mem_i_rd_o_fifo = \fifo_i_rd.r1 ;
  assign \u0.branch_csr_pc_w  = \u0.u_csr.branch_target_q ;
  assign \u0.branch_csr_request_w  = \u0.u_csr.branch_q ;
  assign \u0.branch_d_exec_pc_w  = \u0.u_exec.branch_target_r ;
  assign \u0.branch_d_exec_priv_w  = 2'h0;
  assign \u0.branch_d_exec_request_w  = \u0.u_exec.branch_d_request_o ;
  assign \u0.branch_pc_w  = \u0.u_fetch.branch_pc_i ;
  assign \u0.branch_request_w  = \u0.u_fetch.branch_request_i ;
  assign \u0.clk_i  = clk_i;
  assign \u0.cpu_id_i  = cpu_id_i;
  assign \u0.csr_opcode_invalid_w  = \u0.u_csr.opcode_invalid_i ;
  assign \u0.csr_opcode_opcode_w  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.csr_opcode_pc_w  = \u0.u_exec.opcode_pc_i ;
  assign \u0.csr_opcode_ra_idx_w  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.csr_opcode_ra_operand_w  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.csr_opcode_rb_idx_w  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.csr_opcode_rb_operand_w  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.csr_opcode_rd_idx_w  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.csr_opcode_valid_w  = \u0.u_csr.opcode_valid_i ;
  assign \u0.csr_result_e1_exception_w  = \u0.u_csr.exception_e1_q ;
  assign \u0.csr_result_e1_value_w  = \u0.u_csr.rd_result_e1_q ;
  assign \u0.csr_result_e1_wdata_w  = \u0.u_csr.csr_wdata_e1_q ;
  assign \u0.csr_result_e1_write_w  = \u0.u_csr.rd_valid_e1_q ;
  assign \u0.csr_writeback_exception_addr_w  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.csr_writeback_exception_pc_w  = \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  assign \u0.csr_writeback_exception_w  = \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.csr_writeback_waddr_w  = \u0.u_issue.u_pipe_ctrl.opcode_wb_q [31:20];
  assign \u0.csr_writeback_wdata_w  = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q ;
  assign \u0.csr_writeback_write_w  = \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q ;
  assign \u0.div_opcode_valid_w  = \u0.u_div.opcode_valid_i ;
  assign \u0.exec_hold_w  = \u0.u_exec.hold_i ;
  assign \u0.exec_opcode_valid_w  = \u0.u_div.opcode_valid_i ;
  assign \u0.fetch_accept_w  = \u0.u_fetch.fetch_accept_i ;
  assign \u0.fetch_dec_accept_w  = \u0.u_fetch.fetch_accept_i ;
  assign \u0.fetch_dec_fault_fetch_w  = \u0.u_decode.fetch_in_fault_fetch_i ;
  assign \u0.fetch_dec_fault_page_w  = \u0.u_decode.fetch_in_fault_page_i ;
  assign \u0.fetch_dec_instr_w  = \u0.u_decode.fetch_in_instr_i ;
  assign \u0.fetch_dec_pc_w  = \u0.u_exec.opcode_pc_i ;
  assign \u0.fetch_dec_valid_w  = \u0.u_decode.genblk1.u_dec.valid_i ;
  assign \u0.fetch_fault_fetch_w  = \u0.u_decode.fetch_in_fault_fetch_i ;
  assign \u0.fetch_fault_page_w  = \u0.u_decode.fetch_in_fault_page_i ;
  assign \u0.fetch_in_fault_w  = 1'h0;
  assign \u0.fetch_instr_branch_w  = \u0.u_decode.genblk1.u_dec.branch_o ;
  assign \u0.fetch_instr_csr_w  = \u0.u_decode.genblk1.u_dec.csr_o ;
  assign \u0.fetch_instr_div_w  = \u0.u_decode.genblk1.u_dec.div_o ;
  assign \u0.fetch_instr_exec_w  = \u0.u_decode.genblk1.u_dec.exec_o ;
  assign \u0.fetch_instr_invalid_w  = \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign \u0.fetch_instr_lsu_w  = \u0.u_decode.genblk1.u_dec.lsu_o ;
  assign \u0.fetch_instr_mul_w  = \u0.u_decode.genblk1.u_dec.mul_o ;
  assign \u0.fetch_instr_rd_valid_w  = \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign \u0.fetch_instr_w  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.fetch_pc_w  = \u0.u_exec.opcode_pc_i ;
  assign \u0.fetch_valid_w  = \u0.u_decode.genblk1.u_dec.valid_i ;
  assign \u0.interrupt_inhibit_w  = \u0.u_csr.interrupt_inhibit_i ;
  assign \u0.intr_i  = intr_i;
  assign \u0.lsu_opcode_invalid_w  = 1'h0;
  assign \u0.lsu_opcode_opcode_w  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.lsu_opcode_pc_w  = \u0.u_exec.opcode_pc_i ;
  assign \u0.lsu_opcode_ra_idx_w  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.lsu_opcode_ra_operand_w  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.lsu_opcode_rb_idx_w  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.lsu_opcode_rb_operand_w  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.lsu_opcode_rd_idx_w  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.lsu_opcode_valid_w  = \u0.u_csr.opcode_valid_i ;
  assign \u0.lsu_stall_w  = \u0.u_issue.lsu_stall_i ;
  assign \u0.mem_d_accept_i  = mem_d_accept_i;
  assign \u0.mem_d_ack_i  = mem_d_ack_i;
  assign \u0.mem_d_addr_o  = { \u0.u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u0.mem_d_data_rd_i  = mem_d_data_rd_i;
  assign \u0.mem_d_data_wr_o  = \u0.u_lsu.mem_data_wr_q ;
  assign \u0.mem_d_error_i  = mem_d_error_i;
  assign \u0.mem_d_flush_o  = \u0.u_lsu.mem_flush_q ;
  assign \u0.mem_d_invalidate_o  = \u0.u_lsu.mem_invalidate_q ;
  assign \u0.mem_d_rd_o  = \fifo_d_rd.in ;
  assign \u0.mem_d_req_tag_o  = 11'h000;
  assign \u0.mem_d_resp_tag_i  = mem_d_resp_tag_i;
  assign \u0.mem_d_wr_o  = \u0.u_lsu.mem_wr_o ;
  assign \u0.mem_d_writeback_o  = \u0.u_lsu.mem_writeback_q ;
  assign \u0.mem_i_accept_i  = mem_i_accept_i;
  assign \u0.mem_i_error_i  = mem_i_error_i;
  assign \u0.mem_i_flush_o  = \u0.ifence_w ;
  assign \u0.mem_i_inst_i  = mem_i_inst_i;
  assign \u0.mem_i_invalidate_o  = 1'h0;
  assign \u0.mem_i_pc_o  = { \u0.u_fetch.pc_f_q [31:2], 2'h0 };
  assign \u0.mem_i_rd_o  = \fifo_i_rd.in ;
  assign \u0.mem_i_valid_i  = mem_i_valid_i;
  assign \u0.mmu_ifetch_accept_w  = mem_i_accept_i;
  assign \u0.mmu_ifetch_error_w  = mem_i_error_i;
  assign \u0.mmu_ifetch_flush_w  = \u0.ifence_w ;
  assign \u0.mmu_ifetch_inst_w  = mem_i_inst_i;
  assign \u0.mmu_ifetch_invalidate_w  = 1'h0;
  assign \u0.mmu_ifetch_pc_w  = { \u0.u_fetch.pc_f_q [31:2], 2'h0 };
  assign \u0.mmu_ifetch_rd_w  = \fifo_i_rd.in ;
  assign \u0.mmu_ifetch_valid_w  = mem_i_valid_i;
  assign \u0.mmu_load_fault_w  = 1'h0;
  assign \u0.mmu_lsu_accept_w  = mem_d_accept_i;
  assign \u0.mmu_lsu_ack_w  = mem_d_ack_i;
  assign \u0.mmu_lsu_addr_w  = { \u0.u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u0.mmu_lsu_cacheable_w  = \u0.mem_d_cacheable_o ;
  assign \u0.mmu_lsu_data_rd_w  = mem_d_data_rd_i;
  assign \u0.mmu_lsu_data_wr_w  = \u0.u_lsu.mem_data_wr_q ;
  assign \u0.mmu_lsu_error_w  = mem_d_error_i;
  assign \u0.mmu_lsu_flush_w  = \u0.u_lsu.mem_flush_q ;
  assign \u0.mmu_lsu_invalidate_w  = \u0.u_lsu.mem_invalidate_q ;
  assign \u0.mmu_lsu_rd_w  = \fifo_d_rd.in ;
  assign \u0.mmu_lsu_req_tag_w  = 11'h000;
  assign \u0.mmu_lsu_resp_tag_w  = mem_d_resp_tag_i;
  assign \u0.mmu_lsu_wr_w  = \u0.u_lsu.mem_wr_o ;
  assign \u0.mmu_lsu_writeback_w  = \u0.u_lsu.mem_writeback_q ;
  assign \u0.mmu_mxr_w  = \u0.u_csr.u_csrfile.csr_sr_q [19];
  assign \u0.mmu_satp_w  = 32'h00000000;
  assign \u0.mmu_store_fault_w  = 1'h0;
  assign \u0.mmu_sum_w  = \u0.u_csr.u_csrfile.csr_sr_q [18];
  assign \u0.mul_hold_w  = \u0.u_exec.hold_i ;
  assign \u0.mul_opcode_invalid_w  = 1'h0;
  assign \u0.mul_opcode_opcode_w  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.mul_opcode_pc_w  = \u0.u_exec.opcode_pc_i ;
  assign \u0.mul_opcode_ra_idx_w  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.mul_opcode_ra_operand_w  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.mul_opcode_rb_idx_w  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.mul_opcode_rb_operand_w  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.mul_opcode_rd_idx_w  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.mul_opcode_valid_w  = \u0.u_div.opcode_valid_i ;
  assign \u0.opcode_invalid_w  = 1'h0;
  assign \u0.opcode_opcode_w  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.opcode_pc_w  = \u0.u_exec.opcode_pc_i ;
  assign \u0.opcode_ra_idx_w  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.opcode_ra_operand_w  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.opcode_rb_idx_w  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.opcode_rb_operand_w  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.opcode_rd_idx_w  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.reset_vector_i  = reset_vector_i;
  assign \u0.rst_i  = rst_i;
  assign \u0.squash_decode_w  = \u0.u_fetch.branch_request_i ;
  assign \u0.take_interrupt_w  = \u0.u_csr.take_interrupt_q ;
  assign \u0.u_csr.branch_csr_pc_o  = \u0.u_csr.branch_target_q ;
  assign \u0.u_csr.branch_csr_request_o  = \u0.u_csr.branch_q ;
  assign \u0.u_csr.clk_i  = clk_i;
  assign \u0.u_csr.cpu_id_i  = cpu_id_i;
  assign \u0.u_csr.csr_fault_r  = 1'h0;
  assign \u0.u_csr.csr_priv_r  = \u0.u_csr.opcode_opcode_i [29:28];
  assign \u0.u_csr.csr_result_e1_exception_o  = \u0.u_csr.exception_e1_q ;
  assign \u0.u_csr.csr_result_e1_value_o  = \u0.u_csr.rd_result_e1_q ;
  assign \u0.u_csr.csr_result_e1_wdata_o  = \u0.u_csr.csr_wdata_e1_q ;
  assign \u0.u_csr.csr_result_e1_write_o  = \u0.u_csr.rd_valid_e1_q ;
  assign \u0.u_csr.csr_writeback_exception_addr_i  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.u_csr.csr_writeback_exception_i  = \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.u_csr.csr_writeback_exception_pc_i  = \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  assign \u0.u_csr.csr_writeback_waddr_i  = \u0.u_issue.u_pipe_ctrl.opcode_wb_q [31:20];
  assign \u0.u_csr.csr_writeback_wdata_i  = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q ;
  assign \u0.u_csr.csr_writeback_write_i  = \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q ;
  assign \u0.u_csr.current_priv_w  = { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] };
  assign \u0.u_csr.ifence_o  = \u0.ifence_w ;
  assign \u0.u_csr.ifence_q  = \u0.ifence_w ;
  assign \u0.u_csr.intr_i  = intr_i;
  assign \u0.u_csr.misa_w  = 32'h40001100;
  assign \u0.u_csr.mmu_mxr_o  = \u0.u_csr.u_csrfile.csr_sr_q [19];
  assign \u0.u_csr.mmu_satp_o  = 32'h00000000;
  assign \u0.u_csr.mmu_sum_o  = \u0.u_csr.u_csrfile.csr_sr_q [18];
  assign \u0.u_csr.opcode_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_csr.opcode_ra_idx_i  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_csr.opcode_rb_idx_i  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_csr.opcode_rb_operand_i  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_csr.opcode_rd_idx_i  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_csr.reset_vector_i  = reset_vector_i;
  assign \u0.u_csr.rst_i  = rst_i;
  assign \u0.u_csr.satp_reg_w  = 32'h00000000;
  assign \u0.u_csr.status_reg_w  = \u0.u_csr.u_csrfile.csr_sr_q ;
  assign \u0.u_csr.take_interrupt_o  = \u0.u_csr.take_interrupt_q ;
  assign \u0.u_csr.timer_irq_w  = 1'h0;
  assign \u0.u_csr.u_csrfile.branch_r  = \u0.u_csr.csr_branch_w ;
  assign \u0.u_csr.u_csrfile.branch_target_r  = \u0.u_csr.csr_target_w ;
  assign \u0.u_csr.u_csrfile.clk_i  = clk_i;
  assign \u0.u_csr.u_csrfile.cpu_id_i  = cpu_id_i;
  assign \u0.u_csr.u_csrfile.csr_branch_o  = \u0.u_csr.csr_branch_w ;
  assign \u0.u_csr.u_csrfile.csr_mideleg_q  = 32'h00000000;
  assign { \u0.u_csr.u_csrfile.csr_mip_next_r [31:12], \u0.u_csr.u_csrfile.csr_mip_next_r [10:8], \u0.u_csr.u_csrfile.csr_mip_next_r [6:0] } = { \u0.u_csr.u_csrfile.csr_mip_next_q [31:12], \u0.u_csr.u_csrfile.csr_mip_next_q [10:8], \u0.u_csr.u_csrfile.csr_mip_next_q [6:0] };
  assign \u0.u_csr.u_csrfile.csr_mpriv_q [1] = \u0.u_csr.u_csrfile.csr_mpriv_q [0];
  assign \u0.u_csr.u_csrfile.csr_raddr_i  = \u0.u_csr.opcode_opcode_i [31:20];
  assign \u0.u_csr.u_csrfile.csr_rdata_o  = \u0.u_csr.csr_rdata_w ;
  assign \u0.u_csr.u_csrfile.csr_ren_i  = \u0.u_csr.opcode_valid_i ;
  assign \u0.u_csr.u_csrfile.csr_satp_q  = 32'h00000000;
  assign \u0.u_csr.u_csrfile.csr_sepc_q  = 32'h00000000;
  assign \u0.u_csr.u_csrfile.csr_stvec_q  = 32'h00000000;
  assign \u0.u_csr.u_csrfile.csr_target_o  = \u0.u_csr.csr_target_w ;
  assign \u0.u_csr.u_csrfile.csr_wdata_i  = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q ;
  assign \u0.u_csr.u_csrfile.exception_addr_i  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.u_csr.u_csrfile.exception_i  = \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.u_csr.u_csrfile.exception_pc_i  = \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  assign \u0.u_csr.u_csrfile.exception_s_w  = 1'h0;
  assign \u0.u_csr.u_csrfile.ext_intr_i  = intr_i;
  assign \u0.u_csr.u_csrfile.interrupt_o  = \u0.u_csr.interrupt_w ;
  assign \u0.u_csr.u_csrfile.irq_masked_r  = \u0.u_csr.interrupt_w ;
  assign \u0.u_csr.u_csrfile.irq_priv_r  = 2'h3;
  assign \u0.u_csr.u_csrfile.misa_i  = 32'h40001100;
  assign \u0.u_csr.u_csrfile.priv_o  = { \u0.u_csr.u_csrfile.csr_mpriv_q [0], \u0.u_csr.u_csrfile.csr_mpriv_q [0] };
  assign \u0.u_csr.u_csrfile.rdata_r  = \u0.u_csr.csr_rdata_w ;
  assign \u0.u_csr.u_csrfile.rst_i  = rst_i;
  assign \u0.u_csr.u_csrfile.satp_o  = 32'h00000000;
  assign \u0.u_csr.u_csrfile.status_o  = \u0.u_csr.u_csrfile.csr_sr_q ;
  assign \u0.u_csr.u_csrfile.timer_intr_i  = 1'h0;
  assign \u0.u_decode.clk_i  = clk_i;
  assign \u0.u_decode.enable_muldiv_w  = 1'h1;
  assign \u0.u_decode.fetch_in_accept_o  = \u0.u_fetch.fetch_accept_i ;
  assign \u0.u_decode.fetch_in_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_decode.fetch_in_valid_i  = \u0.u_decode.genblk1.u_dec.valid_i ;
  assign \u0.u_decode.fetch_out_accept_i  = \u0.u_fetch.fetch_accept_i ;
  assign \u0.u_decode.fetch_out_fault_fetch_o  = \u0.u_decode.fetch_in_fault_fetch_i ;
  assign \u0.u_decode.fetch_out_fault_page_o  = \u0.u_decode.fetch_in_fault_page_i ;
  assign \u0.u_decode.fetch_out_instr_branch_o  = \u0.u_decode.genblk1.u_dec.branch_o ;
  assign \u0.u_decode.fetch_out_instr_csr_o  = \u0.u_decode.genblk1.u_dec.csr_o ;
  assign \u0.u_decode.fetch_out_instr_div_o  = \u0.u_decode.genblk1.u_dec.div_o ;
  assign \u0.u_decode.fetch_out_instr_exec_o  = \u0.u_decode.genblk1.u_dec.exec_o ;
  assign \u0.u_decode.fetch_out_instr_invalid_o  = \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign \u0.u_decode.fetch_out_instr_lsu_o  = \u0.u_decode.genblk1.u_dec.lsu_o ;
  assign \u0.u_decode.fetch_out_instr_mul_o  = \u0.u_decode.genblk1.u_dec.mul_o ;
  assign \u0.u_decode.fetch_out_instr_o  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_decode.fetch_out_instr_rd_valid_o  = \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign \u0.u_decode.fetch_out_pc_o  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_decode.fetch_out_valid_o  = \u0.u_decode.genblk1.u_dec.valid_i ;
  assign \u0.u_decode.genblk1.fetch_in_instr_w  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_decode.genblk1.u_dec.enable_muldiv_i  = 1'h1;
  assign \u0.u_decode.genblk1.u_dec.invalid_o  = \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign \u0.u_decode.genblk1.u_dec.opcode_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_decode.rst_i  = rst_i;
  assign \u0.u_decode.squash_decode_i  = \u0.u_fetch.branch_request_i ;
  assign \u0.u_div.clk_i  = clk_i;
  assign \u0.u_div.opcode_invalid_i  = 1'h0;
  assign \u0.u_div.opcode_opcode_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_div.opcode_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_div.opcode_ra_idx_i  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_div.opcode_ra_operand_i  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_div.opcode_rb_idx_i  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_div.opcode_rd_idx_i  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_div.rst_i  = rst_i;
  assign \u0.u_div.writeback_valid_o  = \u0.u_div.valid_q ;
  assign \u0.u_div.writeback_value_o  = \u0.u_div.wb_result_q ;
  assign \u0.u_exec.bimm_r  = { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [7], \u0.u_csr.opcode_opcode_i [30:25], \u0.u_csr.opcode_opcode_i [11:8], 1'h0 };
  assign \u0.u_exec.branch_d_pc_o  = \u0.u_exec.branch_target_r ;
  assign \u0.u_exec.branch_d_priv_o  = 2'h0;
  assign \u0.u_exec.clk_i  = clk_i;
  assign \u0.u_exec.greater_than_signed$func$../../core/riscv/riscv_exec.v:362$760.v  = 32'hxxxxxxxx;
  assign \u0.u_exec.greater_than_signed$func$../../core/riscv/riscv_exec.v:362$760.x  = 32'hxxxxxxxx;
  assign \u0.u_exec.greater_than_signed$func$../../core/riscv/riscv_exec.v:362$760.y  = 32'hxxxxxxxx;
  assign \u0.u_exec.imm12_r  = { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31:20] };
  assign \u0.u_exec.imm20_r  = { \u0.u_csr.opcode_opcode_i [31:12], 12'h000 };
  assign \u0.u_exec.jimm20_r  = { \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [31], \u0.u_csr.opcode_opcode_i [19:12], \u0.u_csr.opcode_opcode_i [20], \u0.u_csr.opcode_opcode_i [30:21], 1'h0 };
  assign \u0.u_exec.less_than_signed$func$../../core/riscv/riscv_exec.v:357$759.v  = 32'hxxxxxxxx;
  assign \u0.u_exec.less_than_signed$func$../../core/riscv/riscv_exec.v:357$759.x  = 32'hxxxxxxxx;
  assign \u0.u_exec.less_than_signed$func$../../core/riscv/riscv_exec.v:357$759.y  = 32'hxxxxxxxx;
  assign \u0.u_exec.opcode_invalid_i  = 1'h0;
  assign \u0.u_exec.opcode_opcode_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_exec.opcode_ra_idx_i  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_exec.opcode_ra_operand_i  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_exec.opcode_rb_idx_i  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_exec.opcode_rb_operand_i  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_exec.opcode_rd_idx_i  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_exec.opcode_valid_i  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_exec.rst_i  = rst_i;
  assign \u0.u_exec.shamt_r  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_exec.u_alu.alu_a_i  = \u0.u_exec.alu_input_a_r ;
  assign \u0.u_exec.u_alu.alu_b_i  = \u0.u_exec.alu_input_b_r ;
  assign \u0.u_exec.u_alu.alu_op_i  = \u0.u_exec.alu_func_r ;
  assign \u0.u_exec.u_alu.alu_p_o  = \u0.u_exec.alu_p_w ;
  assign \u0.u_exec.u_alu.result_r  = \u0.u_exec.alu_p_w ;
  assign \u0.u_exec.writeback_value_o  = \u0.u_exec.result_q ;
  assign \u0.u_fetch.branch_pc_w  = \u0.u_fetch.branch_pc_q ;
  assign \u0.u_fetch.branch_w  = \u0.u_fetch.branch_q ;
  assign \u0.u_fetch.clk_i  = clk_i;
  assign \u0.u_fetch.fetch_fault_fetch_o  = \u0.u_decode.fetch_in_fault_fetch_i ;
  assign \u0.u_fetch.fetch_fault_page_o  = \u0.u_decode.fetch_in_fault_page_i ;
  assign \u0.u_fetch.fetch_instr_o  = \u0.u_decode.fetch_in_instr_i ;
  assign \u0.u_fetch.fetch_invalidate_i  = \u0.ifence_w ;
  assign \u0.u_fetch.fetch_pc_o  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_fetch.fetch_valid_o  = \u0.u_decode.genblk1.u_dec.valid_i ;
  assign \u0.u_fetch.icache_accept_i  = mem_i_accept_i;
  assign \u0.u_fetch.icache_error_i  = mem_i_error_i;
  assign \u0.u_fetch.icache_flush_o  = \u0.ifence_w ;
  assign \u0.u_fetch.icache_inst_i  = mem_i_inst_i;
  assign \u0.u_fetch.icache_invalidate_o  = 1'h0;
  assign \u0.u_fetch.icache_invalidate_q  = 1'h0;
  assign \u0.u_fetch.icache_page_fault_i  = 1'h0;
  assign \u0.u_fetch.icache_pc_o  = { \u0.u_fetch.pc_f_q [31:2], 2'h0 };
  assign \u0.u_fetch.icache_pc_w  = \u0.u_fetch.pc_f_q ;
  assign \u0.u_fetch.icache_rd_o  = \fifo_i_rd.in ;
  assign \u0.u_fetch.icache_valid_i  = mem_i_valid_i;
  assign \u0.u_fetch.rst_i  = rst_i;
  assign \u0.u_fetch.squash_decode_o  = \u0.u_fetch.branch_request_i ;
  assign \u0.u_issue.branch_csr_pc_i  = \u0.u_csr.branch_target_q ;
  assign \u0.u_issue.branch_csr_request_i  = \u0.u_csr.branch_q ;
  assign \u0.u_issue.branch_d_exec_pc_i  = \u0.u_exec.branch_target_r ;
  assign \u0.u_issue.branch_d_exec_priv_i  = 2'h0;
  assign \u0.u_issue.branch_d_exec_request_i  = \u0.u_exec.branch_d_request_o ;
  assign \u0.u_issue.branch_pc_o  = \u0.u_fetch.branch_pc_i ;
  assign \u0.u_issue.branch_request_o  = \u0.u_fetch.branch_request_i ;
  assign \u0.u_issue.clk_i  = clk_i;
  assign \u0.u_issue.csr_opcode_invalid_o  = \u0.u_csr.opcode_invalid_i ;
  assign \u0.u_issue.csr_opcode_opcode_o  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_issue.csr_opcode_pc_o  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_issue.csr_opcode_ra_idx_o  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_issue.csr_opcode_ra_operand_o  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_issue.csr_opcode_rb_idx_o  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_issue.csr_opcode_rb_operand_o  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_issue.csr_opcode_rd_idx_o  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_issue.csr_opcode_valid_o  = \u0.u_csr.opcode_valid_i ;
  assign \u0.u_issue.csr_result_e1_exception_i  = \u0.u_csr.exception_e1_q ;
  assign \u0.u_issue.csr_result_e1_value_i  = \u0.u_csr.rd_result_e1_q ;
  assign \u0.u_issue.csr_result_e1_wdata_i  = \u0.u_csr.csr_wdata_e1_q ;
  assign \u0.u_issue.csr_result_e1_write_i  = \u0.u_csr.rd_valid_e1_q ;
  assign \u0.u_issue.csr_writeback_exception_addr_o  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.u_issue.csr_writeback_exception_o  = \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.u_issue.csr_writeback_exception_pc_o  = \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  assign \u0.u_issue.csr_writeback_waddr_o  = \u0.u_issue.u_pipe_ctrl.opcode_wb_q [31:20];
  assign \u0.u_issue.csr_writeback_wdata_o  = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q ;
  assign \u0.u_issue.csr_writeback_write_o  = \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q ;
  assign \u0.u_issue.div_opcode_valid_o  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.enable_mul_bypass_w  = 1'h1;
  assign \u0.u_issue.enable_muldiv_w  = 1'h1;
  assign \u0.u_issue.exec_hold_o  = \u0.u_exec.hold_i ;
  assign \u0.u_issue.exec_opcode_valid_o  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.fetch_accept_o  = \u0.u_fetch.fetch_accept_i ;
  assign \u0.u_issue.fetch_fault_fetch_i  = \u0.u_decode.fetch_in_fault_fetch_i ;
  assign \u0.u_issue.fetch_fault_page_i  = \u0.u_decode.fetch_in_fault_page_i ;
  assign \u0.u_issue.fetch_instr_branch_i  = \u0.u_decode.genblk1.u_dec.branch_o ;
  assign \u0.u_issue.fetch_instr_csr_i  = \u0.u_decode.genblk1.u_dec.csr_o ;
  assign \u0.u_issue.fetch_instr_div_i  = \u0.u_decode.genblk1.u_dec.div_o ;
  assign \u0.u_issue.fetch_instr_exec_i  = \u0.u_decode.genblk1.u_dec.exec_o ;
  assign \u0.u_issue.fetch_instr_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_issue.fetch_instr_invalid_i  = \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign \u0.u_issue.fetch_instr_lsu_i  = \u0.u_decode.genblk1.u_dec.lsu_o ;
  assign \u0.u_issue.fetch_instr_mul_i  = \u0.u_decode.genblk1.u_dec.mul_o ;
  assign \u0.u_issue.fetch_instr_rd_valid_i  = \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign \u0.u_issue.fetch_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_issue.fetch_valid_i  = \u0.u_decode.genblk1.u_dec.valid_i ;
  assign \u0.u_issue.interrupt_inhibit_o  = \u0.u_csr.interrupt_inhibit_i ;
  assign \u0.u_issue.issue_branch_w  = \u0.u_decode.genblk1.u_dec.branch_o ;
  assign \u0.u_issue.issue_csr_w  = \u0.u_decode.genblk1.u_dec.csr_o ;
  assign \u0.u_issue.issue_div_w  = \u0.u_decode.genblk1.u_dec.div_o ;
  assign \u0.u_issue.issue_exec_w  = \u0.u_decode.genblk1.u_dec.exec_o ;
  assign \u0.u_issue.issue_invalid_w  = \u0.u_decode.genblk1.u_dec.invalid_w ;
  assign \u0.u_issue.issue_lsu_w  = \u0.u_decode.genblk1.u_dec.lsu_o ;
  assign \u0.u_issue.issue_mul_w  = \u0.u_decode.genblk1.u_dec.mul_o ;
  assign \u0.u_issue.issue_ra_idx_w  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_issue.issue_ra_value_r  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_issue.issue_rb_idx_w  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_issue.issue_rb_value_r  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_issue.issue_rd_idx_w  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_issue.issue_sb_alloc_w  = \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign \u0.u_issue.lsu_opcode_invalid_o  = 1'h0;
  assign \u0.u_issue.lsu_opcode_opcode_o  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_issue.lsu_opcode_pc_o  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_issue.lsu_opcode_ra_idx_o  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_issue.lsu_opcode_ra_operand_o  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_issue.lsu_opcode_rb_idx_o  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_issue.lsu_opcode_rb_operand_o  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_issue.lsu_opcode_rd_idx_o  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_issue.lsu_opcode_valid_o  = \u0.u_csr.opcode_valid_i ;
  assign \u0.u_issue.mul_hold_o  = \u0.u_exec.hold_i ;
  assign \u0.u_issue.mul_opcode_invalid_o  = 1'h0;
  assign \u0.u_issue.mul_opcode_opcode_o  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_issue.mul_opcode_pc_o  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_issue.mul_opcode_ra_idx_o  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_issue.mul_opcode_ra_operand_o  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_issue.mul_opcode_rb_idx_o  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_issue.mul_opcode_rb_operand_o  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_issue.mul_opcode_rd_idx_o  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_issue.mul_opcode_valid_o  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.opcode_accept_r  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.opcode_invalid_o  = 1'h0;
  assign \u0.u_issue.opcode_issue_r  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.opcode_opcode_o  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_issue.opcode_pc_o  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_issue.opcode_ra_idx_o  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_issue.opcode_ra_operand_o  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_issue.opcode_rb_idx_o  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_issue.opcode_rb_operand_o  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_issue.opcode_rd_idx_o  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_issue.pipe_branch_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [6];
  assign \u0.u_issue.pipe_exception_wb_w  = \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.u_issue.pipe_load_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [1];
  assign \u0.u_issue.pipe_load_e2_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [1];
  assign \u0.u_issue.pipe_mul_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [5];
  assign \u0.u_issue.pipe_mul_e2_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [5];
  assign \u0.u_issue.pipe_opc_wb_w  = \u0.u_issue.u_pipe_ctrl.opcode_wb_q ;
  assign \u0.u_issue.pipe_opcode_e1_w  = \u0.u_issue.u_pipe_ctrl.opcode_e1_q ;
  assign \u0.u_issue.pipe_pc_e1_w  = \u0.u_issue.u_pipe_ctrl.pc_e1_q ;
  assign \u0.u_issue.pipe_pc_wb_w  = \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  assign \u0.u_issue.pipe_result_wb_w  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.u_issue.pipe_stall_raw_w  = \u0.u_exec.hold_i ;
  assign \u0.u_issue.pipe_store_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [2];
  assign \u0.u_issue.pipe_valid_wb_w  = \u0.u_issue.u_pipe_ctrl.valid_wb_o ;
  assign \u0.u_issue.rst_i  = rst_i;
  assign \u0.u_issue.squash_w  = \u0.u_issue.pipe_squash_e1_e2_w ;
  assign \u0.u_issue.stall_w  = \u0.u_exec.hold_i ;
  assign \u0.u_issue.take_interrupt_i  = \u0.u_csr.take_interrupt_q ;
  assign \u0.u_issue.u_pipe_ctrl.alu_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [0];
  assign \u0.u_issue.u_pipe_ctrl.alu_result_e1_i  = \u0.u_exec.result_q ;
  assign \u0.u_issue.u_pipe_ctrl.branch_e1_o  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [6];
  assign \u0.u_issue.u_pipe_ctrl.clk_i  = clk_i;
  assign \u0.u_issue.u_pipe_ctrl.csr_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [3];
  assign \u0.u_issue.u_pipe_ctrl.csr_result_exception_e1_i  = \u0.u_csr.exception_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.csr_result_value_e1_i  = \u0.u_csr.rd_result_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.csr_result_wdata_e1_i  = \u0.u_csr.csr_wdata_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.csr_result_write_e1_i  = \u0.u_csr.rd_valid_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.csr_waddr_wb_o  = \u0.u_issue.u_pipe_ctrl.opcode_wb_q [31:20];
  assign \u0.u_issue.u_pipe_ctrl.csr_wb_o  = \u0.u_issue.pipe_csr_wb_w ;
  assign \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_o  = \u0.u_issue.u_pipe_ctrl.csr_wdata_wb_q ;
  assign \u0.u_issue.u_pipe_ctrl.csr_write_wb_o  = \u0.u_issue.u_pipe_ctrl.csr_wr_wb_q ;
  assign \u0.u_issue.u_pipe_ctrl.div_complete_i  = \u0.u_div.valid_q ;
  assign \u0.u_issue.u_pipe_ctrl.div_e1_w  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [4];
  assign \u0.u_issue.u_pipe_ctrl.div_result_i  = \u0.u_div.wb_result_q ;
  assign \u0.u_issue.u_pipe_ctrl.exception_wb_o  = \u0.u_issue.u_pipe_ctrl.exception_wb_q ;
  assign \u0.u_issue.u_pipe_ctrl.issue_accept_i  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.u_pipe_ctrl.issue_branch_i  = \u0.u_decode.genblk1.u_dec.branch_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_branch_taken_i  = \u0.u_exec.branch_d_request_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_branch_target_i  = \u0.u_exec.branch_target_r ;
  assign \u0.u_issue.u_pipe_ctrl.issue_csr_i  = \u0.u_decode.genblk1.u_dec.csr_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_div_i  = \u0.u_decode.genblk1.u_dec.div_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_exception_i  = { 1'h0, \u0.u_issue.issue_fault_w  };
  assign \u0.u_issue.u_pipe_ctrl.issue_lsu_i  = \u0.u_decode.genblk1.u_dec.lsu_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_mul_i  = \u0.u_decode.genblk1.u_dec.mul_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_opcode_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_issue.u_pipe_ctrl.issue_operand_ra_i  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_issue.u_pipe_ctrl.issue_operand_rb_i  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_issue.u_pipe_ctrl.issue_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_issue.u_pipe_ctrl.issue_rd_i  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_issue.u_pipe_ctrl.issue_rd_valid_i  = \u0.u_decode.genblk1.u_dec.rd_valid_o ;
  assign \u0.u_issue.u_pipe_ctrl.issue_stall_i  = \u0.u_exec.hold_i ;
  assign \u0.u_issue.u_pipe_ctrl.issue_valid_i  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_issue.u_pipe_ctrl.load_e1_o  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [1];
  assign \u0.u_issue.u_pipe_ctrl.load_e2_o  = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [1];
  assign \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i [5] = 1'h0;
  assign \u0.u_issue.u_pipe_ctrl.mul_e1_o  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [5];
  assign \u0.u_issue.u_pipe_ctrl.mul_e2_o  = \u0.u_issue.u_pipe_ctrl.ctrl_e2_q [5];
  assign \u0.u_issue.u_pipe_ctrl.mul_result_e2_i  = \u0.u_mul.result_e2_q ;
  assign \u0.u_issue.u_pipe_ctrl.opcode_e1_o  = \u0.u_issue.u_pipe_ctrl.opcode_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.opcode_wb_o  = \u0.u_issue.u_pipe_ctrl.opcode_wb_q ;
  assign \u0.u_issue.u_pipe_ctrl.pc_e1_o  = \u0.u_issue.u_pipe_ctrl.pc_e1_q ;
  assign \u0.u_issue.u_pipe_ctrl.pc_wb_o  = \u0.u_issue.u_pipe_ctrl.pc_wb_q ;
  assign \u0.u_issue.u_pipe_ctrl.rd_e1_o  = \u0.u_issue.pipe_rd_e1_w ;
  assign \u0.u_issue.u_pipe_ctrl.rd_e2_o  = \u0.u_issue.pipe_rd_e2_w ;
  assign \u0.u_issue.u_pipe_ctrl.rd_wb_o  = \u0.u_issue.pipe_rd_wb_w ;
  assign \u0.u_issue.u_pipe_ctrl.result_e2_o  = \u0.u_issue.pipe_result_e2_w ;
  assign \u0.u_issue.u_pipe_ctrl.result_e2_r  = \u0.u_issue.pipe_result_e2_w ;
  assign \u0.u_issue.u_pipe_ctrl.result_wb_o  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.u_issue.u_pipe_ctrl.rst_i  = rst_i;
  assign \u0.u_issue.u_pipe_ctrl.squash_e1_e2_i  = 1'h0;
  assign \u0.u_issue.u_pipe_ctrl.squash_e1_e2_o  = \u0.u_issue.pipe_squash_e1_e2_w ;
  assign \u0.u_issue.u_pipe_ctrl.squash_wb_i  = 1'h0;
  assign \u0.u_issue.u_pipe_ctrl.stall_o  = \u0.u_exec.hold_i ;
  assign \u0.u_issue.u_pipe_ctrl.store_e1_o  = \u0.u_issue.u_pipe_ctrl.ctrl_e1_q [2];
  assign \u0.u_issue.u_pipe_ctrl.take_interrupt_i  = \u0.u_csr.take_interrupt_q ;
  assign \u0.u_issue.u_regfile.REGFILE.ra0_value_r  = \u0.u_issue.issue_ra_value_w ;
  assign \u0.u_issue.u_regfile.REGFILE.rb0_value_r  = \u0.u_issue.issue_rb_value_w ;
  assign \u0.u_issue.u_regfile.REGFILE.x0_zero_w  = 32'h00000000;
  assign \u0.u_issue.u_regfile.REGFILE.x10_a0_w  = \u0.u_issue.u_regfile.REGFILE.reg_r10_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x11_a1_w  = \u0.u_issue.u_regfile.REGFILE.reg_r11_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x12_a2_w  = \u0.u_issue.u_regfile.REGFILE.reg_r12_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x13_a3_w  = \u0.u_issue.u_regfile.REGFILE.reg_r13_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x14_a4_w  = \u0.u_issue.u_regfile.REGFILE.reg_r14_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x15_a5_w  = \u0.u_issue.u_regfile.REGFILE.reg_r15_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x16_a6_w  = \u0.u_issue.u_regfile.REGFILE.reg_r16_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x17_a7_w  = \u0.u_issue.u_regfile.REGFILE.reg_r17_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x18_s2_w  = \u0.u_issue.u_regfile.REGFILE.reg_r18_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x19_s3_w  = \u0.u_issue.u_regfile.REGFILE.reg_r19_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x1_ra_w  = \u0.u_issue.u_regfile.REGFILE.reg_r1_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x20_s4_w  = \u0.u_issue.u_regfile.REGFILE.reg_r20_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x21_s5_w  = \u0.u_issue.u_regfile.REGFILE.reg_r21_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x22_s6_w  = \u0.u_issue.u_regfile.REGFILE.reg_r22_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x23_s7_w  = \u0.u_issue.u_regfile.REGFILE.reg_r23_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x24_s8_w  = \u0.u_issue.u_regfile.REGFILE.reg_r24_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x25_s9_w  = \u0.u_issue.u_regfile.REGFILE.reg_r25_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x26_s10_w  = \u0.u_issue.u_regfile.REGFILE.reg_r26_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x27_s11_w  = \u0.u_issue.u_regfile.REGFILE.reg_r27_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x28_t3_w  = \u0.u_issue.u_regfile.REGFILE.reg_r28_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x29_t4_w  = \u0.u_issue.u_regfile.REGFILE.reg_r29_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x2_sp_w  = \u0.u_issue.u_regfile.REGFILE.reg_r2_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x30_t5_w  = \u0.u_issue.u_regfile.REGFILE.reg_r30_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x31_t6_w  = \u0.u_issue.u_regfile.REGFILE.reg_r31_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x3_gp_w  = \u0.u_issue.u_regfile.REGFILE.reg_r3_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x4_tp_w  = \u0.u_issue.u_regfile.REGFILE.reg_r4_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x5_t0_w  = \u0.u_issue.u_regfile.REGFILE.reg_r5_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x6_t1_w  = \u0.u_issue.u_regfile.REGFILE.reg_r6_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x7_t2_w  = \u0.u_issue.u_regfile.REGFILE.reg_r7_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x8_s0_w  = \u0.u_issue.u_regfile.REGFILE.reg_r8_q ;
  assign \u0.u_issue.u_regfile.REGFILE.x9_s1_w  = \u0.u_issue.u_regfile.REGFILE.reg_r9_q ;
  assign \u0.u_issue.u_regfile.clk_i  = clk_i;
  assign \u0.u_issue.u_regfile.ra0_i  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_issue.u_regfile.ra0_value_o  = \u0.u_issue.issue_ra_value_w ;
  assign \u0.u_issue.u_regfile.rb0_i  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_issue.u_regfile.rb0_value_o  = \u0.u_issue.issue_rb_value_w ;
  assign \u0.u_issue.u_regfile.rd0_i  = \u0.u_issue.pipe_rd_wb_w ;
  assign \u0.u_issue.u_regfile.rd0_value_i  = \u0.u_issue.u_pipe_ctrl.result_wb_q ;
  assign \u0.u_issue.u_regfile.rst_i  = rst_i;
  assign \u0.u_issue.writeback_div_valid_i  = \u0.u_div.valid_q ;
  assign \u0.u_issue.writeback_div_value_i  = \u0.u_div.wb_result_q ;
  assign \u0.u_issue.writeback_exec_value_i  = \u0.u_exec.result_q ;
  assign \u0.u_issue.writeback_mem_exception_i  = { 1'h0, \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i [4:0] };
  assign \u0.u_issue.writeback_mem_valid_i  = \u0.u_issue.u_pipe_ctrl.mem_complete_i ;
  assign \u0.u_issue.writeback_mem_value_i  = \u0.u_issue.u_pipe_ctrl.mem_result_e2_i ;
  assign \u0.u_issue.writeback_mul_value_i  = \u0.u_mul.result_e2_q ;
  assign \u0.u_lsu.addr_lsb_r  = \u0.u_lsu.u_lsu_request.data_out_o [5:4];
  assign \u0.u_lsu.clk_i  = clk_i;
  assign \u0.u_lsu.load_byte_r  = \u0.u_lsu.u_lsu_request.data_out_o [1];
  assign \u0.u_lsu.load_half_r  = \u0.u_lsu.u_lsu_request.data_out_o [2];
  assign \u0.u_lsu.load_signed_r  = \u0.u_lsu.u_lsu_request.data_out_o [3];
  assign \u0.u_lsu.mem_accept_i  = mem_d_accept_i;
  assign \u0.u_lsu.mem_ack_i  = mem_d_ack_i;
  assign \u0.u_lsu.mem_addr_o  = { \u0.u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u0.u_lsu.mem_cacheable_o  = \u0.mem_d_cacheable_o ;
  assign \u0.u_lsu.mem_cacheable_q  = \u0.mem_d_cacheable_o ;
  assign \u0.u_lsu.mem_data_rd_i  = mem_d_data_rd_i;
  assign \u0.u_lsu.mem_data_wr_o  = \u0.u_lsu.mem_data_wr_q ;
  assign \u0.u_lsu.mem_error_i  = mem_d_error_i;
  assign \u0.u_lsu.mem_flush_o  = \u0.u_lsu.mem_flush_q ;
  assign \u0.u_lsu.mem_invalidate_o  = \u0.u_lsu.mem_invalidate_q ;
  assign \u0.u_lsu.mem_load_fault_i  = 1'h0;
  assign \u0.u_lsu.mem_rd_o  = \fifo_d_rd.in ;
  assign \u0.u_lsu.mem_req_tag_o  = 11'h000;
  assign \u0.u_lsu.mem_resp_tag_i  = mem_d_resp_tag_i;
  assign \u0.u_lsu.mem_store_fault_i  = 1'h0;
  assign \u0.u_lsu.mem_writeback_o  = \u0.u_lsu.mem_writeback_q ;
  assign \u0.u_lsu.opcode_invalid_i  = 1'h0;
  assign \u0.u_lsu.opcode_opcode_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_lsu.opcode_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_lsu.opcode_ra_idx_i  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_lsu.opcode_ra_operand_i  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_lsu.opcode_rb_idx_i  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_lsu.opcode_rb_operand_i  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_lsu.opcode_rd_idx_i  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_lsu.opcode_valid_i  = \u0.u_csr.opcode_valid_i ;
  assign \u0.u_lsu.resp_addr_w  = \u0.u_lsu.u_lsu_request.data_out_o [35:4];
  assign \u0.u_lsu.resp_byte_w  = \u0.u_lsu.u_lsu_request.data_out_o [1];
  assign \u0.u_lsu.resp_half_w  = \u0.u_lsu.u_lsu_request.data_out_o [2];
  assign \u0.u_lsu.resp_load_w  = \u0.u_lsu.u_lsu_request.data_out_o [0];
  assign \u0.u_lsu.resp_signed_w  = \u0.u_lsu.u_lsu_request.data_out_o [3];
  assign \u0.u_lsu.rst_i  = rst_i;
  assign \u0.u_lsu.stall_o  = \u0.u_issue.lsu_stall_i ;
  assign \u0.u_lsu.u_lsu_request.clk_i  = clk_i;
  assign \u0.u_lsu.u_lsu_request.data_in_i  = { \u0.u_lsu.mem_addr_q , \u0.u_lsu.mem_ls_q , \u0.u_lsu.mem_xh_q , \u0.u_lsu.mem_xb_q , \u0.u_lsu.mem_load_q  };
  assign \u0.u_lsu.u_lsu_request.rst_i  = rst_i;
  assign \u0.u_lsu.wb_result_r  = \u0.u_issue.u_pipe_ctrl.mem_result_e2_i ;
  assign \u0.u_lsu.writeback_exception_o  = { 1'h0, \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i [4:0] };
  assign \u0.u_lsu.writeback_valid_o  = \u0.u_issue.u_pipe_ctrl.mem_complete_i ;
  assign \u0.u_lsu.writeback_value_o  = \u0.u_issue.u_pipe_ctrl.mem_result_e2_i ;
  assign \u0.u_mmu.clk_i  = clk_i;
  assign \u0.u_mmu.fetch_in_accept_o  = mem_i_accept_i;
  assign \u0.u_mmu.fetch_in_error_o  = mem_i_error_i;
  assign \u0.u_mmu.fetch_in_fault_o  = 1'h0;
  assign \u0.u_mmu.fetch_in_flush_i  = \u0.ifence_w ;
  assign \u0.u_mmu.fetch_in_inst_o  = mem_i_inst_i;
  assign \u0.u_mmu.fetch_in_invalidate_i  = 1'h0;
  assign \u0.u_mmu.fetch_in_pc_i  = { \u0.u_fetch.pc_f_q [31:2], 2'h0 };
  assign \u0.u_mmu.fetch_in_rd_i  = \fifo_i_rd.in ;
  assign \u0.u_mmu.fetch_in_valid_o  = mem_i_valid_i;
  assign \u0.u_mmu.fetch_out_accept_i  = mem_i_accept_i;
  assign \u0.u_mmu.fetch_out_error_i  = mem_i_error_i;
  assign \u0.u_mmu.fetch_out_flush_o  = \u0.ifence_w ;
  assign \u0.u_mmu.fetch_out_inst_i  = mem_i_inst_i;
  assign \u0.u_mmu.fetch_out_invalidate_o  = 1'h0;
  assign \u0.u_mmu.fetch_out_pc_o  = { \u0.u_fetch.pc_f_q [31:2], 2'h0 };
  assign \u0.u_mmu.fetch_out_rd_o  = \fifo_i_rd.in ;
  assign \u0.u_mmu.fetch_out_valid_i  = mem_i_valid_i;
  assign \u0.u_mmu.lsu_in_accept_o  = mem_d_accept_i;
  assign \u0.u_mmu.lsu_in_ack_o  = mem_d_ack_i;
  assign \u0.u_mmu.lsu_in_addr_i  = { \u0.u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u0.u_mmu.lsu_in_cacheable_i  = \u0.mem_d_cacheable_o ;
  assign \u0.u_mmu.lsu_in_data_rd_o  = mem_d_data_rd_i;
  assign \u0.u_mmu.lsu_in_data_wr_i  = \u0.u_lsu.mem_data_wr_q ;
  assign \u0.u_mmu.lsu_in_error_o  = mem_d_error_i;
  assign \u0.u_mmu.lsu_in_flush_i  = \u0.u_lsu.mem_flush_q ;
  assign \u0.u_mmu.lsu_in_invalidate_i  = \u0.u_lsu.mem_invalidate_q ;
  assign \u0.u_mmu.lsu_in_load_fault_o  = 1'h0;
  assign \u0.u_mmu.lsu_in_rd_i  = \fifo_d_rd.in ;
  assign \u0.u_mmu.lsu_in_req_tag_i  = 11'h000;
  assign \u0.u_mmu.lsu_in_resp_tag_o  = mem_d_resp_tag_i;
  assign \u0.u_mmu.lsu_in_store_fault_o  = 1'h0;
  assign \u0.u_mmu.lsu_in_wr_i  = \u0.u_lsu.mem_wr_o ;
  assign \u0.u_mmu.lsu_in_writeback_i  = \u0.u_lsu.mem_writeback_q ;
  assign \u0.u_mmu.lsu_out_accept_i  = mem_d_accept_i;
  assign \u0.u_mmu.lsu_out_ack_i  = mem_d_ack_i;
  assign \u0.u_mmu.lsu_out_addr_o  = { \u0.u_lsu.mem_addr_q [31:2], 2'h0 };
  assign \u0.u_mmu.lsu_out_cacheable_o  = \u0.mem_d_cacheable_o ;
  assign \u0.u_mmu.lsu_out_data_rd_i  = mem_d_data_rd_i;
  assign \u0.u_mmu.lsu_out_data_wr_o  = \u0.u_lsu.mem_data_wr_q ;
  assign \u0.u_mmu.lsu_out_error_i  = mem_d_error_i;
  assign \u0.u_mmu.lsu_out_flush_o  = \u0.u_lsu.mem_flush_q ;
  assign \u0.u_mmu.lsu_out_invalidate_o  = \u0.u_lsu.mem_invalidate_q ;
  assign \u0.u_mmu.lsu_out_rd_o  = \fifo_d_rd.in ;
  assign \u0.u_mmu.lsu_out_req_tag_o  = 11'h000;
  assign \u0.u_mmu.lsu_out_resp_tag_i  = mem_d_resp_tag_i;
  assign \u0.u_mmu.lsu_out_wr_o  = \u0.u_lsu.mem_wr_o ;
  assign \u0.u_mmu.lsu_out_writeback_o  = \u0.u_lsu.mem_writeback_q ;
  assign \u0.u_mmu.mxr_i  = \u0.u_csr.u_csrfile.csr_sr_q [19];
  assign \u0.u_mmu.rst_i  = rst_i;
  assign \u0.u_mmu.satp_i  = 32'h00000000;
  assign \u0.u_mmu.sum_i  = \u0.u_csr.u_csrfile.csr_sr_q [18];
  assign \u0.u_mul.clk_i  = clk_i;
  assign \u0.u_mul.hold_i  = \u0.u_exec.hold_i ;
  assign \u0.u_mul.opcode_invalid_i  = 1'h0;
  assign \u0.u_mul.opcode_opcode_i  = \u0.u_csr.opcode_opcode_i ;
  assign \u0.u_mul.opcode_pc_i  = \u0.u_exec.opcode_pc_i ;
  assign \u0.u_mul.opcode_ra_idx_i  = \u0.u_csr.opcode_opcode_i [19:15];
  assign \u0.u_mul.opcode_ra_operand_i  = \u0.u_csr.opcode_ra_operand_i ;
  assign \u0.u_mul.opcode_rb_idx_i  = \u0.u_csr.opcode_opcode_i [24:20];
  assign \u0.u_mul.opcode_rb_operand_i  = \u0.u_div.opcode_rb_operand_i ;
  assign \u0.u_mul.opcode_rd_idx_i  = \u0.u_csr.opcode_opcode_i [11:7];
  assign \u0.u_mul.opcode_valid_i  = \u0.u_div.opcode_valid_i ;
  assign \u0.u_mul.rst_i  = rst_i;
  assign \u0.u_mul.writeback_value_o  = \u0.u_mul.result_e2_q ;
  assign \u0.writeback_div_valid_w  = \u0.u_div.valid_q ;
  assign \u0.writeback_div_value_w  = \u0.u_div.wb_result_q ;
  assign \u0.writeback_exec_value_w  = \u0.u_exec.result_q ;
  assign \u0.writeback_mem_exception_w  = { 1'h0, \u0.u_issue.u_pipe_ctrl.mem_exception_e2_i [4:0] };
  assign \u0.writeback_mem_valid_w  = \u0.u_issue.u_pipe_ctrl.mem_complete_i ;
  assign \u0.writeback_mem_value_w  = \u0.u_issue.u_pipe_ctrl.mem_result_e2_i ;
  assign \u0.writeback_mul_value_w  = \u0.u_mul.result_e2_q ;
  assign wr_d_addr = \fifo_d_addr.wr ;
  assign wr_d_data_wr = \u0.u_lsu.mem_wr_o [0];
  assign wr_d_rd = \fifo_d_rd.in ;
  assign wr_i_rd = \fifo_i_rd.in ;
  assign wri_rd = \fifo_i_pc.wr ;
endmodule
