module SDP_Y_CVT_chn_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_cvt.v:268" *)
  input in_0;
  (* src = "./vmod/nvdla/sdp/NV_NVDLA_SDP_CORE_Y_cvt.v:269" *)
  output outsig;
  assign outsig = in_0;
endmodule
