module FP17_TO_FP16_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:248" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_to_fp16.v:249" *)
  output outsig;
  assign outsig = in_0;
endmodule
