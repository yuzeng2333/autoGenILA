module S(clk, in, out);
  logic [7:0] _000_;
  logic _001_;
  logic _002_;
  logic _003_;
  logic _004_;
  logic _005_;
  logic _006_;
  logic _007_;
  logic _008_;
  logic _009_;
  logic _010_;
  logic _011_;
  logic _012_;
  logic _013_;
  logic _014_;
  logic _015_;
  logic _016_;
  logic _017_;
  logic _018_;
  logic _019_;
  logic _020_;
  logic _021_;
  logic _022_;
  logic _023_;
  logic _024_;
  logic _025_;
  logic _026_;
  logic _027_;
  logic _028_;
  logic _029_;
  logic _030_;
  logic _031_;
  logic _032_;
  logic _033_;
  logic _034_;
  logic _035_;
  logic _036_;
  logic _037_;
  logic _038_;
  logic _039_;
  logic _040_;
  logic _041_;
  logic _042_;
  logic _043_;
  logic _044_;
  logic _045_;
  logic _046_;
  logic _047_;
  logic _048_;
  logic _049_;
  logic _050_;
  logic _051_;
  logic _052_;
  logic _053_;
  logic _054_;
  logic _055_;
  logic _056_;
  logic _057_;
  logic _058_;
  logic _059_;
  logic _060_;
  logic _061_;
  logic _062_;
  logic _063_;
  logic _064_;
  logic _065_;
  logic _066_;
  logic _067_;
  logic _068_;
  logic _069_;
  logic _070_;
  logic _071_;
  logic _072_;
  logic _073_;
  logic _074_;
  logic _075_;
  logic _076_;
  logic _077_;
  logic _078_;
  logic _079_;
  logic _080_;
  logic _081_;
  logic _082_;
  logic _083_;
  logic _084_;
  logic _085_;
  logic _086_;
  logic _087_;
  logic _088_;
  logic _089_;
  logic _090_;
  logic _091_;
  logic _092_;
  logic _093_;
  logic _094_;
  logic _095_;
  logic _096_;
  logic _097_;
  logic _098_;
  logic _099_;
  logic _100_;
  logic _101_;
  logic _102_;
  logic _103_;
  logic _104_;
  logic _105_;
  logic _106_;
  logic _107_;
  logic _108_;
  logic _109_;
  logic _110_;
  logic _111_;
  logic _112_;
  logic _113_;
  logic _114_;
  logic _115_;
  logic _116_;
  logic _117_;
  logic _118_;
  logic _119_;
  logic _120_;
  logic _121_;
  logic _122_;
  logic _123_;
  logic _124_;
  logic _125_;
  logic _126_;
  logic _127_;
  logic _128_;
  logic _129_;
  logic _130_;
  logic _131_;
  logic _132_;
  logic _133_;
  logic _134_;
  logic _135_;
  logic _136_;
  logic _137_;
  logic _138_;
  logic _139_;
  logic _140_;
  logic _141_;
  logic _142_;
  logic _143_;
  logic _144_;
  logic _145_;
  logic _146_;
  logic _147_;
  logic _148_;
  logic _149_;
  logic _150_;
  logic _151_;
  logic _152_;
  logic _153_;
  logic _154_;
  logic _155_;
  logic _156_;
  logic _157_;
  logic _158_;
  logic _159_;
  logic _160_;
  logic _161_;
  logic _162_;
  logic _163_;
  logic _164_;
  logic _165_;
  logic _166_;
  logic _167_;
  logic _168_;
  logic _169_;
  logic _170_;
  logic _171_;
  logic _172_;
  logic _173_;
  logic _174_;
  logic _175_;
  logic _176_;
  logic _177_;
  logic _178_;
  logic _179_;
  logic _180_;
  logic _181_;
  logic _182_;
  logic _183_;
  logic _184_;
  logic _185_;
  logic _186_;
  logic _187_;
  logic _188_;
  logic _189_;
  logic _190_;
  logic _191_;
  logic _192_;
  logic _193_;
  logic _194_;
  logic _195_;
  logic _196_;
  logic _197_;
  logic _198_;
  logic _199_;
  logic _200_;
  logic _201_;
  logic _202_;
  logic _203_;
  logic _204_;
  logic _205_;
  logic _206_;
  logic _207_;
  logic _208_;
  logic _209_;
  logic _210_;
  logic _211_;
  logic _212_;
  logic _213_;
  logic _214_;
  logic _215_;
  logic _216_;
  logic _217_;
  logic _218_;
  logic _219_;
  logic _220_;
  logic _221_;
  logic _222_;
  logic _223_;
  logic _224_;
  logic _225_;
  logic _226_;
  logic _227_;
  logic _228_;
  logic _229_;
  logic _230_;
  logic _231_;
  logic _232_;
  logic _233_;
  logic _234_;
  logic _235_;
  logic _236_;
  logic _237_;
  logic _238_;
  logic _239_;
  logic _240_;
  logic _241_;
  logic _242_;
  logic _243_;
  logic _244_;
  logic _245_;
  logic _246_;
  logic _247_;
  logic _248_;
  logic _249_;
  logic _250_;
  logic _251_;
  logic _252_;
  logic _253_;
  logic _254_;
  logic _255_;
  logic _256_;
  input clk;
  input [7:0] in;
  output [7:0] out;
  logic [7:0] out;
  always @(posedge clk)
      out <= _000_;
  assign _001_ = in == 8'h9e;
  assign _002_ = in == 8'h9d;
  assign _003_ = in == 8'h9c;
  assign _004_ = in == 8'h9b;
  assign _005_ = in == 8'h9a;
  assign _006_ = in == 8'h99;
  assign _007_ = in == 8'h98;
  assign _008_ = in == 8'h97;
  assign _009_ = in == 8'h96;
  assign _010_ = in == 8'h95;
  assign _011_ = in == 8'hf8;
  assign _012_ = in == 8'h94;
  assign _013_ = in == 8'h93;
  assign _014_ = in == 8'h92;
  assign _015_ = in == 8'h91;
  assign _016_ = in == 8'h90;
  assign _017_ = in == 8'h8f;
  assign _018_ = in == 8'h8e;
  assign _019_ = in == 8'h8d;
  assign _020_ = in == 8'h8c;
  assign _021_ = in == 8'h8b;
  assign _022_ = in == 8'hf7;
  assign _023_ = in == 8'h8a;
  assign _024_ = in == 8'h89;
  assign _025_ = in == 8'h88;
  assign _026_ = in == 8'h87;
  assign _027_ = in == 8'h86;
  assign _028_ = in == 8'h85;
  assign _029_ = in == 8'h84;
  assign _030_ = in == 8'h83;
  assign _031_ = in == 8'h82;
  assign _032_ = in == 8'h81;
  assign _033_ = in == 8'hf6;
  assign _034_ = in == 8'h80;
  assign _035_ = in == 7'h7f;
  assign _036_ = in == 7'h7e;
  assign _037_ = in == 7'h7d;
  assign _038_ = in == 7'h7c;
  assign _039_ = in == 7'h7b;
  assign _040_ = in == 7'h7a;
  assign _041_ = in == 7'h79;
  assign _042_ = in == 7'h78;
  assign _043_ = in == 7'h77;
  assign _044_ = in == 8'hf5;
  assign _045_ = in == 7'h76;
  assign _046_ = in == 7'h75;
  assign _047_ = in == 7'h74;
  assign _048_ = in == 7'h73;
  assign _049_ = in == 7'h72;
  assign _050_ = in == 7'h71;
  assign _051_ = in == 7'h70;
  assign _052_ = in == 7'h6f;
  assign _053_ = in == 7'h6e;
  assign _054_ = in == 7'h6d;
  assign _055_ = in == 8'hf4;
  assign _056_ = in == 7'h6c;
  assign _057_ = in == 7'h6b;
  assign _058_ = in == 7'h6a;
  assign _059_ = in == 7'h69;
  assign _060_ = in == 7'h68;
  assign _061_ = in == 7'h67;
  assign _062_ = in == 7'h66;
  assign _063_ = in == 7'h65;
  assign _064_ = in == 7'h64;
  assign _065_ = in == 7'h63;
  assign _066_ = in == 8'hf3;
  assign _067_ = in == 7'h62;
  assign _068_ = in == 7'h61;
  assign _069_ = in == 7'h60;
  assign _070_ = in == 7'h5f;
  assign _071_ = in == 7'h5e;
  assign _072_ = in == 7'h5d;
  assign _073_ = in == 7'h5c;
  assign _074_ = in == 7'h5b;
  assign _075_ = in == 7'h5a;
  assign _076_ = in == 7'h59;
  assign _077_ = in == 8'hf2;
  assign _078_ = in == 7'h58;
  assign _079_ = in == 7'h57;
  assign _080_ = in == 7'h56;
  assign _081_ = in == 7'h55;
  assign _082_ = in == 7'h54;
  assign _083_ = in == 7'h53;
  assign _084_ = in == 7'h52;
  assign _085_ = in == 7'h51;
  assign _086_ = in == 7'h50;
  assign _087_ = in == 7'h4f;
  assign _088_ = in == 8'hf1;
  assign _089_ = in == 7'h4e;
  assign _090_ = in == 7'h4d;
  assign _091_ = in == 7'h4c;
  assign _092_ = in == 7'h4b;
  assign _093_ = in == 7'h4a;
  assign _094_ = in == 7'h49;
  assign _095_ = in == 7'h48;
  assign _096_ = in == 7'h47;
  assign _097_ = in == 7'h46;
  assign _098_ = in == 7'h45;
  assign _099_ = in == 8'hf0;
  assign _100_ = in == 7'h44;
  assign _101_ = in == 7'h43;
  assign _102_ = in == 7'h42;
  assign _103_ = in == 7'h41;
  assign _104_ = in == 7'h40;
  assign _105_ = in == 6'h3f;
  assign _106_ = in == 6'h3e;
  assign _107_ = in == 6'h3d;
  assign _108_ = in == 6'h3c;
  assign _109_ = in == 6'h3b;
  assign _110_ = in == 8'hef;
  logic [255:0] fangyuan0;
  assign fangyuan0 = { _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _131_, _130_, _129_, _128_, _127_, _126_, _125_, _124_, _123_, _122_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_, _098_, _097_, _096_, _095_, _094_, _093_, _092_, _091_, _090_, _089_, _087_, _086_, _085_, _084_, _083_, _082_, _081_, _080_, _079_, _078_, _076_, _075_, _074_, _073_, _072_, _071_, _070_, _069_, _068_, _067_, _065_, _064_, _063_, _062_, _061_, _060_, _059_, _058_, _057_, _056_, _054_, _053_, _052_, _051_, _050_, _049_, _048_, _047_, _046_, _045_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_, _035_, _034_, _032_, _031_, _030_, _029_, _028_, _027_, _026_, _025_, _024_, _023_, _021_, _020_, _019_, _018_, _017_, _016_, _015_, _014_, _013_, _012_, _010_, _009_, _008_, _007_, _006_, _005_, _004_, _003_, _002_, _001_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _165_, _154_, _143_, _132_, _121_, _110_, _099_, _088_, _077_, _066_, _055_, _044_, _033_, _022_, _011_, _256_, _245_, _234_, _223_, _212_, _201_, _190_ };

  always @(out or fangyuan0) begin
    casez (fangyuan0)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1 :
        _000_ = 8'b00010110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1? :
        _000_ = 8'b10111011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?? :
        _000_ = 8'b01010100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??? :
        _000_ = 8'b10110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???? :
        _000_ = 8'b00001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????? :
        _000_ = 8'b00101101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????? :
        _000_ = 8'b10011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????? :
        _000_ = 8'b01000001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????? :
        _000_ = 8'b01101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????? :
        _000_ = 8'b01000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????? :
        _000_ = 8'b11100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????? :
        _000_ = 8'b10111111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????? :
        _000_ = 8'b00001101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????? :
        _000_ = 8'b10001001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????? :
        _000_ = 8'b10100001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????? :
        _000_ = 8'b10001100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????? :
        _000_ = 8'b11011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????? :
        _000_ = 8'b00101000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????? :
        _000_ = 8'b01010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????? :
        _000_ = 8'b11001110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????? :
        _000_ = 8'b11101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????? :
        _000_ = 8'b10000111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????? :
        _000_ = 8'b00011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????? :
        _000_ = 8'b10011011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????? :
        _000_ = 8'b10010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????? :
        _000_ = 8'b10001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????? :
        _000_ = 8'b11011001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????? :
        _000_ = 8'b01101001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????? :
        _000_ = 8'b00010001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????? :
        _000_ = 8'b10011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????? :
        _000_ = 8'b11111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????? :
        _000_ = 8'b11100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????? :
        _000_ = 8'b10011110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????? :
        _000_ = 8'b00011101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????? :
        _000_ = 8'b11000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????? :
        _000_ = 8'b10000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????? :
        _000_ = 8'b10111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????? :
        _000_ = 8'b01010111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????? :
        _000_ = 8'b00110101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????? :
        _000_ = 8'b01100001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????? :
        _000_ = 8'b00001110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????? :
        _000_ = 8'b11110110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????? :
        _000_ = 8'b00000011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????? :
        _000_ = 8'b01001000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????? :
        _000_ = 8'b01100110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????? :
        _000_ = 8'b10110101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????? :
        _000_ = 8'b00111110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????? :
        _000_ = 8'b01110000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????? :
        _000_ = 8'b10001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????? :
        _000_ = 8'b10001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????? :
        _000_ = 8'b10111101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????? :
        _000_ = 8'b01001011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????? :
        _000_ = 8'b00011111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????? :
        _000_ = 8'b01110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????? :
        _000_ = 8'b11011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????? :
        _000_ = 8'b11101000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????? :
        _000_ = 8'b11000110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????? :
        _000_ = 8'b10110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????? :
        _000_ = 8'b10100110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????? :
        _000_ = 8'b00011100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????? :
        _000_ = 8'b00101110 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100101 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001000 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000110 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10001000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101010 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000100 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011111 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101100 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010010 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110110 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111100 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010001 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101000 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011111 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111001 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000101 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110011 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001101 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000011 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101010 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101111 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001111 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01001010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111001 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10111110 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001011 ;
      256'b????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101010 ;
      256'b???????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011011 ;
      256'b??????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110001 ;
      256'b?????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111100 ;
      256'b????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100000 ;
      256'b???????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101101 ;
      256'b??????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000000 ;
      256'b?????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010001 ;
      256'b????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010011 ;
      256'b???????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000100 ;
      256'b??????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101111 ;
      256'b?????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100011 ;
      256'b????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101001 ;
      256'b???????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110011 ;
      256'b??????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010110 ;
      256'b?????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111011 ;
      256'b????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01010010 ;
      256'b???????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100000 ;
      256'b??????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011010 ;
      256'b?????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101110 ;
      256'b????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011011 ;
      256'b???????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011010 ;
      256'b??????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101100 ;
      256'b?????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000011 ;
      256'b????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00001001 ;
      256'b???????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110101 ;
      256'b??????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110010 ;
      256'b?????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100111 ;
      256'b????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11101011 ;
      256'b???????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100010 ;
      256'b??????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000000 ;
      256'b?????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010010 ;
      256'b????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000111 ;
      256'b???????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011010 ;
      256'b??????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000101 ;
      256'b?????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010110 ;
      256'b????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00011000 ;
      256'b???????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000011 ;
      256'b??????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100011 ;
      256'b?????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000111 ;
      256'b????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000100 ;
      256'b???????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00010101 ;
      256'b??????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110001 ;
      256'b?????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11011000 ;
      256'b????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110001 ;
      256'b???????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110001 ;
      256'b??????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11100101 ;
      256'b?????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100101 ;
      256'b????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110100 ;
      256'b???????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001100 ;
      256'b??????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110111 ;
      256'b?????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00111111 ;
      256'b????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110110 ;
      256'b???????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00100110 ;
      256'b??????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10010011 ;
      256'b?????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111101 ;
      256'b????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10110111 ;
      256'b???????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000000 ;
      256'b??????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110010 ;
      256'b?????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100100 ;
      256'b????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10011100 ;
      256'b???????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101111 ;
      256'b??????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10100010 ;
      256'b?????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010100 ;
      256'b????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101101 ;
      256'b???????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110000 ;
      256'b??????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01000111 ;
      256'b?????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01011001 ;
      256'b????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111010 ;
      256'b???????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111101 ;
      256'b??????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001001 ;
      256'b?????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10000010 ;
      256'b????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11001010 ;
      256'b???????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110110 ;
      256'b??????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b10101011 ;
      256'b?????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11010111 ;
      256'b????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11111110 ;
      256'b???????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00101011 ;
      256'b??????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100111 ;
      256'b?????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00000001 ;
      256'b????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b00110000 ;
      256'b???????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11000101 ;
      256'b??????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101111 ;
      256'b?????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01101011 ;
      256'b????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b11110010 ;
      256'b???1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111011 ;
      256'b??1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01110111 ;
      256'b?1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01111100 ;
      256'b1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????? :
        _000_ = 8'b01100011 ;
      default:
        _000_ = out ;
    endcase
  end
  assign _111_ = in == 6'h3a;
  assign _112_ = in == 6'h39;
  assign _113_ = in == 6'h38;
  assign _114_ = in == 6'h37;
  assign _115_ = in == 6'h36;
  assign _116_ = in == 6'h35;
  assign _117_ = in == 6'h34;
  assign _118_ = in == 6'h33;
  assign _119_ = in == 6'h32;
  assign _120_ = in == 6'h31;
  assign _121_ = in == 8'hee;
  assign _122_ = in == 6'h30;
  assign _123_ = in == 6'h2f;
  assign _124_ = in == 6'h2e;
  assign _125_ = in == 6'h2d;
  assign _126_ = in == 6'h2c;
  assign _127_ = in == 6'h2b;
  assign _128_ = in == 6'h2a;
  assign _129_ = in == 6'h29;
  assign _130_ = in == 6'h28;
  assign _131_ = in == 6'h27;
  assign _132_ = in == 8'hed;
  assign _133_ = in == 6'h26;
  assign _134_ = in == 6'h25;
  assign _135_ = in == 6'h24;
  assign _136_ = in == 6'h23;
  assign _137_ = in == 6'h22;
  assign _138_ = in == 6'h21;
  assign _139_ = in == 6'h20;
  assign _140_ = in == 5'h1f;
  assign _141_ = in == 5'h1e;
  assign _142_ = in == 5'h1d;
  assign _143_ = in == 8'hec;
  assign _144_ = in == 5'h1c;
  assign _145_ = in == 5'h1b;
  assign _146_ = in == 5'h1a;
  assign _147_ = in == 5'h19;
  assign _148_ = in == 5'h18;
  assign _149_ = in == 5'h17;
  assign _150_ = in == 5'h16;
  assign _151_ = in == 5'h15;
  assign _152_ = in == 5'h14;
  assign _153_ = in == 5'h13;
  assign _154_ = in == 8'heb;
  assign _155_ = in == 5'h12;
  assign _156_ = in == 5'h11;
  assign _157_ = in == 5'h10;
  assign _158_ = in == 4'hf;
  assign _159_ = in == 4'he;
  assign _160_ = in == 4'hd;
  assign _161_ = in == 4'hc;
  assign _162_ = in == 4'hb;
  assign _163_ = in == 4'ha;
  assign _164_ = in == 4'h9;
  assign _165_ = in == 8'hea;
  assign _166_ = in == 4'h8;
  assign _167_ = in == 3'h7;
  assign _168_ = in == 3'h6;
  assign _169_ = in == 3'h5;
  assign _170_ = in == 3'h4;
  assign _171_ = in == 2'h3;
  assign _172_ = in == 2'h2;
  assign _173_ = in == 1'h1;
  assign _174_ = ! in;
  assign _175_ = in == 8'he9;
  assign _176_ = in == 8'he8;
  assign _177_ = in == 8'he7;
  assign _178_ = in == 8'he6;
  assign _179_ = in == 8'he5;
  assign _180_ = in == 8'he4;
  assign _181_ = in == 8'he3;
  assign _182_ = in == 8'he2;
  assign _183_ = in == 8'he1;
  assign _184_ = in == 8'he0;
  assign _185_ = in == 8'hdf;
  assign _186_ = in == 8'hde;
  assign _187_ = in == 8'hdd;
  assign _188_ = in == 8'hdc;
  assign _189_ = in == 8'hdb;
  assign _190_ = in == 8'hff;
  assign _191_ = in == 8'hda;
  assign _192_ = in == 8'hd9;
  assign _193_ = in == 8'hd8;
  assign _194_ = in == 8'hd7;
  assign _195_ = in == 8'hd6;
  assign _196_ = in == 8'hd5;
  assign _197_ = in == 8'hd4;
  assign _198_ = in == 8'hd3;
  assign _199_ = in == 8'hd2;
  assign _200_ = in == 8'hd1;
  assign _201_ = in == 8'hfe;
  assign _202_ = in == 8'hd0;
  assign _203_ = in == 8'hcf;
  assign _204_ = in == 8'hce;
  assign _205_ = in == 8'hcd;
  assign _206_ = in == 8'hcc;
  assign _207_ = in == 8'hcb;
  assign _208_ = in == 8'hca;
  assign _209_ = in == 8'hc9;
  assign _210_ = in == 8'hc8;
  assign _211_ = in == 8'hc7;
  assign _212_ = in == 8'hfd;
  assign _213_ = in == 8'hc6;
  assign _214_ = in == 8'hc5;
  assign _215_ = in == 8'hc4;
  assign _216_ = in == 8'hc3;
  assign _217_ = in == 8'hc2;
  assign _218_ = in == 8'hc1;
  assign _219_ = in == 8'hc0;
  assign _220_ = in == 8'hbf;
  assign _221_ = in == 8'hbe;
  assign _222_ = in == 8'hbd;
  assign _223_ = in == 8'hfc;
  assign _224_ = in == 8'hbc;
  assign _225_ = in == 8'hbb;
  assign _226_ = in == 8'hba;
  assign _227_ = in == 8'hb9;
  assign _228_ = in == 8'hb8;
  assign _229_ = in == 8'hb7;
  assign _230_ = in == 8'hb6;
  assign _231_ = in == 8'hb5;
  assign _232_ = in == 8'hb4;
  assign _233_ = in == 8'hb3;
  assign _234_ = in == 8'hfb;
  assign _235_ = in == 8'hb2;
  assign _236_ = in == 8'hb1;
  assign _237_ = in == 8'hb0;
  assign _238_ = in == 8'haf;
  assign _239_ = in == 8'hae;
  assign _240_ = in == 8'had;
  assign _241_ = in == 8'hac;
  assign _242_ = in == 8'hab;
  assign _243_ = in == 8'haa;
  assign _244_ = in == 8'ha9;
  assign _245_ = in == 8'hfa;
  assign _246_ = in == 8'ha8;
  assign _247_ = in == 8'ha7;
  assign _248_ = in == 8'ha6;
  assign _249_ = in == 8'ha5;
  assign _250_ = in == 8'ha4;
  assign _251_ = in == 8'ha3;
  assign _252_ = in == 8'ha2;
  assign _253_ = in == 8'ha1;
  assign _254_ = in == 8'ha0;
  assign _255_ = in == 8'h9f;
  assign _256_ = in == 8'hf9;
endmodule
