module AesCombined(clock, reset, io_encDataIn, io_encIvIn, io_encDataValid, io_decDataIn, io_decIvIn, io_decDataValid, io_aes256, io_keyIn, io_keyShift, io_keyValid, io_encReady, io_decReady, io_encDataOut, io_encIvOut, io_encOutputValid, io_decDataOut, io_decIvOut, io_decOutputValid);
  (* src = "crypto_accelerator.v:8041" *)
  wire [5:0] _000_;
  (* src = "crypto_accelerator.v:8041" *)
  wire _001_;
  (* src = "crypto_accelerator.v:7345" *)
  wire _002_;
  (* src = "crypto_accelerator.v:7346" *)
  wire _003_;
  (* src = "crypto_accelerator.v:7347" *)
  wire _004_;
  (* src = "crypto_accelerator.v:7348" *)
  wire _005_;
  (* src = "crypto_accelerator.v:7349" *)
  wire _006_;
  (* src = "crypto_accelerator.v:7350" *)
  wire _007_;
  (* src = "crypto_accelerator.v:7351" *)
  wire _008_;
  (* src = "crypto_accelerator.v:7352" *)
  wire _009_;
  (* src = "crypto_accelerator.v:7353" *)
  wire _010_;
  (* src = "crypto_accelerator.v:7354" *)
  wire _011_;
  (* src = "crypto_accelerator.v:7355" *)
  wire _012_;
  (* src = "crypto_accelerator.v:7356" *)
  wire _013_;
  (* src = "crypto_accelerator.v:7357" *)
  wire _014_;
  (* src = "crypto_accelerator.v:7358" *)
  wire _015_;
  (* src = "crypto_accelerator.v:7360" *)
  wire _016_;
  (* src = "crypto_accelerator.v:7361" *)
  wire _017_;
  (* src = "crypto_accelerator.v:7362" *)
  wire _018_;
  (* src = "crypto_accelerator.v:7363" *)
  wire _019_;
  (* src = "crypto_accelerator.v:7364" *)
  wire _020_;
  (* src = "crypto_accelerator.v:7365" *)
  wire _021_;
  (* src = "crypto_accelerator.v:7366" *)
  wire _022_;
  (* src = "crypto_accelerator.v:7367" *)
  wire _023_;
  (* src = "crypto_accelerator.v:7368" *)
  wire _024_;
  (* src = "crypto_accelerator.v:7369" *)
  wire _025_;
  (* src = "crypto_accelerator.v:7370" *)
  wire _026_;
  (* src = "crypto_accelerator.v:7371" *)
  wire _027_;
  (* src = "crypto_accelerator.v:7372" *)
  wire _028_;
  (* src = "crypto_accelerator.v:7373" *)
  wire _029_;
  wire [5:0] _030_;
  wire [5:0] _031_;
  wire _032_;
  wire _033_;
  (* src = "crypto_accelerator.v:6798" *)
  wire _GEN_0;
  wire [4:0] _GEN_10;
  wire [5:0] _GEN_11;
  wire [6:0] _GEN_12;
  (* src = "crypto_accelerator.v:7351" *)
  wire [7:0] _GEN_13;
  (* src = "crypto_accelerator.v:7352" *)
  wire [7:0] _GEN_14;
  (* src = "crypto_accelerator.v:7353" *)
  wire [7:0] _GEN_15;
  (* src = "crypto_accelerator.v:7354" *)
  wire [7:0] _GEN_16;
  (* src = "crypto_accelerator.v:7355" *)
  wire [7:0] _GEN_17;
  (* src = "crypto_accelerator.v:7356" *)
  wire [7:0] _GEN_18;
  (* src = "crypto_accelerator.v:7357" *)
  wire [7:0] _GEN_19;
  (* src = "crypto_accelerator.v:7358" *)
  wire [7:0] _GEN_20;
  wire _GEN_22;
  wire [1:0] _GEN_23;
  wire [2:0] _GEN_24;
  wire [3:0] _GEN_25;
  wire [4:0] _GEN_26;
  wire [5:0] _GEN_27;
  wire [6:0] _GEN_28;
  (* src = "crypto_accelerator.v:7366" *)
  wire [7:0] _GEN_29;
  (* src = "crypto_accelerator.v:6800" *)
  wire [127:0] _GEN_3;
  (* src = "crypto_accelerator.v:7367" *)
  wire [7:0] _GEN_30;
  (* src = "crypto_accelerator.v:7368" *)
  wire [7:0] _GEN_31;
  (* src = "crypto_accelerator.v:7369" *)
  wire [7:0] _GEN_32;
  (* src = "crypto_accelerator.v:7370" *)
  wire [7:0] _GEN_33;
  (* src = "crypto_accelerator.v:7371" *)
  wire [7:0] _GEN_34;
  (* src = "crypto_accelerator.v:7372" *)
  wire [7:0] _GEN_35;
  (* src = "crypto_accelerator.v:7373" *)
  wire [7:0] _GEN_36;
  (* src = "crypto_accelerator.v:7399" *)
  wire _GEN_39;
  wire _GEN_42;
  wire _GEN_6;
  wire [1:0] _GEN_7;
  wire [2:0] _GEN_8;
  wire [3:0] _GEN_9;
  (* src = "crypto_accelerator.v:6799" *)
  wire _T;
  (* src = "crypto_accelerator.v:6822" *)
  wire _T_100;
  (* src = "crypto_accelerator.v:7259" *)
  wire _T_1001;
  (* src = "crypto_accelerator.v:7260" *)
  wire _T_1003;
  (* src = "crypto_accelerator.v:7261" *)
  wire _T_1005;
  (* src = "crypto_accelerator.v:7262" *)
  wire _T_1007;
  (* src = "crypto_accelerator.v:7263" *)
  wire _T_1009;
  (* src = "crypto_accelerator.v:7264" *)
  wire _T_1011;
  (* src = "crypto_accelerator.v:7265" *)
  wire _T_1013;
  (* src = "crypto_accelerator.v:7266" *)
  wire _T_1015;
  (* src = "crypto_accelerator.v:7267" *)
  wire _T_1017;
  (* src = "crypto_accelerator.v:7268" *)
  wire _T_1019;
  (* src = "crypto_accelerator.v:6823" *)
  wire _T_102;
  (* src = "crypto_accelerator.v:7269" *)
  wire _T_1021;
  (* src = "crypto_accelerator.v:7270" *)
  wire _T_1023;
  (* src = "crypto_accelerator.v:7271" *)
  wire _T_1025;
  (* src = "crypto_accelerator.v:7272" *)
  wire _T_1027;
  (* src = "crypto_accelerator.v:7273" *)
  wire _T_1029;
  (* src = "crypto_accelerator.v:7274" *)
  wire _T_1031;
  (* src = "crypto_accelerator.v:7275" *)
  wire _T_1033;
  (* src = "crypto_accelerator.v:7276" *)
  wire _T_1035;
  (* src = "crypto_accelerator.v:7277" *)
  wire _T_1037;
  (* src = "crypto_accelerator.v:7278" *)
  wire _T_1039;
  (* src = "crypto_accelerator.v:6824" *)
  wire _T_104;
  (* src = "crypto_accelerator.v:7279" *)
  wire _T_1041;
  (* src = "crypto_accelerator.v:7280" *)
  wire _T_1043;
  (* src = "crypto_accelerator.v:7281" *)
  wire _T_1045;
  (* src = "crypto_accelerator.v:7282" *)
  wire _T_1047;
  (* src = "crypto_accelerator.v:7283" *)
  wire _T_1049;
  (* src = "crypto_accelerator.v:7284" *)
  wire _T_1051;
  (* src = "crypto_accelerator.v:7285" *)
  wire _T_1053;
  (* src = "crypto_accelerator.v:7286" *)
  wire _T_1055;
  (* src = "crypto_accelerator.v:7287" *)
  wire _T_1057;
  (* src = "crypto_accelerator.v:7288" *)
  wire _T_1059;
  (* src = "crypto_accelerator.v:6825" *)
  wire _T_106;
  (* src = "crypto_accelerator.v:7289" *)
  wire _T_1061;
  (* src = "crypto_accelerator.v:7290" *)
  wire _T_1063;
  (* src = "crypto_accelerator.v:7291" *)
  wire _T_1065;
  (* src = "crypto_accelerator.v:7292" *)
  wire _T_1067;
  (* src = "crypto_accelerator.v:7293" *)
  wire _T_1069;
  (* src = "crypto_accelerator.v:7294" *)
  wire _T_1071;
  (* src = "crypto_accelerator.v:7295" *)
  wire _T_1073;
  (* src = "crypto_accelerator.v:7296" *)
  wire _T_1075;
  (* src = "crypto_accelerator.v:7297" *)
  wire _T_1077;
  (* src = "crypto_accelerator.v:7298" *)
  wire _T_1079;
  (* src = "crypto_accelerator.v:6826" *)
  wire _T_108;
  (* src = "crypto_accelerator.v:7299" *)
  wire _T_1081;
  (* src = "crypto_accelerator.v:7300" *)
  wire _T_1083;
  (* src = "crypto_accelerator.v:7301" *)
  wire _T_1085;
  (* src = "crypto_accelerator.v:7302" *)
  wire _T_1087;
  (* src = "crypto_accelerator.v:7303" *)
  wire _T_1089;
  (* src = "crypto_accelerator.v:7304" *)
  wire _T_1091;
  (* src = "crypto_accelerator.v:7305" *)
  wire _T_1093;
  (* src = "crypto_accelerator.v:7306" *)
  wire _T_1094;
  (* src = "crypto_accelerator.v:7307" *)
  wire _T_1095;
  (* src = "crypto_accelerator.v:7308" *)
  wire _T_1096;
  (* src = "crypto_accelerator.v:7309" *)
  wire _T_1098;
  (* src = "crypto_accelerator.v:7310" *)
  wire _T_1099;
  (* src = "crypto_accelerator.v:6827" *)
  wire _T_110;
  (* src = "crypto_accelerator.v:7311" *)
  wire _T_1100;
  (* src = "crypto_accelerator.v:7312" *)
  wire _T_1102;
  (* src = "crypto_accelerator.v:7313" *)
  wire _T_1104;
  (* src = "crypto_accelerator.v:7314" *)
  wire _T_1105;
  (* src = "crypto_accelerator.v:7315" *)
  wire _T_1106;
  (* src = "crypto_accelerator.v:7316" *)
  wire _T_1108;
  (* src = "crypto_accelerator.v:7317" *)
  wire _T_1110;
  (* src = "crypto_accelerator.v:7318" *)
  wire _T_1112;
  (* src = "crypto_accelerator.v:7319" *)
  wire _T_1113;
  (* src = "crypto_accelerator.v:7320" *)
  wire _T_1114;
  (* src = "crypto_accelerator.v:7321" *)
  wire _T_1116;
  (* src = "crypto_accelerator.v:7322" *)
  wire _T_1117;
  (* src = "crypto_accelerator.v:7323" *)
  wire _T_1119;
  (* src = "crypto_accelerator.v:6828" *)
  wire _T_112;
  (* src = "crypto_accelerator.v:7324" *)
  wire _T_1120;
  (* src = "crypto_accelerator.v:7325" *)
  wire _T_1121;
  (* src = "crypto_accelerator.v:7326" *)
  wire [7:0] _T_1128;
  (* src = "crypto_accelerator.v:7327" *)
  wire [7:0] _T_1129_0_0;
  (* src = "crypto_accelerator.v:7328" *)
  wire [7:0] _T_1129_0_1;
  (* src = "crypto_accelerator.v:7329" *)
  wire [7:0] _T_1129_0_2;
  (* src = "crypto_accelerator.v:7330" *)
  wire [7:0] _T_1129_0_3;
  (* src = "crypto_accelerator.v:7331" *)
  wire [7:0] _T_1129_1_0;
  (* src = "crypto_accelerator.v:7332" *)
  wire [7:0] _T_1129_1_1;
  (* src = "crypto_accelerator.v:7333" *)
  wire [7:0] _T_1129_1_2;
  (* src = "crypto_accelerator.v:7334" *)
  wire [7:0] _T_1129_1_3;
  (* src = "crypto_accelerator.v:7335" *)
  wire [7:0] _T_1129_2_0;
  (* src = "crypto_accelerator.v:7336" *)
  wire [7:0] _T_1129_2_1;
  (* src = "crypto_accelerator.v:7337" *)
  wire [7:0] _T_1129_2_2;
  (* src = "crypto_accelerator.v:7338" *)
  wire [7:0] _T_1129_2_3;
  (* src = "crypto_accelerator.v:7339" *)
  wire [7:0] _T_1129_3_0;
  (* src = "crypto_accelerator.v:7340" *)
  wire [7:0] _T_1129_3_1;
  (* src = "crypto_accelerator.v:7341" *)
  wire [7:0] _T_1129_3_2;
  (* src = "crypto_accelerator.v:7342" *)
  wire [7:0] _T_1129_3_3;
  wire [3:0] _T_1133;
  (* src = "crypto_accelerator.v:7374" *)
  wire [7:0] _T_1137;
  (* src = "crypto_accelerator.v:7375" *)
  wire [7:0] _T_1138;
  (* src = "crypto_accelerator.v:7376" *)
  wire [7:0] _T_1139;
  (* src = "crypto_accelerator.v:6829" *)
  wire _T_114;
  (* src = "crypto_accelerator.v:7377" *)
  wire [7:0] _T_1140;
  (* src = "crypto_accelerator.v:7378" *)
  wire [7:0] _T_1141;
  (* src = "crypto_accelerator.v:7379" *)
  wire [7:0] _T_1142;
  (* src = "crypto_accelerator.v:7380" *)
  wire [7:0] _T_1143;
  (* src = "crypto_accelerator.v:7381" *)
  wire [7:0] _T_1144;
  (* src = "crypto_accelerator.v:7382" *)
  wire [7:0] _T_1145;
  (* src = "crypto_accelerator.v:7383" *)
  wire [7:0] _T_1146;
  (* src = "crypto_accelerator.v:7384" *)
  wire [7:0] _T_1147;
  (* src = "crypto_accelerator.v:7385" *)
  wire [7:0] _T_1149;
  (* src = "crypto_accelerator.v:7386" *)
  wire [7:0] _T_1150;
  (* src = "crypto_accelerator.v:7387" *)
  wire [7:0] _T_1151;
  (* src = "crypto_accelerator.v:7388" *)
  wire [7:0] _T_1152;
  (* src = "crypto_accelerator.v:7389" *)
  wire [7:0] _T_1154;
  (* src = "crypto_accelerator.v:7390" *)
  wire [7:0] _T_1155;
  (* src = "crypto_accelerator.v:7391" *)
  wire [7:0] _T_1156;
  (* src = "crypto_accelerator.v:7392" *)
  wire [7:0] _T_1157;
  (* src = "crypto_accelerator.v:7393" *)
  wire [7:0] _T_1159;
  (* src = "crypto_accelerator.v:6830" *)
  wire _T_116;
  (* src = "crypto_accelerator.v:7394" *)
  wire [7:0] _T_1160;
  (* src = "crypto_accelerator.v:7395" *)
  wire [7:0] _T_1161;
  (* src = "crypto_accelerator.v:7396" *)
  wire [7:0] _T_1162;
  (* src = "crypto_accelerator.v:7397" *)
  wire [63:0] _T_1170;
  (* src = "crypto_accelerator.v:7398" *)
  wire [127:0] _T_1178;
  (* src = "crypto_accelerator.v:6831" *)
  wire _T_118;
  (* src = "crypto_accelerator.v:6832" *)
  wire _T_120;
  (* src = "crypto_accelerator.v:6833" *)
  wire _T_122;
  (* src = "crypto_accelerator.v:6834" *)
  wire _T_124;
  (* src = "crypto_accelerator.v:6835" *)
  wire _T_126;
  (* src = "crypto_accelerator.v:6836" *)
  wire _T_128;
  (* src = "crypto_accelerator.v:6837" *)
  wire _T_130;
  (* src = "crypto_accelerator.v:6838" *)
  wire _T_132;
  (* src = "crypto_accelerator.v:6839" *)
  wire _T_134;
  (* src = "crypto_accelerator.v:6840" *)
  wire _T_136;
  (* src = "crypto_accelerator.v:6841" *)
  wire _T_138;
  (* src = "crypto_accelerator.v:6842" *)
  wire _T_140;
  (* src = "crypto_accelerator.v:6843" *)
  wire _T_142;
  (* src = "crypto_accelerator.v:6844" *)
  wire _T_144;
  (* src = "crypto_accelerator.v:6845" *)
  wire _T_146;
  (* src = "crypto_accelerator.v:6846" *)
  wire _T_148;
  (* src = "crypto_accelerator.v:7400" *)
  wire _T_1494;
  (* src = "crypto_accelerator.v:7401" *)
  wire _T_1495;
  (* src = "crypto_accelerator.v:7402" *)
  wire _T_1496;
  (* src = "crypto_accelerator.v:7403" *)
  wire _T_1499;
  (* src = "crypto_accelerator.v:6847" *)
  wire _T_150;
  (* src = "crypto_accelerator.v:7404" *)
  wire _T_1504;
  (* src = "crypto_accelerator.v:6848" *)
  wire _T_152;
  (* src = "crypto_accelerator.v:6849" *)
  wire _T_154;
  (* src = "crypto_accelerator.v:6850" *)
  wire _T_156;
  (* src = "crypto_accelerator.v:6851" *)
  wire _T_158;
  (* src = "crypto_accelerator.v:6852" *)
  wire _T_160;
  (* src = "crypto_accelerator.v:6853" *)
  wire _T_162;
  (* src = "crypto_accelerator.v:6854" *)
  wire _T_164;
  (* src = "crypto_accelerator.v:6855" *)
  wire _T_166;
  (* src = "crypto_accelerator.v:6856" *)
  wire _T_168;
  (* src = "crypto_accelerator.v:6857" *)
  wire _T_170;
  (* src = "crypto_accelerator.v:6858" *)
  wire _T_172;
  (* src = "crypto_accelerator.v:6859" *)
  wire _T_174;
  (* src = "crypto_accelerator.v:6860" *)
  wire _T_176;
  (* src = "crypto_accelerator.v:6861" *)
  wire _T_178;
  (* src = "crypto_accelerator.v:6862" *)
  wire _T_180;
  (* src = "crypto_accelerator.v:6863" *)
  wire _T_182;
  (* src = "crypto_accelerator.v:6864" *)
  wire _T_184;
  (* src = "crypto_accelerator.v:6865" *)
  wire _T_186;
  (* src = "crypto_accelerator.v:6866" *)
  wire _T_188;
  (* src = "crypto_accelerator.v:6867" *)
  wire _T_190;
  (* src = "crypto_accelerator.v:6868" *)
  wire _T_192;
  (* src = "crypto_accelerator.v:6869" *)
  wire _T_194;
  (* src = "crypto_accelerator.v:6870" *)
  wire _T_196;
  (* src = "crypto_accelerator.v:6871" *)
  wire _T_198;
  (* src = "crypto_accelerator.v:6801" *)
  wire [5:0] _T_2;
  (* src = "crypto_accelerator.v:6872" *)
  wire _T_200;
  (* src = "crypto_accelerator.v:6873" *)
  wire _T_202;
  (* src = "crypto_accelerator.v:6874" *)
  wire _T_204;
  (* src = "crypto_accelerator.v:6875" *)
  wire _T_206;
  (* src = "crypto_accelerator.v:6876" *)
  wire _T_208;
  (* src = "crypto_accelerator.v:6877" *)
  wire _T_210;
  (* src = "crypto_accelerator.v:6878" *)
  wire _T_212;
  (* src = "crypto_accelerator.v:6879" *)
  wire _T_214;
  (* src = "crypto_accelerator.v:6880" *)
  wire _T_216;
  (* src = "crypto_accelerator.v:6881" *)
  wire _T_218;
  (* src = "crypto_accelerator.v:6882" *)
  wire _T_220;
  (* src = "crypto_accelerator.v:6883" *)
  wire _T_222;
  (* src = "crypto_accelerator.v:6884" *)
  wire _T_224;
  (* src = "crypto_accelerator.v:6885" *)
  wire _T_226;
  (* src = "crypto_accelerator.v:6886" *)
  wire _T_228;
  (* src = "crypto_accelerator.v:6887" *)
  wire _T_230;
  (* src = "crypto_accelerator.v:6888" *)
  wire _T_232;
  (* src = "crypto_accelerator.v:6889" *)
  wire _T_234;
  (* src = "crypto_accelerator.v:6890" *)
  wire _T_236;
  (* src = "crypto_accelerator.v:6891" *)
  wire _T_238;
  (* src = "crypto_accelerator.v:6892" *)
  wire _T_240;
  (* src = "crypto_accelerator.v:6893" *)
  wire _T_242;
  (* src = "crypto_accelerator.v:6894" *)
  wire _T_244;
  (* src = "crypto_accelerator.v:6895" *)
  wire _T_246;
  (* src = "crypto_accelerator.v:6896" *)
  wire _T_248;
  (* src = "crypto_accelerator.v:6897" *)
  wire _T_250;
  (* src = "crypto_accelerator.v:6898" *)
  wire _T_252;
  (* src = "crypto_accelerator.v:6899" *)
  wire _T_254;
  (* src = "crypto_accelerator.v:6900" *)
  wire _T_256;
  (* src = "crypto_accelerator.v:6901" *)
  wire _T_258;
  (* src = "crypto_accelerator.v:6902" *)
  wire _T_260;
  (* src = "crypto_accelerator.v:6903" *)
  wire _T_262;
  (* src = "crypto_accelerator.v:6904" *)
  wire _T_264;
  (* src = "crypto_accelerator.v:6905" *)
  wire _T_266;
  (* src = "crypto_accelerator.v:6906" *)
  wire _T_268;
  (* src = "crypto_accelerator.v:6907" *)
  wire _T_270;
  (* src = "crypto_accelerator.v:6908" *)
  wire _T_272;
  (* src = "crypto_accelerator.v:6909" *)
  wire _T_274;
  (* src = "crypto_accelerator.v:6910" *)
  wire _T_276;
  (* src = "crypto_accelerator.v:6911" *)
  wire _T_278;
  (* src = "crypto_accelerator.v:6912" *)
  wire _T_280;
  (* src = "crypto_accelerator.v:6913" *)
  wire _T_282;
  (* src = "crypto_accelerator.v:6914" *)
  wire _T_284;
  (* src = "crypto_accelerator.v:6915" *)
  wire _T_286;
  (* src = "crypto_accelerator.v:6916" *)
  wire _T_287;
  (* src = "crypto_accelerator.v:6917" *)
  wire _T_288;
  (* src = "crypto_accelerator.v:6918" *)
  wire _T_289;
  (* src = "crypto_accelerator.v:6919" *)
  wire _T_291;
  (* src = "crypto_accelerator.v:6920" *)
  wire _T_292;
  (* src = "crypto_accelerator.v:6921" *)
  wire _T_293;
  (* src = "crypto_accelerator.v:6922" *)
  wire _T_295;
  (* src = "crypto_accelerator.v:6923" *)
  wire _T_297;
  (* src = "crypto_accelerator.v:6924" *)
  wire _T_298;
  (* src = "crypto_accelerator.v:6925" *)
  wire _T_299;
  (* src = "crypto_accelerator.v:6926" *)
  wire _T_301;
  (* src = "crypto_accelerator.v:6927" *)
  wire _T_303;
  (* src = "crypto_accelerator.v:6928" *)
  wire _T_305;
  (* src = "crypto_accelerator.v:6929" *)
  wire _T_306;
  (* src = "crypto_accelerator.v:6930" *)
  wire _T_307;
  (* src = "crypto_accelerator.v:6931" *)
  wire _T_309;
  (* src = "crypto_accelerator.v:6932" *)
  wire _T_310;
  (* src = "crypto_accelerator.v:6933" *)
  wire _T_312;
  (* src = "crypto_accelerator.v:6934" *)
  wire _T_313;
  (* src = "crypto_accelerator.v:6935" *)
  wire _T_314;
  (* src = "crypto_accelerator.v:6936" *)
  wire [7:0] _T_321;
  (* src = "crypto_accelerator.v:6937" *)
  wire _T_339;
  (* src = "crypto_accelerator.v:6938" *)
  wire _T_341;
  (* src = "crypto_accelerator.v:6939" *)
  wire _T_343;
  (* src = "crypto_accelerator.v:6940" *)
  wire _T_345;
  (* src = "crypto_accelerator.v:6941" *)
  wire _T_347;
  (* src = "crypto_accelerator.v:6942" *)
  wire _T_349;
  (* src = "crypto_accelerator.v:6943" *)
  wire _T_351;
  (* src = "crypto_accelerator.v:6944" *)
  wire _T_353;
  (* src = "crypto_accelerator.v:6945" *)
  wire _T_355;
  (* src = "crypto_accelerator.v:6946" *)
  wire _T_357;
  (* src = "crypto_accelerator.v:6947" *)
  wire _T_359;
  (* src = "crypto_accelerator.v:6948" *)
  wire _T_361;
  (* src = "crypto_accelerator.v:6949" *)
  wire _T_363;
  (* src = "crypto_accelerator.v:6950" *)
  wire _T_365;
  (* src = "crypto_accelerator.v:6951" *)
  wire _T_367;
  (* src = "crypto_accelerator.v:6952" *)
  wire _T_369;
  (* src = "crypto_accelerator.v:6953" *)
  wire _T_371;
  (* src = "crypto_accelerator.v:6954" *)
  wire _T_373;
  (* src = "crypto_accelerator.v:6955" *)
  wire _T_375;
  (* src = "crypto_accelerator.v:6956" *)
  wire _T_377;
  (* src = "crypto_accelerator.v:6957" *)
  wire _T_379;
  (* src = "crypto_accelerator.v:6958" *)
  wire _T_381;
  (* src = "crypto_accelerator.v:6959" *)
  wire _T_383;
  (* src = "crypto_accelerator.v:6960" *)
  wire _T_385;
  (* src = "crypto_accelerator.v:6961" *)
  wire _T_387;
  (* src = "crypto_accelerator.v:6962" *)
  wire _T_389;
  (* src = "crypto_accelerator.v:6963" *)
  wire _T_391;
  (* src = "crypto_accelerator.v:6964" *)
  wire _T_393;
  (* src = "crypto_accelerator.v:6965" *)
  wire _T_395;
  (* src = "crypto_accelerator.v:6966" *)
  wire _T_397;
  (* src = "crypto_accelerator.v:6967" *)
  wire _T_399;
  (* src = "crypto_accelerator.v:6968" *)
  wire _T_401;
  (* src = "crypto_accelerator.v:6969" *)
  wire _T_403;
  (* src = "crypto_accelerator.v:6970" *)
  wire _T_405;
  (* src = "crypto_accelerator.v:6971" *)
  wire _T_407;
  (* src = "crypto_accelerator.v:6972" *)
  wire _T_409;
  (* src = "crypto_accelerator.v:6973" *)
  wire _T_411;
  (* src = "crypto_accelerator.v:6974" *)
  wire _T_413;
  (* src = "crypto_accelerator.v:6975" *)
  wire _T_415;
  (* src = "crypto_accelerator.v:6976" *)
  wire _T_417;
  (* src = "crypto_accelerator.v:6977" *)
  wire _T_419;
  (* src = "crypto_accelerator.v:6978" *)
  wire _T_421;
  (* src = "crypto_accelerator.v:6979" *)
  wire _T_423;
  (* src = "crypto_accelerator.v:6980" *)
  wire _T_425;
  (* src = "crypto_accelerator.v:6981" *)
  wire _T_427;
  (* src = "crypto_accelerator.v:6982" *)
  wire _T_429;
  (* src = "crypto_accelerator.v:6983" *)
  wire _T_431;
  (* src = "crypto_accelerator.v:6984" *)
  wire _T_433;
  (* src = "crypto_accelerator.v:6985" *)
  wire _T_435;
  (* src = "crypto_accelerator.v:6986" *)
  wire _T_437;
  (* src = "crypto_accelerator.v:6987" *)
  wire _T_439;
  (* src = "crypto_accelerator.v:6988" *)
  wire _T_441;
  (* src = "crypto_accelerator.v:6989" *)
  wire _T_443;
  (* src = "crypto_accelerator.v:6990" *)
  wire _T_445;
  (* src = "crypto_accelerator.v:6991" *)
  wire _T_447;
  (* src = "crypto_accelerator.v:6992" *)
  wire _T_449;
  (* src = "crypto_accelerator.v:6993" *)
  wire _T_451;
  (* src = "crypto_accelerator.v:6994" *)
  wire _T_453;
  (* src = "crypto_accelerator.v:6995" *)
  wire _T_455;
  (* src = "crypto_accelerator.v:6996" *)
  wire _T_457;
  (* src = "crypto_accelerator.v:6997" *)
  wire _T_459;
  (* src = "crypto_accelerator.v:6998" *)
  wire _T_461;
  (* src = "crypto_accelerator.v:6999" *)
  wire _T_463;
  (* src = "crypto_accelerator.v:7000" *)
  wire _T_465;
  (* src = "crypto_accelerator.v:7001" *)
  wire _T_467;
  (* src = "crypto_accelerator.v:7002" *)
  wire _T_469;
  (* src = "crypto_accelerator.v:7003" *)
  wire _T_471;
  (* src = "crypto_accelerator.v:7004" *)
  wire _T_473;
  (* src = "crypto_accelerator.v:7005" *)
  wire _T_475;
  (* src = "crypto_accelerator.v:7006" *)
  wire _T_477;
  (* src = "crypto_accelerator.v:7007" *)
  wire _T_479;
  (* src = "crypto_accelerator.v:7008" *)
  wire _T_481;
  (* src = "crypto_accelerator.v:7009" *)
  wire _T_483;
  (* src = "crypto_accelerator.v:7010" *)
  wire _T_485;
  (* src = "crypto_accelerator.v:7011" *)
  wire _T_487;
  (* src = "crypto_accelerator.v:7012" *)
  wire _T_489;
  (* src = "crypto_accelerator.v:7013" *)
  wire _T_491;
  (* src = "crypto_accelerator.v:7014" *)
  wire _T_493;
  (* src = "crypto_accelerator.v:7015" *)
  wire _T_495;
  (* src = "crypto_accelerator.v:7016" *)
  wire _T_497;
  (* src = "crypto_accelerator.v:7017" *)
  wire _T_499;
  wire _T_5;
  (* src = "crypto_accelerator.v:7018" *)
  wire _T_501;
  (* src = "crypto_accelerator.v:7019" *)
  wire _T_503;
  (* src = "crypto_accelerator.v:7020" *)
  wire _T_505;
  (* src = "crypto_accelerator.v:7021" *)
  wire _T_507;
  (* src = "crypto_accelerator.v:7022" *)
  wire _T_509;
  (* src = "crypto_accelerator.v:6805" *)
  wire _T_51;
  (* src = "crypto_accelerator.v:7023" *)
  wire _T_511;
  (* src = "crypto_accelerator.v:7024" *)
  wire _T_513;
  (* src = "crypto_accelerator.v:7025" *)
  wire _T_515;
  (* src = "crypto_accelerator.v:7026" *)
  wire _T_517;
  (* src = "crypto_accelerator.v:7027" *)
  wire _T_519;
  (* src = "crypto_accelerator.v:6806" *)
  wire _T_52;
  (* src = "crypto_accelerator.v:7028" *)
  wire _T_521;
  (* src = "crypto_accelerator.v:7029" *)
  wire _T_523;
  (* src = "crypto_accelerator.v:7030" *)
  wire _T_525;
  (* src = "crypto_accelerator.v:7031" *)
  wire _T_527;
  (* src = "crypto_accelerator.v:7032" *)
  wire _T_529;
  (* src = "crypto_accelerator.v:7033" *)
  wire _T_531;
  (* src = "crypto_accelerator.v:7034" *)
  wire _T_533;
  (* src = "crypto_accelerator.v:7035" *)
  wire _T_535;
  (* src = "crypto_accelerator.v:7036" *)
  wire _T_537;
  (* src = "crypto_accelerator.v:7037" *)
  wire _T_539;
  (* src = "crypto_accelerator.v:7038" *)
  wire _T_541;
  (* src = "crypto_accelerator.v:7039" *)
  wire _T_543;
  (* src = "crypto_accelerator.v:7040" *)
  wire _T_545;
  (* src = "crypto_accelerator.v:7041" *)
  wire _T_547;
  (* src = "crypto_accelerator.v:7042" *)
  wire _T_549;
  (* src = "crypto_accelerator.v:7043" *)
  wire _T_551;
  (* src = "crypto_accelerator.v:7044" *)
  wire _T_553;
  (* src = "crypto_accelerator.v:7045" *)
  wire _T_555;
  (* src = "crypto_accelerator.v:7046" *)
  wire _T_556;
  (* src = "crypto_accelerator.v:7047" *)
  wire _T_557;
  (* src = "crypto_accelerator.v:7048" *)
  wire _T_558;
  (* src = "crypto_accelerator.v:7049" *)
  wire _T_560;
  (* src = "crypto_accelerator.v:7050" *)
  wire _T_561;
  (* src = "crypto_accelerator.v:7051" *)
  wire _T_562;
  (* src = "crypto_accelerator.v:7052" *)
  wire _T_564;
  (* src = "crypto_accelerator.v:7053" *)
  wire _T_566;
  (* src = "crypto_accelerator.v:7054" *)
  wire _T_567;
  (* src = "crypto_accelerator.v:7055" *)
  wire _T_568;
  (* src = "crypto_accelerator.v:7056" *)
  wire _T_570;
  (* src = "crypto_accelerator.v:7057" *)
  wire _T_572;
  (* src = "crypto_accelerator.v:7058" *)
  wire _T_574;
  (* src = "crypto_accelerator.v:7059" *)
  wire _T_575;
  (* src = "crypto_accelerator.v:7060" *)
  wire _T_576;
  (* src = "crypto_accelerator.v:7061" *)
  wire _T_578;
  (* src = "crypto_accelerator.v:7062" *)
  wire _T_579;
  (* src = "crypto_accelerator.v:7063" *)
  wire _T_581;
  (* src = "crypto_accelerator.v:7064" *)
  wire _T_582;
  (* src = "crypto_accelerator.v:7065" *)
  wire _T_583;
  (* src = "crypto_accelerator.v:7066" *)
  wire [7:0] _T_590;
  (* src = "crypto_accelerator.v:6804" *)
  wire _T_6;
  (* src = "crypto_accelerator.v:7067" *)
  wire _T_608;
  (* src = "crypto_accelerator.v:7068" *)
  wire _T_610;
  (* src = "crypto_accelerator.v:7069" *)
  wire _T_612;
  (* src = "crypto_accelerator.v:7070" *)
  wire _T_614;
  (* src = "crypto_accelerator.v:7071" *)
  wire _T_616;
  (* src = "crypto_accelerator.v:7072" *)
  wire _T_618;
  (* src = "crypto_accelerator.v:7073" *)
  wire _T_620;
  (* src = "crypto_accelerator.v:7074" *)
  wire _T_622;
  (* src = "crypto_accelerator.v:7075" *)
  wire _T_624;
  (* src = "crypto_accelerator.v:7076" *)
  wire _T_626;
  (* src = "crypto_accelerator.v:7077" *)
  wire _T_628;
  (* src = "crypto_accelerator.v:7078" *)
  wire _T_630;
  (* src = "crypto_accelerator.v:7079" *)
  wire _T_632;
  (* src = "crypto_accelerator.v:7080" *)
  wire _T_634;
  (* src = "crypto_accelerator.v:7081" *)
  wire _T_636;
  (* src = "crypto_accelerator.v:7082" *)
  wire _T_638;
  (* src = "crypto_accelerator.v:7083" *)
  wire _T_640;
  (* src = "crypto_accelerator.v:7084" *)
  wire _T_642;
  (* src = "crypto_accelerator.v:7085" *)
  wire _T_644;
  (* src = "crypto_accelerator.v:7086" *)
  wire _T_646;
  (* src = "crypto_accelerator.v:7087" *)
  wire _T_648;
  (* src = "crypto_accelerator.v:7088" *)
  wire _T_650;
  (* src = "crypto_accelerator.v:7089" *)
  wire _T_652;
  (* src = "crypto_accelerator.v:7090" *)
  wire _T_654;
  (* src = "crypto_accelerator.v:7091" *)
  wire _T_656;
  (* src = "crypto_accelerator.v:7092" *)
  wire _T_658;
  (* src = "crypto_accelerator.v:7093" *)
  wire _T_660;
  (* src = "crypto_accelerator.v:7094" *)
  wire _T_662;
  (* src = "crypto_accelerator.v:7095" *)
  wire _T_664;
  (* src = "crypto_accelerator.v:7096" *)
  wire _T_666;
  (* src = "crypto_accelerator.v:7097" *)
  wire _T_668;
  (* src = "crypto_accelerator.v:7098" *)
  wire _T_670;
  (* src = "crypto_accelerator.v:7099" *)
  wire _T_672;
  (* src = "crypto_accelerator.v:7100" *)
  wire _T_674;
  (* src = "crypto_accelerator.v:7101" *)
  wire _T_676;
  (* src = "crypto_accelerator.v:7102" *)
  wire _T_678;
  (* src = "crypto_accelerator.v:7103" *)
  wire _T_680;
  (* src = "crypto_accelerator.v:7104" *)
  wire _T_682;
  (* src = "crypto_accelerator.v:7105" *)
  wire _T_684;
  (* src = "crypto_accelerator.v:7106" *)
  wire _T_686;
  (* src = "crypto_accelerator.v:7107" *)
  wire _T_688;
  (* src = "crypto_accelerator.v:7108" *)
  wire _T_690;
  (* src = "crypto_accelerator.v:7109" *)
  wire _T_692;
  (* src = "crypto_accelerator.v:7110" *)
  wire _T_694;
  (* src = "crypto_accelerator.v:7111" *)
  wire _T_696;
  (* src = "crypto_accelerator.v:7112" *)
  wire _T_698;
  (* src = "crypto_accelerator.v:6807" *)
  wire _T_70;
  (* src = "crypto_accelerator.v:7113" *)
  wire _T_700;
  (* src = "crypto_accelerator.v:7114" *)
  wire _T_702;
  (* src = "crypto_accelerator.v:7115" *)
  wire _T_704;
  (* src = "crypto_accelerator.v:7116" *)
  wire _T_706;
  (* src = "crypto_accelerator.v:7117" *)
  wire _T_708;
  (* src = "crypto_accelerator.v:7118" *)
  wire _T_710;
  (* src = "crypto_accelerator.v:7119" *)
  wire _T_712;
  (* src = "crypto_accelerator.v:7120" *)
  wire _T_714;
  (* src = "crypto_accelerator.v:7121" *)
  wire _T_716;
  (* src = "crypto_accelerator.v:7122" *)
  wire _T_718;
  (* src = "crypto_accelerator.v:6808" *)
  wire _T_72;
  (* src = "crypto_accelerator.v:7123" *)
  wire _T_720;
  (* src = "crypto_accelerator.v:7124" *)
  wire _T_722;
  (* src = "crypto_accelerator.v:7125" *)
  wire _T_724;
  (* src = "crypto_accelerator.v:7126" *)
  wire _T_726;
  (* src = "crypto_accelerator.v:7127" *)
  wire _T_728;
  (* src = "crypto_accelerator.v:7128" *)
  wire _T_730;
  (* src = "crypto_accelerator.v:7129" *)
  wire _T_732;
  (* src = "crypto_accelerator.v:7130" *)
  wire _T_734;
  (* src = "crypto_accelerator.v:7131" *)
  wire _T_736;
  (* src = "crypto_accelerator.v:7132" *)
  wire _T_738;
  (* src = "crypto_accelerator.v:6809" *)
  wire _T_74;
  (* src = "crypto_accelerator.v:7133" *)
  wire _T_740;
  (* src = "crypto_accelerator.v:7134" *)
  wire _T_742;
  (* src = "crypto_accelerator.v:7135" *)
  wire _T_744;
  (* src = "crypto_accelerator.v:7136" *)
  wire _T_746;
  (* src = "crypto_accelerator.v:7137" *)
  wire _T_748;
  (* src = "crypto_accelerator.v:7138" *)
  wire _T_750;
  (* src = "crypto_accelerator.v:7139" *)
  wire _T_752;
  (* src = "crypto_accelerator.v:7140" *)
  wire _T_754;
  (* src = "crypto_accelerator.v:7141" *)
  wire _T_756;
  (* src = "crypto_accelerator.v:7142" *)
  wire _T_758;
  (* src = "crypto_accelerator.v:6810" *)
  wire _T_76;
  (* src = "crypto_accelerator.v:7143" *)
  wire _T_760;
  (* src = "crypto_accelerator.v:7144" *)
  wire _T_762;
  (* src = "crypto_accelerator.v:7145" *)
  wire _T_764;
  (* src = "crypto_accelerator.v:7146" *)
  wire _T_766;
  (* src = "crypto_accelerator.v:7147" *)
  wire _T_768;
  (* src = "crypto_accelerator.v:7148" *)
  wire _T_770;
  (* src = "crypto_accelerator.v:7149" *)
  wire _T_772;
  (* src = "crypto_accelerator.v:7150" *)
  wire _T_774;
  (* src = "crypto_accelerator.v:7151" *)
  wire _T_776;
  (* src = "crypto_accelerator.v:7152" *)
  wire _T_778;
  (* src = "crypto_accelerator.v:6811" *)
  wire _T_78;
  (* src = "crypto_accelerator.v:7153" *)
  wire _T_780;
  (* src = "crypto_accelerator.v:7154" *)
  wire _T_782;
  (* src = "crypto_accelerator.v:7155" *)
  wire _T_784;
  (* src = "crypto_accelerator.v:7156" *)
  wire _T_786;
  (* src = "crypto_accelerator.v:7157" *)
  wire _T_788;
  (* src = "crypto_accelerator.v:7158" *)
  wire _T_790;
  (* src = "crypto_accelerator.v:7159" *)
  wire _T_792;
  (* src = "crypto_accelerator.v:7160" *)
  wire _T_794;
  (* src = "crypto_accelerator.v:7161" *)
  wire _T_796;
  (* src = "crypto_accelerator.v:7162" *)
  wire _T_798;
  (* src = "crypto_accelerator.v:6812" *)
  wire _T_80;
  (* src = "crypto_accelerator.v:7163" *)
  wire _T_800;
  (* src = "crypto_accelerator.v:7164" *)
  wire _T_802;
  (* src = "crypto_accelerator.v:7165" *)
  wire _T_804;
  (* src = "crypto_accelerator.v:7166" *)
  wire _T_806;
  (* src = "crypto_accelerator.v:7167" *)
  wire _T_808;
  (* src = "crypto_accelerator.v:7168" *)
  wire _T_810;
  (* src = "crypto_accelerator.v:7169" *)
  wire _T_812;
  (* src = "crypto_accelerator.v:7170" *)
  wire _T_814;
  (* src = "crypto_accelerator.v:7171" *)
  wire _T_816;
  (* src = "crypto_accelerator.v:7172" *)
  wire _T_818;
  (* src = "crypto_accelerator.v:6813" *)
  wire _T_82;
  (* src = "crypto_accelerator.v:7173" *)
  wire _T_820;
  (* src = "crypto_accelerator.v:7174" *)
  wire _T_822;
  (* src = "crypto_accelerator.v:7175" *)
  wire _T_824;
  (* src = "crypto_accelerator.v:7176" *)
  wire _T_825;
  (* src = "crypto_accelerator.v:7177" *)
  wire _T_826;
  (* src = "crypto_accelerator.v:7178" *)
  wire _T_827;
  (* src = "crypto_accelerator.v:7179" *)
  wire _T_829;
  (* src = "crypto_accelerator.v:7180" *)
  wire _T_830;
  (* src = "crypto_accelerator.v:7181" *)
  wire _T_831;
  (* src = "crypto_accelerator.v:7182" *)
  wire _T_833;
  (* src = "crypto_accelerator.v:7183" *)
  wire _T_835;
  (* src = "crypto_accelerator.v:7184" *)
  wire _T_836;
  (* src = "crypto_accelerator.v:7185" *)
  wire _T_837;
  (* src = "crypto_accelerator.v:7186" *)
  wire _T_839;
  (* src = "crypto_accelerator.v:6814" *)
  wire _T_84;
  (* src = "crypto_accelerator.v:7187" *)
  wire _T_841;
  (* src = "crypto_accelerator.v:7188" *)
  wire _T_843;
  (* src = "crypto_accelerator.v:7189" *)
  wire _T_844;
  (* src = "crypto_accelerator.v:7190" *)
  wire _T_845;
  (* src = "crypto_accelerator.v:7191" *)
  wire _T_847;
  (* src = "crypto_accelerator.v:7192" *)
  wire _T_848;
  (* src = "crypto_accelerator.v:7193" *)
  wire _T_850;
  (* src = "crypto_accelerator.v:7194" *)
  wire _T_851;
  (* src = "crypto_accelerator.v:7195" *)
  wire _T_852;
  (* src = "crypto_accelerator.v:7196" *)
  wire [7:0] _T_859;
  (* src = "crypto_accelerator.v:6815" *)
  wire _T_86;
  (* src = "crypto_accelerator.v:7197" *)
  wire _T_877;
  (* src = "crypto_accelerator.v:7198" *)
  wire _T_879;
  (* src = "crypto_accelerator.v:6816" *)
  wire _T_88;
  (* src = "crypto_accelerator.v:7199" *)
  wire _T_881;
  (* src = "crypto_accelerator.v:7200" *)
  wire _T_883;
  (* src = "crypto_accelerator.v:7201" *)
  wire _T_885;
  (* src = "crypto_accelerator.v:7202" *)
  wire _T_887;
  (* src = "crypto_accelerator.v:7203" *)
  wire _T_889;
  (* src = "crypto_accelerator.v:7204" *)
  wire _T_891;
  (* src = "crypto_accelerator.v:7205" *)
  wire _T_893;
  (* src = "crypto_accelerator.v:7206" *)
  wire _T_895;
  (* src = "crypto_accelerator.v:7207" *)
  wire _T_897;
  (* src = "crypto_accelerator.v:7208" *)
  wire _T_899;
  (* src = "crypto_accelerator.v:6817" *)
  wire _T_90;
  (* src = "crypto_accelerator.v:7209" *)
  wire _T_901;
  (* src = "crypto_accelerator.v:7210" *)
  wire _T_903;
  (* src = "crypto_accelerator.v:7211" *)
  wire _T_905;
  (* src = "crypto_accelerator.v:7212" *)
  wire _T_907;
  (* src = "crypto_accelerator.v:7213" *)
  wire _T_909;
  (* src = "crypto_accelerator.v:7214" *)
  wire _T_911;
  (* src = "crypto_accelerator.v:7215" *)
  wire _T_913;
  (* src = "crypto_accelerator.v:7216" *)
  wire _T_915;
  (* src = "crypto_accelerator.v:7217" *)
  wire _T_917;
  (* src = "crypto_accelerator.v:7218" *)
  wire _T_919;
  (* src = "crypto_accelerator.v:6818" *)
  wire _T_92;
  (* src = "crypto_accelerator.v:7219" *)
  wire _T_921;
  (* src = "crypto_accelerator.v:7220" *)
  wire _T_923;
  (* src = "crypto_accelerator.v:7221" *)
  wire _T_925;
  (* src = "crypto_accelerator.v:7222" *)
  wire _T_927;
  (* src = "crypto_accelerator.v:7223" *)
  wire _T_929;
  (* src = "crypto_accelerator.v:7224" *)
  wire _T_931;
  (* src = "crypto_accelerator.v:7225" *)
  wire _T_933;
  (* src = "crypto_accelerator.v:7226" *)
  wire _T_935;
  (* src = "crypto_accelerator.v:7227" *)
  wire _T_937;
  (* src = "crypto_accelerator.v:7228" *)
  wire _T_939;
  (* src = "crypto_accelerator.v:6819" *)
  wire _T_94;
  (* src = "crypto_accelerator.v:7229" *)
  wire _T_941;
  (* src = "crypto_accelerator.v:7230" *)
  wire _T_943;
  (* src = "crypto_accelerator.v:7231" *)
  wire _T_945;
  (* src = "crypto_accelerator.v:7232" *)
  wire _T_947;
  (* src = "crypto_accelerator.v:7233" *)
  wire _T_949;
  (* src = "crypto_accelerator.v:7234" *)
  wire _T_951;
  (* src = "crypto_accelerator.v:7235" *)
  wire _T_953;
  (* src = "crypto_accelerator.v:7236" *)
  wire _T_955;
  (* src = "crypto_accelerator.v:7237" *)
  wire _T_957;
  (* src = "crypto_accelerator.v:7238" *)
  wire _T_959;
  (* src = "crypto_accelerator.v:6820" *)
  wire _T_96;
  (* src = "crypto_accelerator.v:7239" *)
  wire _T_961;
  (* src = "crypto_accelerator.v:7240" *)
  wire _T_963;
  (* src = "crypto_accelerator.v:7241" *)
  wire _T_965;
  (* src = "crypto_accelerator.v:7242" *)
  wire _T_967;
  (* src = "crypto_accelerator.v:7243" *)
  wire _T_969;
  (* src = "crypto_accelerator.v:7244" *)
  wire _T_971;
  (* src = "crypto_accelerator.v:7245" *)
  wire _T_973;
  (* src = "crypto_accelerator.v:7246" *)
  wire _T_975;
  (* src = "crypto_accelerator.v:7247" *)
  wire _T_977;
  (* src = "crypto_accelerator.v:7248" *)
  wire _T_979;
  (* src = "crypto_accelerator.v:6821" *)
  wire _T_98;
  (* src = "crypto_accelerator.v:7249" *)
  wire _T_981;
  (* src = "crypto_accelerator.v:7250" *)
  wire _T_983;
  (* src = "crypto_accelerator.v:7251" *)
  wire _T_985;
  (* src = "crypto_accelerator.v:7252" *)
  wire _T_987;
  (* src = "crypto_accelerator.v:7253" *)
  wire _T_989;
  (* src = "crypto_accelerator.v:7254" *)
  wire _T_991;
  (* src = "crypto_accelerator.v:7255" *)
  wire _T_993;
  (* src = "crypto_accelerator.v:7256" *)
  wire _T_995;
  (* src = "crypto_accelerator.v:7257" *)
  wire _T_997;
  (* src = "crypto_accelerator.v:7258" *)
  wire _T_999;
  (* src = "crypto_accelerator.v:6469" *)
  input clock;
  (* src = "crypto_accelerator.v:6543" *)
  wire dec_clock;
  (* src = "crypto_accelerator.v:6788" *)
  wire dec_io_aes256;
  (* src = "crypto_accelerator.v:6545" *)
  wire [127:0] dec_io_dataIn;
  (* src = "crypto_accelerator.v:6793" *)
  wire [127:0] dec_io_dataOut;
  (* src = "crypto_accelerator.v:6547" *)
  wire dec_io_dataValid;
  (* src = "crypto_accelerator.v:6546" *)
  wire [127:0] dec_io_ivIn;
  (* src = "crypto_accelerator.v:6794" *)
  wire [127:0] dec_io_ivOut;
  (* src = "crypto_accelerator.v:6548" *)
  wire [7:0] dec_io_keys_0_0_0;
  (* src = "crypto_accelerator.v:6549" *)
  wire [7:0] dec_io_keys_0_0_1;
  (* src = "crypto_accelerator.v:6550" *)
  wire [7:0] dec_io_keys_0_0_2;
  (* src = "crypto_accelerator.v:6551" *)
  wire [7:0] dec_io_keys_0_0_3;
  (* src = "crypto_accelerator.v:6552" *)
  wire [7:0] dec_io_keys_0_1_0;
  (* src = "crypto_accelerator.v:6553" *)
  wire [7:0] dec_io_keys_0_1_1;
  (* src = "crypto_accelerator.v:6554" *)
  wire [7:0] dec_io_keys_0_1_2;
  (* src = "crypto_accelerator.v:6555" *)
  wire [7:0] dec_io_keys_0_1_3;
  (* src = "crypto_accelerator.v:6556" *)
  wire [7:0] dec_io_keys_0_2_0;
  (* src = "crypto_accelerator.v:6557" *)
  wire [7:0] dec_io_keys_0_2_1;
  (* src = "crypto_accelerator.v:6558" *)
  wire [7:0] dec_io_keys_0_2_2;
  (* src = "crypto_accelerator.v:6559" *)
  wire [7:0] dec_io_keys_0_2_3;
  (* src = "crypto_accelerator.v:6560" *)
  wire [7:0] dec_io_keys_0_3_0;
  (* src = "crypto_accelerator.v:6561" *)
  wire [7:0] dec_io_keys_0_3_1;
  (* src = "crypto_accelerator.v:6562" *)
  wire [7:0] dec_io_keys_0_3_2;
  (* src = "crypto_accelerator.v:6563" *)
  wire [7:0] dec_io_keys_0_3_3;
  (* src = "crypto_accelerator.v:6708" *)
  wire [7:0] dec_io_keys_10_0_0;
  (* src = "crypto_accelerator.v:6709" *)
  wire [7:0] dec_io_keys_10_0_1;
  (* src = "crypto_accelerator.v:6710" *)
  wire [7:0] dec_io_keys_10_0_2;
  (* src = "crypto_accelerator.v:6711" *)
  wire [7:0] dec_io_keys_10_0_3;
  (* src = "crypto_accelerator.v:6712" *)
  wire [7:0] dec_io_keys_10_1_0;
  (* src = "crypto_accelerator.v:6713" *)
  wire [7:0] dec_io_keys_10_1_1;
  (* src = "crypto_accelerator.v:6714" *)
  wire [7:0] dec_io_keys_10_1_2;
  (* src = "crypto_accelerator.v:6715" *)
  wire [7:0] dec_io_keys_10_1_3;
  (* src = "crypto_accelerator.v:6716" *)
  wire [7:0] dec_io_keys_10_2_0;
  (* src = "crypto_accelerator.v:6717" *)
  wire [7:0] dec_io_keys_10_2_1;
  (* src = "crypto_accelerator.v:6718" *)
  wire [7:0] dec_io_keys_10_2_2;
  (* src = "crypto_accelerator.v:6719" *)
  wire [7:0] dec_io_keys_10_2_3;
  (* src = "crypto_accelerator.v:6720" *)
  wire [7:0] dec_io_keys_10_3_0;
  (* src = "crypto_accelerator.v:6721" *)
  wire [7:0] dec_io_keys_10_3_1;
  (* src = "crypto_accelerator.v:6722" *)
  wire [7:0] dec_io_keys_10_3_2;
  (* src = "crypto_accelerator.v:6723" *)
  wire [7:0] dec_io_keys_10_3_3;
  (* src = "crypto_accelerator.v:6724" *)
  wire [7:0] dec_io_keys_11_0_0;
  (* src = "crypto_accelerator.v:6725" *)
  wire [7:0] dec_io_keys_11_0_1;
  (* src = "crypto_accelerator.v:6726" *)
  wire [7:0] dec_io_keys_11_0_2;
  (* src = "crypto_accelerator.v:6727" *)
  wire [7:0] dec_io_keys_11_0_3;
  (* src = "crypto_accelerator.v:6728" *)
  wire [7:0] dec_io_keys_11_1_0;
  (* src = "crypto_accelerator.v:6729" *)
  wire [7:0] dec_io_keys_11_1_1;
  (* src = "crypto_accelerator.v:6730" *)
  wire [7:0] dec_io_keys_11_1_2;
  (* src = "crypto_accelerator.v:6731" *)
  wire [7:0] dec_io_keys_11_1_3;
  (* src = "crypto_accelerator.v:6732" *)
  wire [7:0] dec_io_keys_11_2_0;
  (* src = "crypto_accelerator.v:6733" *)
  wire [7:0] dec_io_keys_11_2_1;
  (* src = "crypto_accelerator.v:6734" *)
  wire [7:0] dec_io_keys_11_2_2;
  (* src = "crypto_accelerator.v:6735" *)
  wire [7:0] dec_io_keys_11_2_3;
  (* src = "crypto_accelerator.v:6736" *)
  wire [7:0] dec_io_keys_11_3_0;
  (* src = "crypto_accelerator.v:6737" *)
  wire [7:0] dec_io_keys_11_3_1;
  (* src = "crypto_accelerator.v:6738" *)
  wire [7:0] dec_io_keys_11_3_2;
  (* src = "crypto_accelerator.v:6739" *)
  wire [7:0] dec_io_keys_11_3_3;
  (* src = "crypto_accelerator.v:6740" *)
  wire [7:0] dec_io_keys_12_0_0;
  (* src = "crypto_accelerator.v:6741" *)
  wire [7:0] dec_io_keys_12_0_1;
  (* src = "crypto_accelerator.v:6742" *)
  wire [7:0] dec_io_keys_12_0_2;
  (* src = "crypto_accelerator.v:6743" *)
  wire [7:0] dec_io_keys_12_0_3;
  (* src = "crypto_accelerator.v:6744" *)
  wire [7:0] dec_io_keys_12_1_0;
  (* src = "crypto_accelerator.v:6745" *)
  wire [7:0] dec_io_keys_12_1_1;
  (* src = "crypto_accelerator.v:6746" *)
  wire [7:0] dec_io_keys_12_1_2;
  (* src = "crypto_accelerator.v:6747" *)
  wire [7:0] dec_io_keys_12_1_3;
  (* src = "crypto_accelerator.v:6748" *)
  wire [7:0] dec_io_keys_12_2_0;
  (* src = "crypto_accelerator.v:6749" *)
  wire [7:0] dec_io_keys_12_2_1;
  (* src = "crypto_accelerator.v:6750" *)
  wire [7:0] dec_io_keys_12_2_2;
  (* src = "crypto_accelerator.v:6751" *)
  wire [7:0] dec_io_keys_12_2_3;
  (* src = "crypto_accelerator.v:6752" *)
  wire [7:0] dec_io_keys_12_3_0;
  (* src = "crypto_accelerator.v:6753" *)
  wire [7:0] dec_io_keys_12_3_1;
  (* src = "crypto_accelerator.v:6754" *)
  wire [7:0] dec_io_keys_12_3_2;
  (* src = "crypto_accelerator.v:6755" *)
  wire [7:0] dec_io_keys_12_3_3;
  (* src = "crypto_accelerator.v:6756" *)
  wire [7:0] dec_io_keys_13_0_0;
  (* src = "crypto_accelerator.v:6757" *)
  wire [7:0] dec_io_keys_13_0_1;
  (* src = "crypto_accelerator.v:6758" *)
  wire [7:0] dec_io_keys_13_0_2;
  (* src = "crypto_accelerator.v:6759" *)
  wire [7:0] dec_io_keys_13_0_3;
  (* src = "crypto_accelerator.v:6760" *)
  wire [7:0] dec_io_keys_13_1_0;
  (* src = "crypto_accelerator.v:6761" *)
  wire [7:0] dec_io_keys_13_1_1;
  (* src = "crypto_accelerator.v:6762" *)
  wire [7:0] dec_io_keys_13_1_2;
  (* src = "crypto_accelerator.v:6763" *)
  wire [7:0] dec_io_keys_13_1_3;
  (* src = "crypto_accelerator.v:6764" *)
  wire [7:0] dec_io_keys_13_2_0;
  (* src = "crypto_accelerator.v:6765" *)
  wire [7:0] dec_io_keys_13_2_1;
  (* src = "crypto_accelerator.v:6766" *)
  wire [7:0] dec_io_keys_13_2_2;
  (* src = "crypto_accelerator.v:6767" *)
  wire [7:0] dec_io_keys_13_2_3;
  (* src = "crypto_accelerator.v:6768" *)
  wire [7:0] dec_io_keys_13_3_0;
  (* src = "crypto_accelerator.v:6769" *)
  wire [7:0] dec_io_keys_13_3_1;
  (* src = "crypto_accelerator.v:6770" *)
  wire [7:0] dec_io_keys_13_3_2;
  (* src = "crypto_accelerator.v:6771" *)
  wire [7:0] dec_io_keys_13_3_3;
  (* src = "crypto_accelerator.v:6772" *)
  wire [7:0] dec_io_keys_14_0_0;
  (* src = "crypto_accelerator.v:6773" *)
  wire [7:0] dec_io_keys_14_0_1;
  (* src = "crypto_accelerator.v:6774" *)
  wire [7:0] dec_io_keys_14_0_2;
  (* src = "crypto_accelerator.v:6775" *)
  wire [7:0] dec_io_keys_14_0_3;
  (* src = "crypto_accelerator.v:6776" *)
  wire [7:0] dec_io_keys_14_1_0;
  (* src = "crypto_accelerator.v:6777" *)
  wire [7:0] dec_io_keys_14_1_1;
  (* src = "crypto_accelerator.v:6778" *)
  wire [7:0] dec_io_keys_14_1_2;
  (* src = "crypto_accelerator.v:6779" *)
  wire [7:0] dec_io_keys_14_1_3;
  (* src = "crypto_accelerator.v:6780" *)
  wire [7:0] dec_io_keys_14_2_0;
  (* src = "crypto_accelerator.v:6781" *)
  wire [7:0] dec_io_keys_14_2_1;
  (* src = "crypto_accelerator.v:6782" *)
  wire [7:0] dec_io_keys_14_2_2;
  (* src = "crypto_accelerator.v:6783" *)
  wire [7:0] dec_io_keys_14_2_3;
  (* src = "crypto_accelerator.v:6784" *)
  wire [7:0] dec_io_keys_14_3_0;
  (* src = "crypto_accelerator.v:6785" *)
  wire [7:0] dec_io_keys_14_3_1;
  (* src = "crypto_accelerator.v:6786" *)
  wire [7:0] dec_io_keys_14_3_2;
  (* src = "crypto_accelerator.v:6787" *)
  wire [7:0] dec_io_keys_14_3_3;
  (* src = "crypto_accelerator.v:6564" *)
  wire [7:0] dec_io_keys_1_0_0;
  (* src = "crypto_accelerator.v:6565" *)
  wire [7:0] dec_io_keys_1_0_1;
  (* src = "crypto_accelerator.v:6566" *)
  wire [7:0] dec_io_keys_1_0_2;
  (* src = "crypto_accelerator.v:6567" *)
  wire [7:0] dec_io_keys_1_0_3;
  (* src = "crypto_accelerator.v:6568" *)
  wire [7:0] dec_io_keys_1_1_0;
  (* src = "crypto_accelerator.v:6569" *)
  wire [7:0] dec_io_keys_1_1_1;
  (* src = "crypto_accelerator.v:6570" *)
  wire [7:0] dec_io_keys_1_1_2;
  (* src = "crypto_accelerator.v:6571" *)
  wire [7:0] dec_io_keys_1_1_3;
  (* src = "crypto_accelerator.v:6572" *)
  wire [7:0] dec_io_keys_1_2_0;
  (* src = "crypto_accelerator.v:6573" *)
  wire [7:0] dec_io_keys_1_2_1;
  (* src = "crypto_accelerator.v:6574" *)
  wire [7:0] dec_io_keys_1_2_2;
  (* src = "crypto_accelerator.v:6575" *)
  wire [7:0] dec_io_keys_1_2_3;
  (* src = "crypto_accelerator.v:6576" *)
  wire [7:0] dec_io_keys_1_3_0;
  (* src = "crypto_accelerator.v:6577" *)
  wire [7:0] dec_io_keys_1_3_1;
  (* src = "crypto_accelerator.v:6578" *)
  wire [7:0] dec_io_keys_1_3_2;
  (* src = "crypto_accelerator.v:6579" *)
  wire [7:0] dec_io_keys_1_3_3;
  (* src = "crypto_accelerator.v:6580" *)
  wire [7:0] dec_io_keys_2_0_0;
  (* src = "crypto_accelerator.v:6581" *)
  wire [7:0] dec_io_keys_2_0_1;
  (* src = "crypto_accelerator.v:6582" *)
  wire [7:0] dec_io_keys_2_0_2;
  (* src = "crypto_accelerator.v:6583" *)
  wire [7:0] dec_io_keys_2_0_3;
  (* src = "crypto_accelerator.v:6584" *)
  wire [7:0] dec_io_keys_2_1_0;
  (* src = "crypto_accelerator.v:6585" *)
  wire [7:0] dec_io_keys_2_1_1;
  (* src = "crypto_accelerator.v:6586" *)
  wire [7:0] dec_io_keys_2_1_2;
  (* src = "crypto_accelerator.v:6587" *)
  wire [7:0] dec_io_keys_2_1_3;
  (* src = "crypto_accelerator.v:6588" *)
  wire [7:0] dec_io_keys_2_2_0;
  (* src = "crypto_accelerator.v:6589" *)
  wire [7:0] dec_io_keys_2_2_1;
  (* src = "crypto_accelerator.v:6590" *)
  wire [7:0] dec_io_keys_2_2_2;
  (* src = "crypto_accelerator.v:6591" *)
  wire [7:0] dec_io_keys_2_2_3;
  (* src = "crypto_accelerator.v:6592" *)
  wire [7:0] dec_io_keys_2_3_0;
  (* src = "crypto_accelerator.v:6593" *)
  wire [7:0] dec_io_keys_2_3_1;
  (* src = "crypto_accelerator.v:6594" *)
  wire [7:0] dec_io_keys_2_3_2;
  (* src = "crypto_accelerator.v:6595" *)
  wire [7:0] dec_io_keys_2_3_3;
  (* src = "crypto_accelerator.v:6596" *)
  wire [7:0] dec_io_keys_3_0_0;
  (* src = "crypto_accelerator.v:6597" *)
  wire [7:0] dec_io_keys_3_0_1;
  (* src = "crypto_accelerator.v:6598" *)
  wire [7:0] dec_io_keys_3_0_2;
  (* src = "crypto_accelerator.v:6599" *)
  wire [7:0] dec_io_keys_3_0_3;
  (* src = "crypto_accelerator.v:6600" *)
  wire [7:0] dec_io_keys_3_1_0;
  (* src = "crypto_accelerator.v:6601" *)
  wire [7:0] dec_io_keys_3_1_1;
  (* src = "crypto_accelerator.v:6602" *)
  wire [7:0] dec_io_keys_3_1_2;
  (* src = "crypto_accelerator.v:6603" *)
  wire [7:0] dec_io_keys_3_1_3;
  (* src = "crypto_accelerator.v:6604" *)
  wire [7:0] dec_io_keys_3_2_0;
  (* src = "crypto_accelerator.v:6605" *)
  wire [7:0] dec_io_keys_3_2_1;
  (* src = "crypto_accelerator.v:6606" *)
  wire [7:0] dec_io_keys_3_2_2;
  (* src = "crypto_accelerator.v:6607" *)
  wire [7:0] dec_io_keys_3_2_3;
  (* src = "crypto_accelerator.v:6608" *)
  wire [7:0] dec_io_keys_3_3_0;
  (* src = "crypto_accelerator.v:6609" *)
  wire [7:0] dec_io_keys_3_3_1;
  (* src = "crypto_accelerator.v:6610" *)
  wire [7:0] dec_io_keys_3_3_2;
  (* src = "crypto_accelerator.v:6611" *)
  wire [7:0] dec_io_keys_3_3_3;
  (* src = "crypto_accelerator.v:6612" *)
  wire [7:0] dec_io_keys_4_0_0;
  (* src = "crypto_accelerator.v:6613" *)
  wire [7:0] dec_io_keys_4_0_1;
  (* src = "crypto_accelerator.v:6614" *)
  wire [7:0] dec_io_keys_4_0_2;
  (* src = "crypto_accelerator.v:6615" *)
  wire [7:0] dec_io_keys_4_0_3;
  (* src = "crypto_accelerator.v:6616" *)
  wire [7:0] dec_io_keys_4_1_0;
  (* src = "crypto_accelerator.v:6617" *)
  wire [7:0] dec_io_keys_4_1_1;
  (* src = "crypto_accelerator.v:6618" *)
  wire [7:0] dec_io_keys_4_1_2;
  (* src = "crypto_accelerator.v:6619" *)
  wire [7:0] dec_io_keys_4_1_3;
  (* src = "crypto_accelerator.v:6620" *)
  wire [7:0] dec_io_keys_4_2_0;
  (* src = "crypto_accelerator.v:6621" *)
  wire [7:0] dec_io_keys_4_2_1;
  (* src = "crypto_accelerator.v:6622" *)
  wire [7:0] dec_io_keys_4_2_2;
  (* src = "crypto_accelerator.v:6623" *)
  wire [7:0] dec_io_keys_4_2_3;
  (* src = "crypto_accelerator.v:6624" *)
  wire [7:0] dec_io_keys_4_3_0;
  (* src = "crypto_accelerator.v:6625" *)
  wire [7:0] dec_io_keys_4_3_1;
  (* src = "crypto_accelerator.v:6626" *)
  wire [7:0] dec_io_keys_4_3_2;
  (* src = "crypto_accelerator.v:6627" *)
  wire [7:0] dec_io_keys_4_3_3;
  (* src = "crypto_accelerator.v:6628" *)
  wire [7:0] dec_io_keys_5_0_0;
  (* src = "crypto_accelerator.v:6629" *)
  wire [7:0] dec_io_keys_5_0_1;
  (* src = "crypto_accelerator.v:6630" *)
  wire [7:0] dec_io_keys_5_0_2;
  (* src = "crypto_accelerator.v:6631" *)
  wire [7:0] dec_io_keys_5_0_3;
  (* src = "crypto_accelerator.v:6632" *)
  wire [7:0] dec_io_keys_5_1_0;
  (* src = "crypto_accelerator.v:6633" *)
  wire [7:0] dec_io_keys_5_1_1;
  (* src = "crypto_accelerator.v:6634" *)
  wire [7:0] dec_io_keys_5_1_2;
  (* src = "crypto_accelerator.v:6635" *)
  wire [7:0] dec_io_keys_5_1_3;
  (* src = "crypto_accelerator.v:6636" *)
  wire [7:0] dec_io_keys_5_2_0;
  (* src = "crypto_accelerator.v:6637" *)
  wire [7:0] dec_io_keys_5_2_1;
  (* src = "crypto_accelerator.v:6638" *)
  wire [7:0] dec_io_keys_5_2_2;
  (* src = "crypto_accelerator.v:6639" *)
  wire [7:0] dec_io_keys_5_2_3;
  (* src = "crypto_accelerator.v:6640" *)
  wire [7:0] dec_io_keys_5_3_0;
  (* src = "crypto_accelerator.v:6641" *)
  wire [7:0] dec_io_keys_5_3_1;
  (* src = "crypto_accelerator.v:6642" *)
  wire [7:0] dec_io_keys_5_3_2;
  (* src = "crypto_accelerator.v:6643" *)
  wire [7:0] dec_io_keys_5_3_3;
  (* src = "crypto_accelerator.v:6644" *)
  wire [7:0] dec_io_keys_6_0_0;
  (* src = "crypto_accelerator.v:6645" *)
  wire [7:0] dec_io_keys_6_0_1;
  (* src = "crypto_accelerator.v:6646" *)
  wire [7:0] dec_io_keys_6_0_2;
  (* src = "crypto_accelerator.v:6647" *)
  wire [7:0] dec_io_keys_6_0_3;
  (* src = "crypto_accelerator.v:6648" *)
  wire [7:0] dec_io_keys_6_1_0;
  (* src = "crypto_accelerator.v:6649" *)
  wire [7:0] dec_io_keys_6_1_1;
  (* src = "crypto_accelerator.v:6650" *)
  wire [7:0] dec_io_keys_6_1_2;
  (* src = "crypto_accelerator.v:6651" *)
  wire [7:0] dec_io_keys_6_1_3;
  (* src = "crypto_accelerator.v:6652" *)
  wire [7:0] dec_io_keys_6_2_0;
  (* src = "crypto_accelerator.v:6653" *)
  wire [7:0] dec_io_keys_6_2_1;
  (* src = "crypto_accelerator.v:6654" *)
  wire [7:0] dec_io_keys_6_2_2;
  (* src = "crypto_accelerator.v:6655" *)
  wire [7:0] dec_io_keys_6_2_3;
  (* src = "crypto_accelerator.v:6656" *)
  wire [7:0] dec_io_keys_6_3_0;
  (* src = "crypto_accelerator.v:6657" *)
  wire [7:0] dec_io_keys_6_3_1;
  (* src = "crypto_accelerator.v:6658" *)
  wire [7:0] dec_io_keys_6_3_2;
  (* src = "crypto_accelerator.v:6659" *)
  wire [7:0] dec_io_keys_6_3_3;
  (* src = "crypto_accelerator.v:6660" *)
  wire [7:0] dec_io_keys_7_0_0;
  (* src = "crypto_accelerator.v:6661" *)
  wire [7:0] dec_io_keys_7_0_1;
  (* src = "crypto_accelerator.v:6662" *)
  wire [7:0] dec_io_keys_7_0_2;
  (* src = "crypto_accelerator.v:6663" *)
  wire [7:0] dec_io_keys_7_0_3;
  (* src = "crypto_accelerator.v:6664" *)
  wire [7:0] dec_io_keys_7_1_0;
  (* src = "crypto_accelerator.v:6665" *)
  wire [7:0] dec_io_keys_7_1_1;
  (* src = "crypto_accelerator.v:6666" *)
  wire [7:0] dec_io_keys_7_1_2;
  (* src = "crypto_accelerator.v:6667" *)
  wire [7:0] dec_io_keys_7_1_3;
  (* src = "crypto_accelerator.v:6668" *)
  wire [7:0] dec_io_keys_7_2_0;
  (* src = "crypto_accelerator.v:6669" *)
  wire [7:0] dec_io_keys_7_2_1;
  (* src = "crypto_accelerator.v:6670" *)
  wire [7:0] dec_io_keys_7_2_2;
  (* src = "crypto_accelerator.v:6671" *)
  wire [7:0] dec_io_keys_7_2_3;
  (* src = "crypto_accelerator.v:6672" *)
  wire [7:0] dec_io_keys_7_3_0;
  (* src = "crypto_accelerator.v:6673" *)
  wire [7:0] dec_io_keys_7_3_1;
  (* src = "crypto_accelerator.v:6674" *)
  wire [7:0] dec_io_keys_7_3_2;
  (* src = "crypto_accelerator.v:6675" *)
  wire [7:0] dec_io_keys_7_3_3;
  (* src = "crypto_accelerator.v:6676" *)
  wire [7:0] dec_io_keys_8_0_0;
  (* src = "crypto_accelerator.v:6677" *)
  wire [7:0] dec_io_keys_8_0_1;
  (* src = "crypto_accelerator.v:6678" *)
  wire [7:0] dec_io_keys_8_0_2;
  (* src = "crypto_accelerator.v:6679" *)
  wire [7:0] dec_io_keys_8_0_3;
  (* src = "crypto_accelerator.v:6680" *)
  wire [7:0] dec_io_keys_8_1_0;
  (* src = "crypto_accelerator.v:6681" *)
  wire [7:0] dec_io_keys_8_1_1;
  (* src = "crypto_accelerator.v:6682" *)
  wire [7:0] dec_io_keys_8_1_2;
  (* src = "crypto_accelerator.v:6683" *)
  wire [7:0] dec_io_keys_8_1_3;
  (* src = "crypto_accelerator.v:6684" *)
  wire [7:0] dec_io_keys_8_2_0;
  (* src = "crypto_accelerator.v:6685" *)
  wire [7:0] dec_io_keys_8_2_1;
  (* src = "crypto_accelerator.v:6686" *)
  wire [7:0] dec_io_keys_8_2_2;
  (* src = "crypto_accelerator.v:6687" *)
  wire [7:0] dec_io_keys_8_2_3;
  (* src = "crypto_accelerator.v:6688" *)
  wire [7:0] dec_io_keys_8_3_0;
  (* src = "crypto_accelerator.v:6689" *)
  wire [7:0] dec_io_keys_8_3_1;
  (* src = "crypto_accelerator.v:6690" *)
  wire [7:0] dec_io_keys_8_3_2;
  (* src = "crypto_accelerator.v:6691" *)
  wire [7:0] dec_io_keys_8_3_3;
  (* src = "crypto_accelerator.v:6692" *)
  wire [7:0] dec_io_keys_9_0_0;
  (* src = "crypto_accelerator.v:6693" *)
  wire [7:0] dec_io_keys_9_0_1;
  (* src = "crypto_accelerator.v:6694" *)
  wire [7:0] dec_io_keys_9_0_2;
  (* src = "crypto_accelerator.v:6695" *)
  wire [7:0] dec_io_keys_9_0_3;
  (* src = "crypto_accelerator.v:6696" *)
  wire [7:0] dec_io_keys_9_1_0;
  (* src = "crypto_accelerator.v:6697" *)
  wire [7:0] dec_io_keys_9_1_1;
  (* src = "crypto_accelerator.v:6698" *)
  wire [7:0] dec_io_keys_9_1_2;
  (* src = "crypto_accelerator.v:6699" *)
  wire [7:0] dec_io_keys_9_1_3;
  (* src = "crypto_accelerator.v:6700" *)
  wire [7:0] dec_io_keys_9_2_0;
  (* src = "crypto_accelerator.v:6701" *)
  wire [7:0] dec_io_keys_9_2_1;
  (* src = "crypto_accelerator.v:6702" *)
  wire [7:0] dec_io_keys_9_2_2;
  (* src = "crypto_accelerator.v:6703" *)
  wire [7:0] dec_io_keys_9_2_3;
  (* src = "crypto_accelerator.v:6704" *)
  wire [7:0] dec_io_keys_9_3_0;
  (* src = "crypto_accelerator.v:6705" *)
  wire [7:0] dec_io_keys_9_3_1;
  (* src = "crypto_accelerator.v:6706" *)
  wire [7:0] dec_io_keys_9_3_2;
  (* src = "crypto_accelerator.v:6707" *)
  wire [7:0] dec_io_keys_9_3_3;
  (* src = "crypto_accelerator.v:6795" *)
  wire dec_io_outputValid;
  (* src = "crypto_accelerator.v:6792" *)
  wire dec_io_ready;
  (* src = "crypto_accelerator.v:6791" *)
  wire dec_io_shift;
  (* src = "crypto_accelerator.v:6789" *)
  wire dec_io_shiftCyc;
  (* src = "crypto_accelerator.v:6790" *)
  wire dec_io_shiftRev;
  (* src = "crypto_accelerator.v:6544" *)
  wire dec_reset;
  (* src = "crypto_accelerator.v:6515" *)
  wire enc_clock;
  (* src = "crypto_accelerator.v:6536" *)
  wire enc_io_aes256;
  (* src = "crypto_accelerator.v:6517" *)
  wire [127:0] enc_io_dataIn;
  (* src = "crypto_accelerator.v:6540" *)
  wire [127:0] enc_io_dataOut;
  (* src = "crypto_accelerator.v:6519" *)
  wire enc_io_dataValid;
  (* src = "crypto_accelerator.v:6518" *)
  wire [127:0] enc_io_ivIn;
  (* src = "crypto_accelerator.v:6541" *)
  wire [127:0] enc_io_ivOut;
  (* src = "crypto_accelerator.v:6520" *)
  wire [7:0] enc_io_keys_0_0_0;
  (* src = "crypto_accelerator.v:6521" *)
  wire [7:0] enc_io_keys_0_0_1;
  (* src = "crypto_accelerator.v:6522" *)
  wire [7:0] enc_io_keys_0_0_2;
  (* src = "crypto_accelerator.v:6523" *)
  wire [7:0] enc_io_keys_0_0_3;
  (* src = "crypto_accelerator.v:6524" *)
  wire [7:0] enc_io_keys_0_1_0;
  (* src = "crypto_accelerator.v:6525" *)
  wire [7:0] enc_io_keys_0_1_1;
  (* src = "crypto_accelerator.v:6526" *)
  wire [7:0] enc_io_keys_0_1_2;
  (* src = "crypto_accelerator.v:6527" *)
  wire [7:0] enc_io_keys_0_1_3;
  (* src = "crypto_accelerator.v:6528" *)
  wire [7:0] enc_io_keys_0_2_0;
  (* src = "crypto_accelerator.v:6529" *)
  wire [7:0] enc_io_keys_0_2_1;
  (* src = "crypto_accelerator.v:6530" *)
  wire [7:0] enc_io_keys_0_2_2;
  (* src = "crypto_accelerator.v:6531" *)
  wire [7:0] enc_io_keys_0_2_3;
  (* src = "crypto_accelerator.v:6532" *)
  wire [7:0] enc_io_keys_0_3_0;
  (* src = "crypto_accelerator.v:6533" *)
  wire [7:0] enc_io_keys_0_3_1;
  (* src = "crypto_accelerator.v:6534" *)
  wire [7:0] enc_io_keys_0_3_2;
  (* src = "crypto_accelerator.v:6535" *)
  wire [7:0] enc_io_keys_0_3_3;
  (* src = "crypto_accelerator.v:6542" *)
  wire enc_io_outputValid;
  (* src = "crypto_accelerator.v:6539" *)
  wire enc_io_ready;
  (* src = "crypto_accelerator.v:6538" *)
  wire enc_io_shift;
  (* src = "crypto_accelerator.v:6537" *)
  wire enc_io_shiftCyc;
  (* src = "crypto_accelerator.v:6516" *)
  wire enc_reset;
  (* src = "crypto_accelerator.v:6477" *)
  input io_aes256;
  (* src = "crypto_accelerator.v:6474" *)
  input [127:0] io_decDataIn;
  (* src = "crypto_accelerator.v:6486" *)
  output [127:0] io_decDataOut;
  (* src = "crypto_accelerator.v:6476" *)
  input io_decDataValid;
  (* src = "crypto_accelerator.v:6475" *)
  input [127:0] io_decIvIn;
  (* src = "crypto_accelerator.v:6487" *)
  output [127:0] io_decIvOut;
  (* src = "crypto_accelerator.v:6488" *)
  output io_decOutputValid;
  (* src = "crypto_accelerator.v:6482" *)
  output io_decReady;
  (* src = "crypto_accelerator.v:6471" *)
  input [127:0] io_encDataIn;
  (* src = "crypto_accelerator.v:6483" *)
  output [127:0] io_encDataOut;
  (* src = "crypto_accelerator.v:6473" *)
  input io_encDataValid;
  (* src = "crypto_accelerator.v:6472" *)
  input [127:0] io_encIvIn;
  (* src = "crypto_accelerator.v:6484" *)
  output [127:0] io_encIvOut;
  (* src = "crypto_accelerator.v:6485" *)
  output io_encOutputValid;
  (* src = "crypto_accelerator.v:6481" *)
  output io_encReady;
  (* src = "crypto_accelerator.v:6478" *)
  input [127:0] io_keyIn;
  (* src = "crypto_accelerator.v:6479" *)
  input io_keyShift;
  (* src = "crypto_accelerator.v:6480" *)
  input io_keyValid;
  (* src = "crypto_accelerator.v:6797" *)
  reg [5:0] keyInd;
  (* src = "crypto_accelerator.v:6796" *)
  reg keyUpdate;
  (* src = "crypto_accelerator.v:6470" *)
  input reset;
  (* src = "crypto_accelerator.v:6494" *)
  wire shreg_clock;
  (* src = "crypto_accelerator.v:6498" *)
  wire shreg_io_cyc;
  (* src = "crypto_accelerator.v:6496" *)
  wire shreg_io_enable;
  (* src = "crypto_accelerator.v:6495" *)
  wire [127:0] shreg_io_input;
  (* src = "crypto_accelerator.v:6500" *)
  wire [127:0] shreg_io_output_0;
  (* src = "crypto_accelerator.v:6501" *)
  wire [127:0] shreg_io_output_1;
  (* src = "crypto_accelerator.v:6510" *)
  wire [127:0] shreg_io_output_10;
  (* src = "crypto_accelerator.v:6511" *)
  wire [127:0] shreg_io_output_11;
  (* src = "crypto_accelerator.v:6512" *)
  wire [127:0] shreg_io_output_12;
  (* src = "crypto_accelerator.v:6513" *)
  wire [127:0] shreg_io_output_13;
  (* src = "crypto_accelerator.v:6514" *)
  wire [127:0] shreg_io_output_14;
  (* src = "crypto_accelerator.v:6502" *)
  wire [127:0] shreg_io_output_2;
  (* src = "crypto_accelerator.v:6503" *)
  wire [127:0] shreg_io_output_3;
  (* src = "crypto_accelerator.v:6504" *)
  wire [127:0] shreg_io_output_4;
  (* src = "crypto_accelerator.v:6505" *)
  wire [127:0] shreg_io_output_5;
  (* src = "crypto_accelerator.v:6506" *)
  wire [127:0] shreg_io_output_6;
  (* src = "crypto_accelerator.v:6507" *)
  wire [127:0] shreg_io_output_7;
  (* src = "crypto_accelerator.v:6508" *)
  wire [127:0] shreg_io_output_8;
  (* src = "crypto_accelerator.v:6509" *)
  wire [127:0] shreg_io_output_9;
  (* src = "crypto_accelerator.v:6497" *)
  wire shreg_io_rev;
  (* src = "crypto_accelerator.v:6499" *)
  wire shreg_io_tap;
  assign _T_2 = keyInd + (* src = "crypto_accelerator.v:6801" *) 1'b1;
  assign _T_1133 = keyInd[4:1] + (* src = "crypto_accelerator.v:7343" *) 1'b1;
  assign _T_52 = _T_51 & (* src = "crypto_accelerator.v:6806" *) io_aes256;
  assign _T_124 = _T_106 & (* src = "crypto_accelerator.v:6834" *) _T_78;
  assign _T_126 = _T_108 & (* src = "crypto_accelerator.v:6835" *) _T_90;
  assign _T_130 = _T_88 & (* src = "crypto_accelerator.v:6837" *) shreg_io_output_0[24];
  assign _T_134 = _T_82 & (* src = "crypto_accelerator.v:6839" *) _T_110;
  assign _T_136 = _T_86 & (* src = "crypto_accelerator.v:6840" *) _T_76;
  assign _T_140 = _T_112 & (* src = "crypto_accelerator.v:6842" *) _T_102;
  assign _T_144 = _T_72 & (* src = "crypto_accelerator.v:6844" *) _T_84;
  assign _T_146 = _T_118 & (* src = "crypto_accelerator.v:6845" *) _T_114;
  assign _T_150 = _T_100 & (* src = "crypto_accelerator.v:6847" *) _T_96;
  assign _T_172 = _T_166 & (* src = "crypto_accelerator.v:6858" *) _T_162;
  assign _T_180 = _T_178 & (* src = "crypto_accelerator.v:6862" *) _T_176;
  assign _T_182 = _T_174 & (* src = "crypto_accelerator.v:6863" *) _T_170;
  assign _T_184 = _T_162 & (* src = "crypto_accelerator.v:6864" *) _T_168;
  assign _T_186 = _T_176 & (* src = "crypto_accelerator.v:6865" *) _T_184;
  assign _T_190 = _T_164 & (* src = "crypto_accelerator.v:6867" *) _T_166;
  assign _T_192 = _T_170 & (* src = "crypto_accelerator.v:6868" *) _T_190;
  assign _T_214 = _T_210 & (* src = "crypto_accelerator.v:6879" *) _T_78;
  assign _T_216 = _T_202 & (* src = "crypto_accelerator.v:6880" *) _T_90;
  assign _T_218 = _T_200 & (* src = "crypto_accelerator.v:6881" *) shreg_io_output_0[24];
  assign _T_220 = _T_208 & (* src = "crypto_accelerator.v:6882" *) _T_110;
  assign _T_222 = _T_198 & (* src = "crypto_accelerator.v:6883" *) _T_76;
  assign _T_224 = _T_196 & (* src = "crypto_accelerator.v:6884" *) _T_102;
  assign _T_226 = _T_206 & (* src = "crypto_accelerator.v:6885" *) _T_84;
  assign _T_228 = _T_212 & (* src = "crypto_accelerator.v:6886" *) _T_114;
  assign _T_230 = _T_204 & (* src = "crypto_accelerator.v:6887" *) _T_96;
  assign _T_232 = _T_210 & (* src = "crypto_accelerator.v:6888" *) _T_106;
  assign _T_234 = _T_202 & (* src = "crypto_accelerator.v:6889" *) _T_108;
  assign _T_236 = _T_200 & (* src = "crypto_accelerator.v:6890" *) _T_88;
  assign _T_238 = _T_208 & (* src = "crypto_accelerator.v:6891" *) _T_82;
  assign _T_240 = _T_198 & (* src = "crypto_accelerator.v:6892" *) _T_86;
  assign _T_242 = _T_196 & (* src = "crypto_accelerator.v:6893" *) _T_112;
  assign _T_244 = _T_206 & (* src = "crypto_accelerator.v:6894" *) _T_72;
  assign _T_246 = _T_212 & (* src = "crypto_accelerator.v:6895" *) _T_118;
  assign _T_248 = _T_204 & (* src = "crypto_accelerator.v:6896" *) _T_100;
  assign _T_393 = _T_375 & (* src = "crypto_accelerator.v:6964" *) _T_347;
  assign _T_395 = _T_377 & (* src = "crypto_accelerator.v:6965" *) _T_359;
  assign _T_399 = _T_357 & (* src = "crypto_accelerator.v:6967" *) shreg_io_output_0[16];
  assign _T_403 = _T_351 & (* src = "crypto_accelerator.v:6969" *) _T_379;
  assign _T_405 = _T_355 & (* src = "crypto_accelerator.v:6970" *) _T_345;
  assign _T_409 = _T_381 & (* src = "crypto_accelerator.v:6972" *) _T_371;
  assign _T_413 = _T_341 & (* src = "crypto_accelerator.v:6974" *) _T_353;
  assign _T_415 = _T_387 & (* src = "crypto_accelerator.v:6975" *) _T_383;
  assign _T_419 = _T_369 & (* src = "crypto_accelerator.v:6977" *) _T_365;
  assign _T_441 = _T_435 & (* src = "crypto_accelerator.v:6988" *) _T_431;
  assign _T_449 = _T_447 & (* src = "crypto_accelerator.v:6992" *) _T_445;
  assign _T_451 = _T_443 & (* src = "crypto_accelerator.v:6993" *) _T_439;
  assign _T_453 = _T_431 & (* src = "crypto_accelerator.v:6994" *) _T_437;
  assign _T_455 = _T_445 & (* src = "crypto_accelerator.v:6995" *) _T_453;
  assign _T_459 = _T_433 & (* src = "crypto_accelerator.v:6997" *) _T_435;
  assign _T_461 = _T_439 & (* src = "crypto_accelerator.v:6998" *) _T_459;
  assign _T_483 = _T_479 & (* src = "crypto_accelerator.v:7009" *) _T_347;
  assign _T_485 = _T_471 & (* src = "crypto_accelerator.v:7010" *) _T_359;
  assign _T_487 = _T_469 & (* src = "crypto_accelerator.v:7011" *) shreg_io_output_0[16];
  assign _T_489 = _T_477 & (* src = "crypto_accelerator.v:7012" *) _T_379;
  assign _T_491 = _T_467 & (* src = "crypto_accelerator.v:7013" *) _T_345;
  assign _T_493 = _T_465 & (* src = "crypto_accelerator.v:7014" *) _T_371;
  assign _T_495 = _T_475 & (* src = "crypto_accelerator.v:7015" *) _T_353;
  assign _T_497 = _T_481 & (* src = "crypto_accelerator.v:7016" *) _T_383;
  assign _T_499 = _T_473 & (* src = "crypto_accelerator.v:7017" *) _T_365;
  assign _T_501 = _T_479 & (* src = "crypto_accelerator.v:7018" *) _T_375;
  assign _T_503 = _T_471 & (* src = "crypto_accelerator.v:7019" *) _T_377;
  assign _T_505 = _T_469 & (* src = "crypto_accelerator.v:7020" *) _T_357;
  assign _T_507 = _T_477 & (* src = "crypto_accelerator.v:7021" *) _T_351;
  assign _T_509 = _T_467 & (* src = "crypto_accelerator.v:7022" *) _T_355;
  assign _T_511 = _T_465 & (* src = "crypto_accelerator.v:7023" *) _T_381;
  assign _T_513 = _T_475 & (* src = "crypto_accelerator.v:7024" *) _T_341;
  assign _T_515 = _T_481 & (* src = "crypto_accelerator.v:7025" *) _T_387;
  assign _T_517 = _T_473 & (* src = "crypto_accelerator.v:7026" *) _T_369;
  assign _T_662 = _T_644 & (* src = "crypto_accelerator.v:7094" *) _T_616;
  assign _T_664 = _T_646 & (* src = "crypto_accelerator.v:7095" *) _T_628;
  assign _T_668 = _T_626 & (* src = "crypto_accelerator.v:7097" *) shreg_io_output_0[8];
  assign _T_672 = _T_620 & (* src = "crypto_accelerator.v:7099" *) _T_648;
  assign _T_674 = _T_624 & (* src = "crypto_accelerator.v:7100" *) _T_614;
  assign _T_678 = _T_650 & (* src = "crypto_accelerator.v:7102" *) _T_640;
  assign _T_682 = _T_610 & (* src = "crypto_accelerator.v:7104" *) _T_622;
  assign _T_684 = _T_656 & (* src = "crypto_accelerator.v:7105" *) _T_652;
  assign _T_688 = _T_638 & (* src = "crypto_accelerator.v:7107" *) _T_634;
  assign _T_710 = _T_704 & (* src = "crypto_accelerator.v:7118" *) _T_700;
  assign _T_718 = _T_716 & (* src = "crypto_accelerator.v:7122" *) _T_714;
  assign _T_720 = _T_712 & (* src = "crypto_accelerator.v:7123" *) _T_708;
  assign _T_722 = _T_700 & (* src = "crypto_accelerator.v:7124" *) _T_706;
  assign _T_724 = _T_714 & (* src = "crypto_accelerator.v:7125" *) _T_722;
  assign _T_728 = _T_702 & (* src = "crypto_accelerator.v:7127" *) _T_704;
  assign _T_730 = _T_708 & (* src = "crypto_accelerator.v:7128" *) _T_728;
  assign _T_752 = _T_748 & (* src = "crypto_accelerator.v:7139" *) _T_616;
  assign _T_754 = _T_740 & (* src = "crypto_accelerator.v:7140" *) _T_628;
  assign _T_756 = _T_738 & (* src = "crypto_accelerator.v:7141" *) shreg_io_output_0[8];
  assign _T_758 = _T_746 & (* src = "crypto_accelerator.v:7142" *) _T_648;
  assign _T_760 = _T_736 & (* src = "crypto_accelerator.v:7143" *) _T_614;
  assign _T_762 = _T_734 & (* src = "crypto_accelerator.v:7144" *) _T_640;
  assign _T_764 = _T_744 & (* src = "crypto_accelerator.v:7145" *) _T_622;
  assign _T_766 = _T_750 & (* src = "crypto_accelerator.v:7146" *) _T_652;
  assign _T_768 = _T_742 & (* src = "crypto_accelerator.v:7147" *) _T_634;
  assign _T_770 = _T_748 & (* src = "crypto_accelerator.v:7148" *) _T_644;
  assign _T_772 = _T_740 & (* src = "crypto_accelerator.v:7149" *) _T_646;
  assign _T_774 = _T_738 & (* src = "crypto_accelerator.v:7150" *) _T_626;
  assign _T_776 = _T_746 & (* src = "crypto_accelerator.v:7151" *) _T_620;
  assign _T_778 = _T_736 & (* src = "crypto_accelerator.v:7152" *) _T_624;
  assign _T_780 = _T_734 & (* src = "crypto_accelerator.v:7153" *) _T_650;
  assign _T_782 = _T_744 & (* src = "crypto_accelerator.v:7154" *) _T_610;
  assign _T_784 = _T_750 & (* src = "crypto_accelerator.v:7155" *) _T_656;
  assign _T_786 = _T_742 & (* src = "crypto_accelerator.v:7156" *) _T_638;
  assign _T_931 = _T_913 & (* src = "crypto_accelerator.v:7224" *) _T_885;
  assign _T_933 = _T_915 & (* src = "crypto_accelerator.v:7225" *) _T_897;
  assign _T_937 = _T_895 & (* src = "crypto_accelerator.v:7227" *) shreg_io_output_0[0];
  assign _T_941 = _T_889 & (* src = "crypto_accelerator.v:7229" *) _T_917;
  assign _T_943 = _T_893 & (* src = "crypto_accelerator.v:7230" *) _T_883;
  assign _T_947 = _T_919 & (* src = "crypto_accelerator.v:7232" *) _T_909;
  assign _T_951 = _T_879 & (* src = "crypto_accelerator.v:7234" *) _T_891;
  assign _T_953 = _T_925 & (* src = "crypto_accelerator.v:7235" *) _T_921;
  assign _T_957 = _T_907 & (* src = "crypto_accelerator.v:7237" *) _T_903;
  assign _T_979 = _T_973 & (* src = "crypto_accelerator.v:7248" *) _T_969;
  assign _T_987 = _T_985 & (* src = "crypto_accelerator.v:7252" *) _T_983;
  assign _T_989 = _T_981 & (* src = "crypto_accelerator.v:7253" *) _T_977;
  assign _T_991 = _T_969 & (* src = "crypto_accelerator.v:7254" *) _T_975;
  assign _T_993 = _T_983 & (* src = "crypto_accelerator.v:7255" *) _T_991;
  assign _T_997 = _T_971 & (* src = "crypto_accelerator.v:7257" *) _T_973;
  assign _T_999 = _T_977 & (* src = "crypto_accelerator.v:7258" *) _T_997;
  assign _T_1021 = _T_1017 & (* src = "crypto_accelerator.v:7269" *) _T_885;
  assign _T_1023 = _T_1009 & (* src = "crypto_accelerator.v:7270" *) _T_897;
  assign _T_1025 = _T_1007 & (* src = "crypto_accelerator.v:7271" *) shreg_io_output_0[0];
  assign _T_1027 = _T_1015 & (* src = "crypto_accelerator.v:7272" *) _T_917;
  assign _T_1029 = _T_1005 & (* src = "crypto_accelerator.v:7273" *) _T_883;
  assign _T_1031 = _T_1003 & (* src = "crypto_accelerator.v:7274" *) _T_909;
  assign _T_1033 = _T_1013 & (* src = "crypto_accelerator.v:7275" *) _T_891;
  assign _T_1035 = _T_1019 & (* src = "crypto_accelerator.v:7276" *) _T_921;
  assign _T_1037 = _T_1011 & (* src = "crypto_accelerator.v:7277" *) _T_903;
  assign _T_1039 = _T_1017 & (* src = "crypto_accelerator.v:7278" *) _T_913;
  assign _T_1041 = _T_1009 & (* src = "crypto_accelerator.v:7279" *) _T_915;
  assign _T_1043 = _T_1007 & (* src = "crypto_accelerator.v:7280" *) _T_895;
  assign _T_1045 = _T_1015 & (* src = "crypto_accelerator.v:7281" *) _T_889;
  assign _T_1047 = _T_1005 & (* src = "crypto_accelerator.v:7282" *) _T_893;
  assign _T_1049 = _T_1003 & (* src = "crypto_accelerator.v:7283" *) _T_919;
  assign _T_1051 = _T_1013 & (* src = "crypto_accelerator.v:7284" *) _T_879;
  assign _T_1053 = _T_1019 & (* src = "crypto_accelerator.v:7285" *) _T_925;
  assign _T_1055 = _T_1011 & (* src = "crypto_accelerator.v:7286" *) _T_907;
  assign _T_1495 = enc_io_ready & (* src = "crypto_accelerator.v:7401" *) _T_1494;
  assign _T_1499 = dec_io_ready & (* src = "crypto_accelerator.v:7403" *) _T_1494;
  assign io_encReady = _T_1495 & (* src = "crypto_accelerator.v:7713" *) _T_1496;
  assign io_decReady = _T_1499 & (* src = "crypto_accelerator.v:7714" *) _T_1496;
  assign _T_6 = _T_2 == (* src = "crypto_accelerator.v:6804" *) { 3'b111, _GEN_42 };
  assign _GEN_6 = 1'b1 == (* src = "crypto_accelerator.v:7344" *) _T_1133;
  assign _002_ = 2'b10 == (* src = "crypto_accelerator.v:7345" *) _T_1133;
  assign _003_ = 2'b11 == (* src = "crypto_accelerator.v:7346" *) _T_1133;
  assign _004_ = 3'b100 == (* src = "crypto_accelerator.v:7347" *) _T_1133;
  assign _005_ = 3'b101 == (* src = "crypto_accelerator.v:7348" *) _T_1133;
  assign _006_ = 3'b110 == (* src = "crypto_accelerator.v:7349" *) _T_1133;
  assign _007_ = 3'b111 == (* src = "crypto_accelerator.v:7350" *) _T_1133;
  assign _008_ = 4'b1000 == (* src = "crypto_accelerator.v:7351" *) _T_1133;
  assign _009_ = 4'b1001 == (* src = "crypto_accelerator.v:7352" *) _T_1133;
  assign _010_ = 4'b1010 == (* src = "crypto_accelerator.v:7353" *) _T_1133;
  assign _011_ = 4'b1011 == (* src = "crypto_accelerator.v:7354" *) _T_1133;
  assign _012_ = 4'b1100 == (* src = "crypto_accelerator.v:7355" *) _T_1133;
  assign _013_ = 4'b1101 == (* src = "crypto_accelerator.v:7356" *) _T_1133;
  assign _014_ = 4'b1110 == (* src = "crypto_accelerator.v:7357" *) _T_1133;
  assign _015_ = 4'b1111 == (* src = "crypto_accelerator.v:7358" *) _T_1133;
  assign _GEN_22 = 1'b1 == (* src = "crypto_accelerator.v:7359" *) keyInd[3:0];
  assign _016_ = 2'b10 == (* src = "crypto_accelerator.v:7360" *) keyInd[3:0];
  assign _017_ = 2'b11 == (* src = "crypto_accelerator.v:7361" *) keyInd[3:0];
  assign _018_ = 3'b100 == (* src = "crypto_accelerator.v:7362" *) keyInd[3:0];
  assign _019_ = 3'b101 == (* src = "crypto_accelerator.v:7363" *) keyInd[3:0];
  assign _020_ = 3'b110 == (* src = "crypto_accelerator.v:7364" *) keyInd[3:0];
  assign _021_ = 3'b111 == (* src = "crypto_accelerator.v:7365" *) keyInd[3:0];
  assign _022_ = 4'b1000 == (* src = "crypto_accelerator.v:7366" *) keyInd[3:0];
  assign _023_ = 4'b1001 == (* src = "crypto_accelerator.v:7367" *) keyInd[3:0];
  assign _024_ = 4'b1010 == (* src = "crypto_accelerator.v:7368" *) keyInd[3:0];
  assign _025_ = 4'b1011 == (* src = "crypto_accelerator.v:7369" *) keyInd[3:0];
  assign _026_ = 4'b1100 == (* src = "crypto_accelerator.v:7370" *) keyInd[3:0];
  assign _027_ = 4'b1101 == (* src = "crypto_accelerator.v:7371" *) keyInd[3:0];
  assign _028_ = 4'b1110 == (* src = "crypto_accelerator.v:7372" *) keyInd[3:0];
  assign _029_ = 4'b1111 == (* src = "crypto_accelerator.v:7373" *) keyInd[3:0];
  assign _T_51 = ~ (* src = "crypto_accelerator.v:6805" *) keyInd[0];
  assign _T_289 = ~ (* src = "crypto_accelerator.v:6918" *) _T_288;
  assign _T_299 = ~ (* src = "crypto_accelerator.v:6925" *) _T_298;
  assign _T_307 = ~ (* src = "crypto_accelerator.v:6930" *) _T_306;
  assign _T_314 = ~ (* src = "crypto_accelerator.v:6935" *) _T_313;
  assign _T_558 = ~ (* src = "crypto_accelerator.v:7048" *) _T_557;
  assign _T_568 = ~ (* src = "crypto_accelerator.v:7055" *) _T_567;
  assign _T_576 = ~ (* src = "crypto_accelerator.v:7060" *) _T_575;
  assign _T_583 = ~ (* src = "crypto_accelerator.v:7065" *) _T_582;
  assign _T_827 = ~ (* src = "crypto_accelerator.v:7178" *) _T_826;
  assign _T_837 = ~ (* src = "crypto_accelerator.v:7185" *) _T_836;
  assign _T_845 = ~ (* src = "crypto_accelerator.v:7190" *) _T_844;
  assign _T_852 = ~ (* src = "crypto_accelerator.v:7195" *) _T_851;
  assign _T_1096 = ~ (* src = "crypto_accelerator.v:7308" *) _T_1095;
  assign _T_1106 = ~ (* src = "crypto_accelerator.v:7315" *) _T_1105;
  assign _T_1114 = ~ (* src = "crypto_accelerator.v:7320" *) _T_1113;
  assign _T_1121 = ~ (* src = "crypto_accelerator.v:7325" *) _T_1120;
  assign _T_1494 = ~ (* src = "crypto_accelerator.v:7400" *) keyUpdate;
  assign _T_1496 = ~ (* src = "crypto_accelerator.v:7402" *) io_keyValid;
  assign _GEN_0 = io_keyValid | (* src = "crypto_accelerator.v:6798" *) keyUpdate;
  assign _T = io_keyValid | (* src = "crypto_accelerator.v:6799" *) io_keyShift;
  assign _GEN_39 = keyUpdate | (* src = "crypto_accelerator.v:7399" *) _T;
  assign _T_1504 = enc_io_shift | (* src = "crypto_accelerator.v:7404" *) dec_io_shift;
  assign shreg_io_enable = _T_1504 | (* src = "crypto_accelerator.v:7723" *) _GEN_39;
  assign shreg_io_cyc = enc_io_shiftCyc | (* src = "crypto_accelerator.v:7725" *) dec_io_shiftCyc;
  always @(posedge clock)
      keyUpdate <= _001_;
  always @(posedge clock)
      keyInd <= _000_;
  assign _030_ = io_keyValid ? (* src = "crypto_accelerator.v:8057" *) 6'b000001 : keyInd;
  assign _031_ = keyUpdate ? (* src = "crypto_accelerator.v:8055" *) _T_2 : _030_;
  assign _000_ = reset ? (* src = "crypto_accelerator.v:8053" *) 6'b000000 : _031_;
  assign _032_ = _T_6 ? (* src = "crypto_accelerator.v:8045" *) 1'b0 : _GEN_0;
  assign _033_ = keyUpdate ? (* src = "crypto_accelerator.v:8044" *) _032_ : _GEN_0;
  assign _001_ = reset ? (* src = "crypto_accelerator.v:8042" *) 1'b0 : _033_;
  assign _GEN_3 = _T ? (* src = "crypto_accelerator.v:6800" *) io_keyIn : 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
  assign _GEN_42 = io_aes256 ? (* src = "crypto_accelerator.v:6802" *) 1'b0 : 1'b1;
  assign _T_1129_0_0 = io_aes256 ? (* src = "crypto_accelerator.v:7327" *) shreg_io_output_1[127:120] : shreg_io_output_0[127:120];
  assign _T_1129_0_1 = io_aes256 ? (* src = "crypto_accelerator.v:7328" *) shreg_io_output_1[119:112] : shreg_io_output_0[119:112];
  assign _T_1129_0_2 = io_aes256 ? (* src = "crypto_accelerator.v:7329" *) shreg_io_output_1[111:104] : shreg_io_output_0[111:104];
  assign _T_1129_0_3 = io_aes256 ? (* src = "crypto_accelerator.v:7330" *) shreg_io_output_1[103:96] : shreg_io_output_0[103:96];
  assign _T_1129_1_0 = io_aes256 ? (* src = "crypto_accelerator.v:7331" *) shreg_io_output_1[95:88] : shreg_io_output_0[95:88];
  assign _T_1129_1_1 = io_aes256 ? (* src = "crypto_accelerator.v:7332" *) shreg_io_output_1[87:80] : shreg_io_output_0[87:80];
  assign _T_1129_1_2 = io_aes256 ? (* src = "crypto_accelerator.v:7333" *) shreg_io_output_1[79:72] : shreg_io_output_0[79:72];
  assign _T_1129_1_3 = io_aes256 ? (* src = "crypto_accelerator.v:7334" *) shreg_io_output_1[71:64] : shreg_io_output_0[71:64];
  assign _T_1129_2_0 = io_aes256 ? (* src = "crypto_accelerator.v:7335" *) shreg_io_output_1[63:56] : shreg_io_output_0[63:56];
  assign _T_1129_2_1 = io_aes256 ? (* src = "crypto_accelerator.v:7336" *) shreg_io_output_1[55:48] : shreg_io_output_0[55:48];
  assign _T_1129_2_2 = io_aes256 ? (* src = "crypto_accelerator.v:7337" *) shreg_io_output_1[47:40] : shreg_io_output_0[47:40];
  assign _T_1129_2_3 = io_aes256 ? (* src = "crypto_accelerator.v:7338" *) shreg_io_output_1[39:32] : shreg_io_output_0[39:32];
  assign _T_1129_3_0 = io_aes256 ? (* src = "crypto_accelerator.v:7339" *) shreg_io_output_1[31:24] : shreg_io_output_0[31:24];
  assign _T_1129_3_1 = io_aes256 ? (* src = "crypto_accelerator.v:7340" *) shreg_io_output_1[23:16] : shreg_io_output_0[23:16];
  assign _T_1129_3_2 = io_aes256 ? (* src = "crypto_accelerator.v:7341" *) shreg_io_output_1[15:8] : shreg_io_output_0[15:8];
  assign _T_1129_3_3 = io_aes256 ? (* src = "crypto_accelerator.v:7342" *) shreg_io_output_1[7:0] : shreg_io_output_0[7:0];
  assign _GEN_7 = _002_ ? (* src = "crypto_accelerator.v:7345" *) 2'b10 : { 1'b0, _GEN_6 };
  assign _GEN_8 = _003_ ? (* src = "crypto_accelerator.v:7346" *) 3'b100 : { 1'b0, _GEN_7 };
  assign _GEN_9 = _004_ ? (* src = "crypto_accelerator.v:7347" *) 4'b1000 : { 1'b0, _GEN_8 };
  assign _GEN_10 = _005_ ? (* src = "crypto_accelerator.v:7348" *) 5'b10000 : { 1'b0, _GEN_9 };
  assign _GEN_11 = _006_ ? (* src = "crypto_accelerator.v:7349" *) 6'b100000 : { 1'b0, _GEN_10 };
  assign _GEN_12 = _007_ ? (* src = "crypto_accelerator.v:7350" *) 7'b1000000 : { 1'b0, _GEN_11 };
  assign _GEN_13 = _008_ ? (* src = "crypto_accelerator.v:7351" *) 8'b10000000 : { 1'b0, _GEN_12 };
  assign _GEN_14 = _009_ ? (* src = "crypto_accelerator.v:7352" *) 8'b00011011 : _GEN_13;
  assign _GEN_15 = _010_ ? (* src = "crypto_accelerator.v:7353" *) 8'b00110110 : _GEN_14;
  assign _GEN_16 = _011_ ? (* src = "crypto_accelerator.v:7354" *) 8'b01101100 : _GEN_15;
  assign _GEN_17 = _012_ ? (* src = "crypto_accelerator.v:7355" *) 8'b11011000 : _GEN_16;
  assign _GEN_18 = _013_ ? (* src = "crypto_accelerator.v:7356" *) 8'b10101011 : _GEN_17;
  assign _GEN_19 = _014_ ? (* src = "crypto_accelerator.v:7357" *) 8'b01001101 : _GEN_18;
  assign _GEN_20 = _015_ ? (* src = "crypto_accelerator.v:7358" *) 8'b10011010 : _GEN_19;
  assign _GEN_23 = _016_ ? (* src = "crypto_accelerator.v:7360" *) 2'b10 : { 1'b0, _GEN_22 };
  assign _GEN_24 = _017_ ? (* src = "crypto_accelerator.v:7361" *) 3'b100 : { 1'b0, _GEN_23 };
  assign _GEN_25 = _018_ ? (* src = "crypto_accelerator.v:7362" *) 4'b1000 : { 1'b0, _GEN_24 };
  assign _GEN_26 = _019_ ? (* src = "crypto_accelerator.v:7363" *) 5'b10000 : { 1'b0, _GEN_25 };
  assign _GEN_27 = _020_ ? (* src = "crypto_accelerator.v:7364" *) 6'b100000 : { 1'b0, _GEN_26 };
  assign _GEN_28 = _021_ ? (* src = "crypto_accelerator.v:7365" *) 7'b1000000 : { 1'b0, _GEN_27 };
  assign _GEN_29 = _022_ ? (* src = "crypto_accelerator.v:7366" *) 8'b10000000 : { 1'b0, _GEN_28 };
  assign _GEN_30 = _023_ ? (* src = "crypto_accelerator.v:7367" *) 8'b00011011 : _GEN_29;
  assign _GEN_31 = _024_ ? (* src = "crypto_accelerator.v:7368" *) 8'b00110110 : _GEN_30;
  assign _GEN_32 = _025_ ? (* src = "crypto_accelerator.v:7369" *) 8'b01101100 : _GEN_31;
  assign _GEN_33 = _026_ ? (* src = "crypto_accelerator.v:7370" *) 8'b11011000 : _GEN_32;
  assign _GEN_34 = _027_ ? (* src = "crypto_accelerator.v:7371" *) 8'b10101011 : _GEN_33;
  assign _GEN_35 = _028_ ? (* src = "crypto_accelerator.v:7372" *) 8'b01001101 : _GEN_34;
  assign _GEN_36 = _029_ ? (* src = "crypto_accelerator.v:7373" *) 8'b10011010 : _GEN_35;
  assign _T_1137 = io_aes256 ? (* src = "crypto_accelerator.v:7374" *) _GEN_20 : _GEN_36;
  assign _T_1138 = _T_52 ? (* src = "crypto_accelerator.v:7375" *) { _T_287, _T_314, _T_289, _T_292, _T_293, _T_310, _T_307, _T_299 } : { _T_556, _T_583, _T_558, _T_561, _T_562, _T_579, _T_576, _T_568 };
  assign _T_1140 = _T_52 ? (* src = "crypto_accelerator.v:7377" *) 8'b00000000 : _T_1137;
  assign _T_1142 = _T_52 ? (* src = "crypto_accelerator.v:7379" *) { _T_556, _T_583, _T_558, _T_561, _T_562, _T_579, _T_576, _T_568 } : { _T_825, _T_852, _T_827, _T_830, _T_831, _T_848, _T_845, _T_837 };
  assign _T_1144 = _T_52 ? (* src = "crypto_accelerator.v:7381" *) { _T_825, _T_852, _T_827, _T_830, _T_831, _T_848, _T_845, _T_837 } : { _T_1094, _T_1121, _T_1096, _T_1099, _T_1100, _T_1117, _T_1114, _T_1106 };
  assign _T_1146 = _T_52 ? (* src = "crypto_accelerator.v:7383" *) { _T_1094, _T_1121, _T_1096, _T_1099, _T_1100, _T_1117, _T_1114, _T_1106 } : { _T_287, _T_314, _T_289, _T_292, _T_293, _T_310, _T_307, _T_299 };
  assign shreg_io_input = keyUpdate ? (* src = "crypto_accelerator.v:7722" *) { _T_1141, _T_1143, _T_1145, _T_1147, _T_1149, _T_1150, _T_1151, _T_1152, _T_1154, _T_1155, _T_1156, _T_1157, _T_1159, _T_1160, _T_1161, _T_1162 } : _GEN_3;
  assign _T_70 = shreg_io_output_0[25] ^ (* src = "crypto_accelerator.v:6807" *) shreg_io_output_0[27];
  assign _T_72 = shreg_io_output_0[28] ^ (* src = "crypto_accelerator.v:6808" *) shreg_io_output_0[31];
  assign _T_74 = shreg_io_output_0[30] ^ (* src = "crypto_accelerator.v:6809" *) shreg_io_output_0[29];
  assign _T_76 = shreg_io_output_0[24] ^ (* src = "crypto_accelerator.v:6810" *) _T_74;
  assign _T_78 = _T_70 ^ (* src = "crypto_accelerator.v:6811" *) _T_72;
  assign _T_80 = shreg_io_output_0[30] ^ (* src = "crypto_accelerator.v:6812" *) shreg_io_output_0[26];
  assign _T_82 = shreg_io_output_0[31] ^ (* src = "crypto_accelerator.v:6813" *) shreg_io_output_0[25];
  assign _T_84 = _T_70 ^ (* src = "crypto_accelerator.v:6814" *) _T_80;
  assign _T_86 = shreg_io_output_0[25] ^ (* src = "crypto_accelerator.v:6815" *) _T_76;
  assign _T_88 = shreg_io_output_0[28] ^ (* src = "crypto_accelerator.v:6816" *) _T_76;
  assign _T_90 = shreg_io_output_0[24] ^ (* src = "crypto_accelerator.v:6817" *) _T_78;
  assign _T_92 = _T_78 ^ (* src = "crypto_accelerator.v:6818" *) _T_80;
  assign _T_94 = shreg_io_output_0[29] ^ (* src = "crypto_accelerator.v:6819" *) shreg_io_output_0[26];
  assign _T_96 = _T_74 ^ (* src = "crypto_accelerator.v:6820" *) _T_78;
  assign _T_98 = shreg_io_output_0[26] ^ (* src = "crypto_accelerator.v:6821" *) _T_82;
  assign _T_100 = shreg_io_output_0[31] ^ (* src = "crypto_accelerator.v:6822" *) shreg_io_output_0[26];
  assign _T_102 = shreg_io_output_0[24] ^ (* src = "crypto_accelerator.v:6823" *) _T_84;
  assign _T_104 = shreg_io_output_0[25] ^ (* src = "crypto_accelerator.v:6824" *) shreg_io_output_0[26];
  assign _T_106 = _T_72 ^ (* src = "crypto_accelerator.v:6825" *) _T_104;
  assign _T_108 = _T_76 ^ (* src = "crypto_accelerator.v:6826" *) _T_98;
  assign _T_110 = _T_70 ^ (* src = "crypto_accelerator.v:6827" *) _T_94;
  assign _T_112 = shreg_io_output_0[31] ^ (* src = "crypto_accelerator.v:6828" *) _T_76;
  assign _T_114 = _T_110 ^ (* src = "crypto_accelerator.v:6829" *) _T_78;
  assign _T_116 = _T_110 ^ (* src = "crypto_accelerator.v:6830" *) _T_82;
  assign _T_118 = _T_82 ^ (* src = "crypto_accelerator.v:6831" *) _T_106;
  assign _T_120 = _T_100 ^ (* src = "crypto_accelerator.v:6832" *) _T_96;
  assign _T_122 = _T_112 ^ (* src = "crypto_accelerator.v:6833" *) _T_102;
  assign _T_128 = _T_92 ^ (* src = "crypto_accelerator.v:6836" *) _T_124;
  assign _T_132 = _T_130 ^ (* src = "crypto_accelerator.v:6838" *) _T_124;
  assign _T_138 = _T_116 ^ (* src = "crypto_accelerator.v:6841" *) _T_134;
  assign _T_142 = _T_140 ^ (* src = "crypto_accelerator.v:6843" *) _T_134;
  assign _T_148 = _T_146 ^ (* src = "crypto_accelerator.v:6846" *) _T_144;
  assign _T_152 = _T_150 ^ (* src = "crypto_accelerator.v:6848" *) _T_144;
  assign _T_154 = _T_128 ^ (* src = "crypto_accelerator.v:6849" *) _T_126;
  assign _T_156 = _T_132 ^ (* src = "crypto_accelerator.v:6850" *) _T_120;
  assign _T_158 = _T_138 ^ (* src = "crypto_accelerator.v:6851" *) _T_136;
  assign _T_160 = _T_142 ^ (* src = "crypto_accelerator.v:6852" *) _T_152;
  assign _T_162 = _T_154 ^ (* src = "crypto_accelerator.v:6853" *) _T_148;
  assign _T_164 = _T_156 ^ (* src = "crypto_accelerator.v:6854" *) _T_152;
  assign _T_166 = _T_158 ^ (* src = "crypto_accelerator.v:6855" *) _T_148;
  assign _T_168 = _T_160 ^ (* src = "crypto_accelerator.v:6856" *) _T_122;
  assign _T_170 = _T_166 ^ (* src = "crypto_accelerator.v:6857" *) _T_168;
  assign _T_174 = _T_164 ^ (* src = "crypto_accelerator.v:6859" *) _T_172;
  assign _T_176 = _T_162 ^ (* src = "crypto_accelerator.v:6860" *) _T_164;
  assign _T_178 = _T_168 ^ (* src = "crypto_accelerator.v:6861" *) _T_172;
  assign _T_188 = _T_176 ^ (* src = "crypto_accelerator.v:6866" *) _T_172;
  assign _T_194 = _T_170 ^ (* src = "crypto_accelerator.v:6869" *) _T_172;
  assign _T_196 = _T_164 ^ (* src = "crypto_accelerator.v:6870" *) _T_180;
  assign _T_198 = _T_186 ^ (* src = "crypto_accelerator.v:6871" *) _T_188;
  assign _T_200 = _T_168 ^ (* src = "crypto_accelerator.v:6872" *) _T_182;
  assign _T_202 = _T_192 ^ (* src = "crypto_accelerator.v:6873" *) _T_194;
  assign _T_204 = _T_198 ^ (* src = "crypto_accelerator.v:6874" *) _T_202;
  assign _T_206 = _T_196 ^ (* src = "crypto_accelerator.v:6875" *) _T_200;
  assign _T_208 = _T_196 ^ (* src = "crypto_accelerator.v:6876" *) _T_198;
  assign _T_210 = _T_200 ^ (* src = "crypto_accelerator.v:6877" *) _T_202;
  assign _T_212 = _T_206 ^ (* src = "crypto_accelerator.v:6878" *) _T_204;
  assign _T_250 = _T_244 ^ (* src = "crypto_accelerator.v:6897" *) _T_246;
  assign _T_252 = _T_222 ^ (* src = "crypto_accelerator.v:6898" *) _T_234;
  assign _T_254 = _T_228 ^ (* src = "crypto_accelerator.v:6899" *) _T_250;
  assign _T_256 = _T_232 ^ (* src = "crypto_accelerator.v:6900" *) _T_252;
  assign _T_258 = _T_218 ^ (* src = "crypto_accelerator.v:6901" *) _T_238;
  assign _T_260 = _T_214 ^ (* src = "crypto_accelerator.v:6902" *) _T_220;
  assign _T_262 = _T_250 ^ (* src = "crypto_accelerator.v:6903" *) _T_260;
  assign _T_264 = _T_216 ^ (* src = "crypto_accelerator.v:6904" *) _T_256;
  assign _T_266 = _T_214 ^ (* src = "crypto_accelerator.v:6905" *) _T_226;
  assign _T_268 = _T_224 ^ (* src = "crypto_accelerator.v:6906" *) _T_240;
  assign _T_270 = _T_230 ^ (* src = "crypto_accelerator.v:6907" *) _T_242;
  assign _T_272 = _T_218 ^ (* src = "crypto_accelerator.v:6908" *) _T_264;
  assign _T_274 = _T_258 ^ (* src = "crypto_accelerator.v:6909" *) _T_270;
  assign _T_276 = _T_236 ^ (* src = "crypto_accelerator.v:6910" *) _T_252;
  assign _T_278 = _T_220 ^ (* src = "crypto_accelerator.v:6911" *) _T_226;
  assign _T_280 = _T_256 ^ (* src = "crypto_accelerator.v:6912" *) _T_278;
  assign _T_282 = _T_248 ^ (* src = "crypto_accelerator.v:6913" *) _T_274;
  assign _T_284 = _T_244 ^ (* src = "crypto_accelerator.v:6914" *) _T_266;
  assign _T_286 = _T_258 ^ (* src = "crypto_accelerator.v:6915" *) _T_268;
  assign _T_287 = _T_254 ^ (* src = "crypto_accelerator.v:6916" *) _T_280;
  assign _T_288 = _T_282 ^ (* src = "crypto_accelerator.v:6917" *) _T_284;
  assign _T_291 = _T_224 ^ (* src = "crypto_accelerator.v:6919" *) _T_250;
  assign _T_292 = _T_262 ^ (* src = "crypto_accelerator.v:6920" *) _T_264;
  assign _T_293 = _T_272 ^ (* src = "crypto_accelerator.v:6921" *) _T_291;
  assign _T_295 = _T_222 ^ (* src = "crypto_accelerator.v:6922" *) _T_238;
  assign _T_297 = _T_260 ^ (* src = "crypto_accelerator.v:6923" *) _T_276;
  assign _T_298 = _T_262 ^ (* src = "crypto_accelerator.v:6924" *) _T_286;
  assign _T_301 = _T_230 ^ (* src = "crypto_accelerator.v:6926" *) _T_268;
  assign _T_303 = _T_295 ^ (* src = "crypto_accelerator.v:6927" *) _T_301;
  assign _T_305 = _T_222 ^ (* src = "crypto_accelerator.v:6928" *) _T_266;
  assign _T_306 = _T_254 ^ (* src = "crypto_accelerator.v:6929" *) _T_303;
  assign _T_309 = _T_274 ^ (* src = "crypto_accelerator.v:6931" *) _T_297;
  assign _T_310 = _T_254 ^ (* src = "crypto_accelerator.v:6932" *) _T_309;
  assign _T_312 = _T_264 ^ (* src = "crypto_accelerator.v:6933" *) _T_305;
  assign _T_313 = _T_254 ^ (* src = "crypto_accelerator.v:6934" *) _T_312;
  assign _T_339 = shreg_io_output_0[17] ^ (* src = "crypto_accelerator.v:6937" *) shreg_io_output_0[19];
  assign _T_341 = shreg_io_output_0[20] ^ (* src = "crypto_accelerator.v:6938" *) shreg_io_output_0[23];
  assign _T_343 = shreg_io_output_0[22] ^ (* src = "crypto_accelerator.v:6939" *) shreg_io_output_0[21];
  assign _T_345 = shreg_io_output_0[16] ^ (* src = "crypto_accelerator.v:6940" *) _T_343;
  assign _T_347 = _T_339 ^ (* src = "crypto_accelerator.v:6941" *) _T_341;
  assign _T_349 = shreg_io_output_0[22] ^ (* src = "crypto_accelerator.v:6942" *) shreg_io_output_0[18];
  assign _T_351 = shreg_io_output_0[23] ^ (* src = "crypto_accelerator.v:6943" *) shreg_io_output_0[17];
  assign _T_353 = _T_339 ^ (* src = "crypto_accelerator.v:6944" *) _T_349;
  assign _T_355 = shreg_io_output_0[17] ^ (* src = "crypto_accelerator.v:6945" *) _T_345;
  assign _T_357 = shreg_io_output_0[20] ^ (* src = "crypto_accelerator.v:6946" *) _T_345;
  assign _T_359 = shreg_io_output_0[16] ^ (* src = "crypto_accelerator.v:6947" *) _T_347;
  assign _T_361 = _T_347 ^ (* src = "crypto_accelerator.v:6948" *) _T_349;
  assign _T_363 = shreg_io_output_0[21] ^ (* src = "crypto_accelerator.v:6949" *) shreg_io_output_0[18];
  assign _T_365 = _T_343 ^ (* src = "crypto_accelerator.v:6950" *) _T_347;
  assign _T_367 = shreg_io_output_0[18] ^ (* src = "crypto_accelerator.v:6951" *) _T_351;
  assign _T_369 = shreg_io_output_0[23] ^ (* src = "crypto_accelerator.v:6952" *) shreg_io_output_0[18];
  assign _T_371 = shreg_io_output_0[16] ^ (* src = "crypto_accelerator.v:6953" *) _T_353;
  assign _T_373 = shreg_io_output_0[17] ^ (* src = "crypto_accelerator.v:6954" *) shreg_io_output_0[18];
  assign _T_375 = _T_341 ^ (* src = "crypto_accelerator.v:6955" *) _T_373;
  assign _T_377 = _T_345 ^ (* src = "crypto_accelerator.v:6956" *) _T_367;
  assign _T_379 = _T_339 ^ (* src = "crypto_accelerator.v:6957" *) _T_363;
  assign _T_381 = shreg_io_output_0[23] ^ (* src = "crypto_accelerator.v:6958" *) _T_345;
  assign _T_383 = _T_379 ^ (* src = "crypto_accelerator.v:6959" *) _T_347;
  assign _T_385 = _T_379 ^ (* src = "crypto_accelerator.v:6960" *) _T_351;
  assign _T_387 = _T_351 ^ (* src = "crypto_accelerator.v:6961" *) _T_375;
  assign _T_389 = _T_369 ^ (* src = "crypto_accelerator.v:6962" *) _T_365;
  assign _T_391 = _T_381 ^ (* src = "crypto_accelerator.v:6963" *) _T_371;
  assign _T_397 = _T_361 ^ (* src = "crypto_accelerator.v:6966" *) _T_393;
  assign _T_401 = _T_399 ^ (* src = "crypto_accelerator.v:6968" *) _T_393;
  assign _T_407 = _T_385 ^ (* src = "crypto_accelerator.v:6971" *) _T_403;
  assign _T_411 = _T_409 ^ (* src = "crypto_accelerator.v:6973" *) _T_403;
  assign _T_417 = _T_415 ^ (* src = "crypto_accelerator.v:6976" *) _T_413;
  assign _T_421 = _T_419 ^ (* src = "crypto_accelerator.v:6978" *) _T_413;
  assign _T_423 = _T_397 ^ (* src = "crypto_accelerator.v:6979" *) _T_395;
  assign _T_425 = _T_401 ^ (* src = "crypto_accelerator.v:6980" *) _T_389;
  assign _T_427 = _T_407 ^ (* src = "crypto_accelerator.v:6981" *) _T_405;
  assign _T_429 = _T_411 ^ (* src = "crypto_accelerator.v:6982" *) _T_421;
  assign _T_431 = _T_423 ^ (* src = "crypto_accelerator.v:6983" *) _T_417;
  assign _T_433 = _T_425 ^ (* src = "crypto_accelerator.v:6984" *) _T_421;
  assign _T_435 = _T_427 ^ (* src = "crypto_accelerator.v:6985" *) _T_417;
  assign _T_437 = _T_429 ^ (* src = "crypto_accelerator.v:6986" *) _T_391;
  assign _T_439 = _T_435 ^ (* src = "crypto_accelerator.v:6987" *) _T_437;
  assign _T_443 = _T_433 ^ (* src = "crypto_accelerator.v:6989" *) _T_441;
  assign _T_445 = _T_431 ^ (* src = "crypto_accelerator.v:6990" *) _T_433;
  assign _T_447 = _T_437 ^ (* src = "crypto_accelerator.v:6991" *) _T_441;
  assign _T_457 = _T_445 ^ (* src = "crypto_accelerator.v:6996" *) _T_441;
  assign _T_463 = _T_439 ^ (* src = "crypto_accelerator.v:6999" *) _T_441;
  assign _T_465 = _T_433 ^ (* src = "crypto_accelerator.v:7000" *) _T_449;
  assign _T_467 = _T_455 ^ (* src = "crypto_accelerator.v:7001" *) _T_457;
  assign _T_469 = _T_437 ^ (* src = "crypto_accelerator.v:7002" *) _T_451;
  assign _T_471 = _T_461 ^ (* src = "crypto_accelerator.v:7003" *) _T_463;
  assign _T_473 = _T_467 ^ (* src = "crypto_accelerator.v:7004" *) _T_471;
  assign _T_475 = _T_465 ^ (* src = "crypto_accelerator.v:7005" *) _T_469;
  assign _T_477 = _T_465 ^ (* src = "crypto_accelerator.v:7006" *) _T_467;
  assign _T_479 = _T_469 ^ (* src = "crypto_accelerator.v:7007" *) _T_471;
  assign _T_481 = _T_475 ^ (* src = "crypto_accelerator.v:7008" *) _T_473;
  assign _T_519 = _T_513 ^ (* src = "crypto_accelerator.v:7027" *) _T_515;
  assign _T_521 = _T_491 ^ (* src = "crypto_accelerator.v:7028" *) _T_503;
  assign _T_523 = _T_497 ^ (* src = "crypto_accelerator.v:7029" *) _T_519;
  assign _T_525 = _T_501 ^ (* src = "crypto_accelerator.v:7030" *) _T_521;
  assign _T_527 = _T_487 ^ (* src = "crypto_accelerator.v:7031" *) _T_507;
  assign _T_529 = _T_483 ^ (* src = "crypto_accelerator.v:7032" *) _T_489;
  assign _T_531 = _T_519 ^ (* src = "crypto_accelerator.v:7033" *) _T_529;
  assign _T_533 = _T_485 ^ (* src = "crypto_accelerator.v:7034" *) _T_525;
  assign _T_535 = _T_483 ^ (* src = "crypto_accelerator.v:7035" *) _T_495;
  assign _T_537 = _T_493 ^ (* src = "crypto_accelerator.v:7036" *) _T_509;
  assign _T_539 = _T_499 ^ (* src = "crypto_accelerator.v:7037" *) _T_511;
  assign _T_541 = _T_487 ^ (* src = "crypto_accelerator.v:7038" *) _T_533;
  assign _T_543 = _T_527 ^ (* src = "crypto_accelerator.v:7039" *) _T_539;
  assign _T_545 = _T_505 ^ (* src = "crypto_accelerator.v:7040" *) _T_521;
  assign _T_547 = _T_489 ^ (* src = "crypto_accelerator.v:7041" *) _T_495;
  assign _T_549 = _T_525 ^ (* src = "crypto_accelerator.v:7042" *) _T_547;
  assign _T_551 = _T_517 ^ (* src = "crypto_accelerator.v:7043" *) _T_543;
  assign _T_553 = _T_513 ^ (* src = "crypto_accelerator.v:7044" *) _T_535;
  assign _T_555 = _T_527 ^ (* src = "crypto_accelerator.v:7045" *) _T_537;
  assign _T_556 = _T_523 ^ (* src = "crypto_accelerator.v:7046" *) _T_549;
  assign _T_557 = _T_551 ^ (* src = "crypto_accelerator.v:7047" *) _T_553;
  assign _T_560 = _T_493 ^ (* src = "crypto_accelerator.v:7049" *) _T_519;
  assign _T_561 = _T_531 ^ (* src = "crypto_accelerator.v:7050" *) _T_533;
  assign _T_562 = _T_541 ^ (* src = "crypto_accelerator.v:7051" *) _T_560;
  assign _T_564 = _T_491 ^ (* src = "crypto_accelerator.v:7052" *) _T_507;
  assign _T_566 = _T_529 ^ (* src = "crypto_accelerator.v:7053" *) _T_545;
  assign _T_567 = _T_531 ^ (* src = "crypto_accelerator.v:7054" *) _T_555;
  assign _T_570 = _T_499 ^ (* src = "crypto_accelerator.v:7056" *) _T_537;
  assign _T_572 = _T_564 ^ (* src = "crypto_accelerator.v:7057" *) _T_570;
  assign _T_574 = _T_491 ^ (* src = "crypto_accelerator.v:7058" *) _T_535;
  assign _T_575 = _T_523 ^ (* src = "crypto_accelerator.v:7059" *) _T_572;
  assign _T_578 = _T_543 ^ (* src = "crypto_accelerator.v:7061" *) _T_566;
  assign _T_579 = _T_523 ^ (* src = "crypto_accelerator.v:7062" *) _T_578;
  assign _T_581 = _T_533 ^ (* src = "crypto_accelerator.v:7063" *) _T_574;
  assign _T_582 = _T_523 ^ (* src = "crypto_accelerator.v:7064" *) _T_581;
  assign _T_608 = shreg_io_output_0[9] ^ (* src = "crypto_accelerator.v:7067" *) shreg_io_output_0[11];
  assign _T_610 = shreg_io_output_0[12] ^ (* src = "crypto_accelerator.v:7068" *) shreg_io_output_0[15];
  assign _T_612 = shreg_io_output_0[14] ^ (* src = "crypto_accelerator.v:7069" *) shreg_io_output_0[13];
  assign _T_614 = shreg_io_output_0[8] ^ (* src = "crypto_accelerator.v:7070" *) _T_612;
  assign _T_616 = _T_608 ^ (* src = "crypto_accelerator.v:7071" *) _T_610;
  assign _T_618 = shreg_io_output_0[14] ^ (* src = "crypto_accelerator.v:7072" *) shreg_io_output_0[10];
  assign _T_620 = shreg_io_output_0[15] ^ (* src = "crypto_accelerator.v:7073" *) shreg_io_output_0[9];
  assign _T_622 = _T_608 ^ (* src = "crypto_accelerator.v:7074" *) _T_618;
  assign _T_624 = shreg_io_output_0[9] ^ (* src = "crypto_accelerator.v:7075" *) _T_614;
  assign _T_626 = shreg_io_output_0[12] ^ (* src = "crypto_accelerator.v:7076" *) _T_614;
  assign _T_628 = shreg_io_output_0[8] ^ (* src = "crypto_accelerator.v:7077" *) _T_616;
  assign _T_630 = _T_616 ^ (* src = "crypto_accelerator.v:7078" *) _T_618;
  assign _T_632 = shreg_io_output_0[13] ^ (* src = "crypto_accelerator.v:7079" *) shreg_io_output_0[10];
  assign _T_634 = _T_612 ^ (* src = "crypto_accelerator.v:7080" *) _T_616;
  assign _T_636 = shreg_io_output_0[10] ^ (* src = "crypto_accelerator.v:7081" *) _T_620;
  assign _T_638 = shreg_io_output_0[15] ^ (* src = "crypto_accelerator.v:7082" *) shreg_io_output_0[10];
  assign _T_640 = shreg_io_output_0[8] ^ (* src = "crypto_accelerator.v:7083" *) _T_622;
  assign _T_642 = shreg_io_output_0[9] ^ (* src = "crypto_accelerator.v:7084" *) shreg_io_output_0[10];
  assign _T_644 = _T_610 ^ (* src = "crypto_accelerator.v:7085" *) _T_642;
  assign _T_646 = _T_614 ^ (* src = "crypto_accelerator.v:7086" *) _T_636;
  assign _T_648 = _T_608 ^ (* src = "crypto_accelerator.v:7087" *) _T_632;
  assign _T_650 = shreg_io_output_0[15] ^ (* src = "crypto_accelerator.v:7088" *) _T_614;
  assign _T_652 = _T_648 ^ (* src = "crypto_accelerator.v:7089" *) _T_616;
  assign _T_654 = _T_648 ^ (* src = "crypto_accelerator.v:7090" *) _T_620;
  assign _T_656 = _T_620 ^ (* src = "crypto_accelerator.v:7091" *) _T_644;
  assign _T_658 = _T_638 ^ (* src = "crypto_accelerator.v:7092" *) _T_634;
  assign _T_660 = _T_650 ^ (* src = "crypto_accelerator.v:7093" *) _T_640;
  assign _T_666 = _T_630 ^ (* src = "crypto_accelerator.v:7096" *) _T_662;
  assign _T_670 = _T_668 ^ (* src = "crypto_accelerator.v:7098" *) _T_662;
  assign _T_676 = _T_654 ^ (* src = "crypto_accelerator.v:7101" *) _T_672;
  assign _T_680 = _T_678 ^ (* src = "crypto_accelerator.v:7103" *) _T_672;
  assign _T_686 = _T_684 ^ (* src = "crypto_accelerator.v:7106" *) _T_682;
  assign _T_690 = _T_688 ^ (* src = "crypto_accelerator.v:7108" *) _T_682;
  assign _T_692 = _T_666 ^ (* src = "crypto_accelerator.v:7109" *) _T_664;
  assign _T_694 = _T_670 ^ (* src = "crypto_accelerator.v:7110" *) _T_658;
  assign _T_696 = _T_676 ^ (* src = "crypto_accelerator.v:7111" *) _T_674;
  assign _T_698 = _T_680 ^ (* src = "crypto_accelerator.v:7112" *) _T_690;
  assign _T_700 = _T_692 ^ (* src = "crypto_accelerator.v:7113" *) _T_686;
  assign _T_702 = _T_694 ^ (* src = "crypto_accelerator.v:7114" *) _T_690;
  assign _T_704 = _T_696 ^ (* src = "crypto_accelerator.v:7115" *) _T_686;
  assign _T_706 = _T_698 ^ (* src = "crypto_accelerator.v:7116" *) _T_660;
  assign _T_708 = _T_704 ^ (* src = "crypto_accelerator.v:7117" *) _T_706;
  assign _T_712 = _T_702 ^ (* src = "crypto_accelerator.v:7119" *) _T_710;
  assign _T_714 = _T_700 ^ (* src = "crypto_accelerator.v:7120" *) _T_702;
  assign _T_716 = _T_706 ^ (* src = "crypto_accelerator.v:7121" *) _T_710;
  assign _T_726 = _T_714 ^ (* src = "crypto_accelerator.v:7126" *) _T_710;
  assign _T_732 = _T_708 ^ (* src = "crypto_accelerator.v:7129" *) _T_710;
  assign _T_734 = _T_702 ^ (* src = "crypto_accelerator.v:7130" *) _T_718;
  assign _T_736 = _T_724 ^ (* src = "crypto_accelerator.v:7131" *) _T_726;
  assign _T_738 = _T_706 ^ (* src = "crypto_accelerator.v:7132" *) _T_720;
  assign _T_740 = _T_730 ^ (* src = "crypto_accelerator.v:7133" *) _T_732;
  assign _T_742 = _T_736 ^ (* src = "crypto_accelerator.v:7134" *) _T_740;
  assign _T_744 = _T_734 ^ (* src = "crypto_accelerator.v:7135" *) _T_738;
  assign _T_746 = _T_734 ^ (* src = "crypto_accelerator.v:7136" *) _T_736;
  assign _T_748 = _T_738 ^ (* src = "crypto_accelerator.v:7137" *) _T_740;
  assign _T_750 = _T_744 ^ (* src = "crypto_accelerator.v:7138" *) _T_742;
  assign _T_788 = _T_782 ^ (* src = "crypto_accelerator.v:7157" *) _T_784;
  assign _T_790 = _T_760 ^ (* src = "crypto_accelerator.v:7158" *) _T_772;
  assign _T_792 = _T_766 ^ (* src = "crypto_accelerator.v:7159" *) _T_788;
  assign _T_794 = _T_770 ^ (* src = "crypto_accelerator.v:7160" *) _T_790;
  assign _T_796 = _T_756 ^ (* src = "crypto_accelerator.v:7161" *) _T_776;
  assign _T_798 = _T_752 ^ (* src = "crypto_accelerator.v:7162" *) _T_758;
  assign _T_800 = _T_788 ^ (* src = "crypto_accelerator.v:7163" *) _T_798;
  assign _T_802 = _T_754 ^ (* src = "crypto_accelerator.v:7164" *) _T_794;
  assign _T_804 = _T_752 ^ (* src = "crypto_accelerator.v:7165" *) _T_764;
  assign _T_806 = _T_762 ^ (* src = "crypto_accelerator.v:7166" *) _T_778;
  assign _T_808 = _T_768 ^ (* src = "crypto_accelerator.v:7167" *) _T_780;
  assign _T_810 = _T_756 ^ (* src = "crypto_accelerator.v:7168" *) _T_802;
  assign _T_812 = _T_796 ^ (* src = "crypto_accelerator.v:7169" *) _T_808;
  assign _T_814 = _T_774 ^ (* src = "crypto_accelerator.v:7170" *) _T_790;
  assign _T_816 = _T_758 ^ (* src = "crypto_accelerator.v:7171" *) _T_764;
  assign _T_818 = _T_794 ^ (* src = "crypto_accelerator.v:7172" *) _T_816;
  assign _T_820 = _T_786 ^ (* src = "crypto_accelerator.v:7173" *) _T_812;
  assign _T_822 = _T_782 ^ (* src = "crypto_accelerator.v:7174" *) _T_804;
  assign _T_824 = _T_796 ^ (* src = "crypto_accelerator.v:7175" *) _T_806;
  assign _T_825 = _T_792 ^ (* src = "crypto_accelerator.v:7176" *) _T_818;
  assign _T_826 = _T_820 ^ (* src = "crypto_accelerator.v:7177" *) _T_822;
  assign _T_829 = _T_762 ^ (* src = "crypto_accelerator.v:7179" *) _T_788;
  assign _T_830 = _T_800 ^ (* src = "crypto_accelerator.v:7180" *) _T_802;
  assign _T_831 = _T_810 ^ (* src = "crypto_accelerator.v:7181" *) _T_829;
  assign _T_833 = _T_760 ^ (* src = "crypto_accelerator.v:7182" *) _T_776;
  assign _T_835 = _T_798 ^ (* src = "crypto_accelerator.v:7183" *) _T_814;
  assign _T_836 = _T_800 ^ (* src = "crypto_accelerator.v:7184" *) _T_824;
  assign _T_839 = _T_768 ^ (* src = "crypto_accelerator.v:7186" *) _T_806;
  assign _T_841 = _T_833 ^ (* src = "crypto_accelerator.v:7187" *) _T_839;
  assign _T_843 = _T_760 ^ (* src = "crypto_accelerator.v:7188" *) _T_804;
  assign _T_844 = _T_792 ^ (* src = "crypto_accelerator.v:7189" *) _T_841;
  assign _T_847 = _T_812 ^ (* src = "crypto_accelerator.v:7191" *) _T_835;
  assign _T_848 = _T_792 ^ (* src = "crypto_accelerator.v:7192" *) _T_847;
  assign _T_850 = _T_802 ^ (* src = "crypto_accelerator.v:7193" *) _T_843;
  assign _T_851 = _T_792 ^ (* src = "crypto_accelerator.v:7194" *) _T_850;
  assign _T_877 = shreg_io_output_0[1] ^ (* src = "crypto_accelerator.v:7197" *) shreg_io_output_0[3];
  assign _T_879 = shreg_io_output_0[4] ^ (* src = "crypto_accelerator.v:7198" *) shreg_io_output_0[7];
  assign _T_881 = shreg_io_output_0[6] ^ (* src = "crypto_accelerator.v:7199" *) shreg_io_output_0[5];
  assign _T_883 = shreg_io_output_0[0] ^ (* src = "crypto_accelerator.v:7200" *) _T_881;
  assign _T_885 = _T_877 ^ (* src = "crypto_accelerator.v:7201" *) _T_879;
  assign _T_887 = shreg_io_output_0[6] ^ (* src = "crypto_accelerator.v:7202" *) shreg_io_output_0[2];
  assign _T_889 = shreg_io_output_0[7] ^ (* src = "crypto_accelerator.v:7203" *) shreg_io_output_0[1];
  assign _T_891 = _T_877 ^ (* src = "crypto_accelerator.v:7204" *) _T_887;
  assign _T_893 = shreg_io_output_0[1] ^ (* src = "crypto_accelerator.v:7205" *) _T_883;
  assign _T_895 = shreg_io_output_0[4] ^ (* src = "crypto_accelerator.v:7206" *) _T_883;
  assign _T_897 = shreg_io_output_0[0] ^ (* src = "crypto_accelerator.v:7207" *) _T_885;
  assign _T_899 = _T_885 ^ (* src = "crypto_accelerator.v:7208" *) _T_887;
  assign _T_901 = shreg_io_output_0[5] ^ (* src = "crypto_accelerator.v:7209" *) shreg_io_output_0[2];
  assign _T_903 = _T_881 ^ (* src = "crypto_accelerator.v:7210" *) _T_885;
  assign _T_905 = shreg_io_output_0[2] ^ (* src = "crypto_accelerator.v:7211" *) _T_889;
  assign _T_907 = shreg_io_output_0[7] ^ (* src = "crypto_accelerator.v:7212" *) shreg_io_output_0[2];
  assign _T_909 = shreg_io_output_0[0] ^ (* src = "crypto_accelerator.v:7213" *) _T_891;
  assign _T_911 = shreg_io_output_0[1] ^ (* src = "crypto_accelerator.v:7214" *) shreg_io_output_0[2];
  assign _T_913 = _T_879 ^ (* src = "crypto_accelerator.v:7215" *) _T_911;
  assign _T_915 = _T_883 ^ (* src = "crypto_accelerator.v:7216" *) _T_905;
  assign _T_917 = _T_877 ^ (* src = "crypto_accelerator.v:7217" *) _T_901;
  assign _T_919 = shreg_io_output_0[7] ^ (* src = "crypto_accelerator.v:7218" *) _T_883;
  assign _T_921 = _T_917 ^ (* src = "crypto_accelerator.v:7219" *) _T_885;
  assign _T_923 = _T_917 ^ (* src = "crypto_accelerator.v:7220" *) _T_889;
  assign _T_925 = _T_889 ^ (* src = "crypto_accelerator.v:7221" *) _T_913;
  assign _T_927 = _T_907 ^ (* src = "crypto_accelerator.v:7222" *) _T_903;
  assign _T_929 = _T_919 ^ (* src = "crypto_accelerator.v:7223" *) _T_909;
  assign _T_935 = _T_899 ^ (* src = "crypto_accelerator.v:7226" *) _T_931;
  assign _T_939 = _T_937 ^ (* src = "crypto_accelerator.v:7228" *) _T_931;
  assign _T_945 = _T_923 ^ (* src = "crypto_accelerator.v:7231" *) _T_941;
  assign _T_949 = _T_947 ^ (* src = "crypto_accelerator.v:7233" *) _T_941;
  assign _T_955 = _T_953 ^ (* src = "crypto_accelerator.v:7236" *) _T_951;
  assign _T_959 = _T_957 ^ (* src = "crypto_accelerator.v:7238" *) _T_951;
  assign _T_961 = _T_935 ^ (* src = "crypto_accelerator.v:7239" *) _T_933;
  assign _T_963 = _T_939 ^ (* src = "crypto_accelerator.v:7240" *) _T_927;
  assign _T_965 = _T_945 ^ (* src = "crypto_accelerator.v:7241" *) _T_943;
  assign _T_967 = _T_949 ^ (* src = "crypto_accelerator.v:7242" *) _T_959;
  assign _T_969 = _T_961 ^ (* src = "crypto_accelerator.v:7243" *) _T_955;
  assign _T_971 = _T_963 ^ (* src = "crypto_accelerator.v:7244" *) _T_959;
  assign _T_973 = _T_965 ^ (* src = "crypto_accelerator.v:7245" *) _T_955;
  assign _T_975 = _T_967 ^ (* src = "crypto_accelerator.v:7246" *) _T_929;
  assign _T_977 = _T_973 ^ (* src = "crypto_accelerator.v:7247" *) _T_975;
  assign _T_981 = _T_971 ^ (* src = "crypto_accelerator.v:7249" *) _T_979;
  assign _T_983 = _T_969 ^ (* src = "crypto_accelerator.v:7250" *) _T_971;
  assign _T_985 = _T_975 ^ (* src = "crypto_accelerator.v:7251" *) _T_979;
  assign _T_995 = _T_983 ^ (* src = "crypto_accelerator.v:7256" *) _T_979;
  assign _T_1001 = _T_977 ^ (* src = "crypto_accelerator.v:7259" *) _T_979;
  assign _T_1003 = _T_971 ^ (* src = "crypto_accelerator.v:7260" *) _T_987;
  assign _T_1005 = _T_993 ^ (* src = "crypto_accelerator.v:7261" *) _T_995;
  assign _T_1007 = _T_975 ^ (* src = "crypto_accelerator.v:7262" *) _T_989;
  assign _T_1009 = _T_999 ^ (* src = "crypto_accelerator.v:7263" *) _T_1001;
  assign _T_1011 = _T_1005 ^ (* src = "crypto_accelerator.v:7264" *) _T_1009;
  assign _T_1013 = _T_1003 ^ (* src = "crypto_accelerator.v:7265" *) _T_1007;
  assign _T_1015 = _T_1003 ^ (* src = "crypto_accelerator.v:7266" *) _T_1005;
  assign _T_1017 = _T_1007 ^ (* src = "crypto_accelerator.v:7267" *) _T_1009;
  assign _T_1019 = _T_1013 ^ (* src = "crypto_accelerator.v:7268" *) _T_1011;
  assign _T_1057 = _T_1051 ^ (* src = "crypto_accelerator.v:7287" *) _T_1053;
  assign _T_1059 = _T_1029 ^ (* src = "crypto_accelerator.v:7288" *) _T_1041;
  assign _T_1061 = _T_1035 ^ (* src = "crypto_accelerator.v:7289" *) _T_1057;
  assign _T_1063 = _T_1039 ^ (* src = "crypto_accelerator.v:7290" *) _T_1059;
  assign _T_1065 = _T_1025 ^ (* src = "crypto_accelerator.v:7291" *) _T_1045;
  assign _T_1067 = _T_1021 ^ (* src = "crypto_accelerator.v:7292" *) _T_1027;
  assign _T_1069 = _T_1057 ^ (* src = "crypto_accelerator.v:7293" *) _T_1067;
  assign _T_1071 = _T_1023 ^ (* src = "crypto_accelerator.v:7294" *) _T_1063;
  assign _T_1073 = _T_1021 ^ (* src = "crypto_accelerator.v:7295" *) _T_1033;
  assign _T_1075 = _T_1031 ^ (* src = "crypto_accelerator.v:7296" *) _T_1047;
  assign _T_1077 = _T_1037 ^ (* src = "crypto_accelerator.v:7297" *) _T_1049;
  assign _T_1079 = _T_1025 ^ (* src = "crypto_accelerator.v:7298" *) _T_1071;
  assign _T_1081 = _T_1065 ^ (* src = "crypto_accelerator.v:7299" *) _T_1077;
  assign _T_1083 = _T_1043 ^ (* src = "crypto_accelerator.v:7300" *) _T_1059;
  assign _T_1085 = _T_1027 ^ (* src = "crypto_accelerator.v:7301" *) _T_1033;
  assign _T_1087 = _T_1063 ^ (* src = "crypto_accelerator.v:7302" *) _T_1085;
  assign _T_1089 = _T_1055 ^ (* src = "crypto_accelerator.v:7303" *) _T_1081;
  assign _T_1091 = _T_1051 ^ (* src = "crypto_accelerator.v:7304" *) _T_1073;
  assign _T_1093 = _T_1065 ^ (* src = "crypto_accelerator.v:7305" *) _T_1075;
  assign _T_1094 = _T_1061 ^ (* src = "crypto_accelerator.v:7306" *) _T_1087;
  assign _T_1095 = _T_1089 ^ (* src = "crypto_accelerator.v:7307" *) _T_1091;
  assign _T_1098 = _T_1031 ^ (* src = "crypto_accelerator.v:7309" *) _T_1057;
  assign _T_1099 = _T_1069 ^ (* src = "crypto_accelerator.v:7310" *) _T_1071;
  assign _T_1100 = _T_1079 ^ (* src = "crypto_accelerator.v:7311" *) _T_1098;
  assign _T_1102 = _T_1029 ^ (* src = "crypto_accelerator.v:7312" *) _T_1045;
  assign _T_1104 = _T_1067 ^ (* src = "crypto_accelerator.v:7313" *) _T_1083;
  assign _T_1105 = _T_1069 ^ (* src = "crypto_accelerator.v:7314" *) _T_1093;
  assign _T_1108 = _T_1037 ^ (* src = "crypto_accelerator.v:7316" *) _T_1075;
  assign _T_1110 = _T_1102 ^ (* src = "crypto_accelerator.v:7317" *) _T_1108;
  assign _T_1112 = _T_1029 ^ (* src = "crypto_accelerator.v:7318" *) _T_1073;
  assign _T_1113 = _T_1061 ^ (* src = "crypto_accelerator.v:7319" *) _T_1110;
  assign _T_1116 = _T_1081 ^ (* src = "crypto_accelerator.v:7321" *) _T_1104;
  assign _T_1117 = _T_1061 ^ (* src = "crypto_accelerator.v:7322" *) _T_1116;
  assign _T_1119 = _T_1071 ^ (* src = "crypto_accelerator.v:7323" *) _T_1112;
  assign _T_1120 = _T_1061 ^ (* src = "crypto_accelerator.v:7324" *) _T_1119;
  assign _T_1139 = _T_1129_0_0 ^ (* src = "crypto_accelerator.v:7376" *) _T_1138;
  assign _T_1141 = _T_1139 ^ (* src = "crypto_accelerator.v:7378" *) _T_1140;
  assign _T_1143 = _T_1129_0_1 ^ (* src = "crypto_accelerator.v:7380" *) _T_1142;
  assign _T_1145 = _T_1129_0_2 ^ (* src = "crypto_accelerator.v:7382" *) _T_1144;
  assign _T_1147 = _T_1129_0_3 ^ (* src = "crypto_accelerator.v:7384" *) _T_1146;
  assign _T_1149 = _T_1129_1_0 ^ (* src = "crypto_accelerator.v:7385" *) _T_1141;
  assign _T_1150 = _T_1129_1_1 ^ (* src = "crypto_accelerator.v:7386" *) _T_1143;
  assign _T_1151 = _T_1129_1_2 ^ (* src = "crypto_accelerator.v:7387" *) _T_1145;
  assign _T_1152 = _T_1129_1_3 ^ (* src = "crypto_accelerator.v:7388" *) _T_1147;
  assign _T_1154 = _T_1129_2_0 ^ (* src = "crypto_accelerator.v:7389" *) _T_1149;
  assign _T_1155 = _T_1129_2_1 ^ (* src = "crypto_accelerator.v:7390" *) _T_1150;
  assign _T_1156 = _T_1129_2_2 ^ (* src = "crypto_accelerator.v:7391" *) _T_1151;
  assign _T_1157 = _T_1129_2_3 ^ (* src = "crypto_accelerator.v:7392" *) _T_1152;
  assign _T_1159 = _T_1129_3_0 ^ (* src = "crypto_accelerator.v:7393" *) _T_1154;
  assign _T_1160 = _T_1129_3_1 ^ (* src = "crypto_accelerator.v:7394" *) _T_1155;
  assign _T_1161 = _T_1129_3_2 ^ (* src = "crypto_accelerator.v:7395" *) _T_1156;
  assign _T_1162 = _T_1129_3_3 ^ (* src = "crypto_accelerator.v:7396" *) _T_1157;
  (* src = "crypto_accelerator.v:7458" *)
  AesDecrypt dec (
    .clock(clock),
    .io_aes256(io_aes256),
    .io_dataIn(io_decDataIn),
    .io_dataOut(dec_io_dataOut),
    .io_dataValid(io_decDataValid),
    .io_ivIn(io_decIvIn),
    .io_ivOut(dec_io_ivOut),
    .io_keys_0_0_0(shreg_io_output_14[127:120]),
    .io_keys_0_0_1(shreg_io_output_14[119:112]),
    .io_keys_0_0_2(shreg_io_output_14[111:104]),
    .io_keys_0_0_3(shreg_io_output_14[103:96]),
    .io_keys_0_1_0(shreg_io_output_14[95:88]),
    .io_keys_0_1_1(shreg_io_output_14[87:80]),
    .io_keys_0_1_2(shreg_io_output_14[79:72]),
    .io_keys_0_1_3(shreg_io_output_14[71:64]),
    .io_keys_0_2_0(shreg_io_output_14[63:56]),
    .io_keys_0_2_1(shreg_io_output_14[55:48]),
    .io_keys_0_2_2(shreg_io_output_14[47:40]),
    .io_keys_0_2_3(shreg_io_output_14[39:32]),
    .io_keys_0_3_0(shreg_io_output_14[31:24]),
    .io_keys_0_3_1(shreg_io_output_14[23:16]),
    .io_keys_0_3_2(shreg_io_output_14[15:8]),
    .io_keys_0_3_3(shreg_io_output_14[7:0]),
    .io_keys_10_0_0(shreg_io_output_4[127:120]),
    .io_keys_10_0_1(shreg_io_output_4[119:112]),
    .io_keys_10_0_2(shreg_io_output_4[111:104]),
    .io_keys_10_0_3(shreg_io_output_4[103:96]),
    .io_keys_10_1_0(shreg_io_output_4[95:88]),
    .io_keys_10_1_1(shreg_io_output_4[87:80]),
    .io_keys_10_1_2(shreg_io_output_4[79:72]),
    .io_keys_10_1_3(shreg_io_output_4[71:64]),
    .io_keys_10_2_0(shreg_io_output_4[63:56]),
    .io_keys_10_2_1(shreg_io_output_4[55:48]),
    .io_keys_10_2_2(shreg_io_output_4[47:40]),
    .io_keys_10_2_3(shreg_io_output_4[39:32]),
    .io_keys_10_3_0(shreg_io_output_4[31:24]),
    .io_keys_10_3_1(shreg_io_output_4[23:16]),
    .io_keys_10_3_2(shreg_io_output_4[15:8]),
    .io_keys_10_3_3(shreg_io_output_4[7:0]),
    .io_keys_11_0_0(shreg_io_output_3[127:120]),
    .io_keys_11_0_1(shreg_io_output_3[119:112]),
    .io_keys_11_0_2(shreg_io_output_3[111:104]),
    .io_keys_11_0_3(shreg_io_output_3[103:96]),
    .io_keys_11_1_0(shreg_io_output_3[95:88]),
    .io_keys_11_1_1(shreg_io_output_3[87:80]),
    .io_keys_11_1_2(shreg_io_output_3[79:72]),
    .io_keys_11_1_3(shreg_io_output_3[71:64]),
    .io_keys_11_2_0(shreg_io_output_3[63:56]),
    .io_keys_11_2_1(shreg_io_output_3[55:48]),
    .io_keys_11_2_2(shreg_io_output_3[47:40]),
    .io_keys_11_2_3(shreg_io_output_3[39:32]),
    .io_keys_11_3_0(shreg_io_output_3[31:24]),
    .io_keys_11_3_1(shreg_io_output_3[23:16]),
    .io_keys_11_3_2(shreg_io_output_3[15:8]),
    .io_keys_11_3_3(shreg_io_output_3[7:0]),
    .io_keys_12_0_0(shreg_io_output_2[127:120]),
    .io_keys_12_0_1(shreg_io_output_2[119:112]),
    .io_keys_12_0_2(shreg_io_output_2[111:104]),
    .io_keys_12_0_3(shreg_io_output_2[103:96]),
    .io_keys_12_1_0(shreg_io_output_2[95:88]),
    .io_keys_12_1_1(shreg_io_output_2[87:80]),
    .io_keys_12_1_2(shreg_io_output_2[79:72]),
    .io_keys_12_1_3(shreg_io_output_2[71:64]),
    .io_keys_12_2_0(shreg_io_output_2[63:56]),
    .io_keys_12_2_1(shreg_io_output_2[55:48]),
    .io_keys_12_2_2(shreg_io_output_2[47:40]),
    .io_keys_12_2_3(shreg_io_output_2[39:32]),
    .io_keys_12_3_0(shreg_io_output_2[31:24]),
    .io_keys_12_3_1(shreg_io_output_2[23:16]),
    .io_keys_12_3_2(shreg_io_output_2[15:8]),
    .io_keys_12_3_3(shreg_io_output_2[7:0]),
    .io_keys_13_0_0(shreg_io_output_1[127:120]),
    .io_keys_13_0_1(shreg_io_output_1[119:112]),
    .io_keys_13_0_2(shreg_io_output_1[111:104]),
    .io_keys_13_0_3(shreg_io_output_1[103:96]),
    .io_keys_13_1_0(shreg_io_output_1[95:88]),
    .io_keys_13_1_1(shreg_io_output_1[87:80]),
    .io_keys_13_1_2(shreg_io_output_1[79:72]),
    .io_keys_13_1_3(shreg_io_output_1[71:64]),
    .io_keys_13_2_0(shreg_io_output_1[63:56]),
    .io_keys_13_2_1(shreg_io_output_1[55:48]),
    .io_keys_13_2_2(shreg_io_output_1[47:40]),
    .io_keys_13_2_3(shreg_io_output_1[39:32]),
    .io_keys_13_3_0(shreg_io_output_1[31:24]),
    .io_keys_13_3_1(shreg_io_output_1[23:16]),
    .io_keys_13_3_2(shreg_io_output_1[15:8]),
    .io_keys_13_3_3(shreg_io_output_1[7:0]),
    .io_keys_14_0_0(shreg_io_output_0[127:120]),
    .io_keys_14_0_1(shreg_io_output_0[119:112]),
    .io_keys_14_0_2(shreg_io_output_0[111:104]),
    .io_keys_14_0_3(shreg_io_output_0[103:96]),
    .io_keys_14_1_0(shreg_io_output_0[95:88]),
    .io_keys_14_1_1(shreg_io_output_0[87:80]),
    .io_keys_14_1_2(shreg_io_output_0[79:72]),
    .io_keys_14_1_3(shreg_io_output_0[71:64]),
    .io_keys_14_2_0(shreg_io_output_0[63:56]),
    .io_keys_14_2_1(shreg_io_output_0[55:48]),
    .io_keys_14_2_2(shreg_io_output_0[47:40]),
    .io_keys_14_2_3(shreg_io_output_0[39:32]),
    .io_keys_14_3_0(shreg_io_output_0[31:24]),
    .io_keys_14_3_1(shreg_io_output_0[23:16]),
    .io_keys_14_3_2(shreg_io_output_0[15:8]),
    .io_keys_14_3_3(shreg_io_output_0[7:0]),
    .io_keys_1_0_0(shreg_io_output_13[127:120]),
    .io_keys_1_0_1(shreg_io_output_13[119:112]),
    .io_keys_1_0_2(shreg_io_output_13[111:104]),
    .io_keys_1_0_3(shreg_io_output_13[103:96]),
    .io_keys_1_1_0(shreg_io_output_13[95:88]),
    .io_keys_1_1_1(shreg_io_output_13[87:80]),
    .io_keys_1_1_2(shreg_io_output_13[79:72]),
    .io_keys_1_1_3(shreg_io_output_13[71:64]),
    .io_keys_1_2_0(shreg_io_output_13[63:56]),
    .io_keys_1_2_1(shreg_io_output_13[55:48]),
    .io_keys_1_2_2(shreg_io_output_13[47:40]),
    .io_keys_1_2_3(shreg_io_output_13[39:32]),
    .io_keys_1_3_0(shreg_io_output_13[31:24]),
    .io_keys_1_3_1(shreg_io_output_13[23:16]),
    .io_keys_1_3_2(shreg_io_output_13[15:8]),
    .io_keys_1_3_3(shreg_io_output_13[7:0]),
    .io_keys_2_0_0(shreg_io_output_12[127:120]),
    .io_keys_2_0_1(shreg_io_output_12[119:112]),
    .io_keys_2_0_2(shreg_io_output_12[111:104]),
    .io_keys_2_0_3(shreg_io_output_12[103:96]),
    .io_keys_2_1_0(shreg_io_output_12[95:88]),
    .io_keys_2_1_1(shreg_io_output_12[87:80]),
    .io_keys_2_1_2(shreg_io_output_12[79:72]),
    .io_keys_2_1_3(shreg_io_output_12[71:64]),
    .io_keys_2_2_0(shreg_io_output_12[63:56]),
    .io_keys_2_2_1(shreg_io_output_12[55:48]),
    .io_keys_2_2_2(shreg_io_output_12[47:40]),
    .io_keys_2_2_3(shreg_io_output_12[39:32]),
    .io_keys_2_3_0(shreg_io_output_12[31:24]),
    .io_keys_2_3_1(shreg_io_output_12[23:16]),
    .io_keys_2_3_2(shreg_io_output_12[15:8]),
    .io_keys_2_3_3(shreg_io_output_12[7:0]),
    .io_keys_3_0_0(shreg_io_output_11[127:120]),
    .io_keys_3_0_1(shreg_io_output_11[119:112]),
    .io_keys_3_0_2(shreg_io_output_11[111:104]),
    .io_keys_3_0_3(shreg_io_output_11[103:96]),
    .io_keys_3_1_0(shreg_io_output_11[95:88]),
    .io_keys_3_1_1(shreg_io_output_11[87:80]),
    .io_keys_3_1_2(shreg_io_output_11[79:72]),
    .io_keys_3_1_3(shreg_io_output_11[71:64]),
    .io_keys_3_2_0(shreg_io_output_11[63:56]),
    .io_keys_3_2_1(shreg_io_output_11[55:48]),
    .io_keys_3_2_2(shreg_io_output_11[47:40]),
    .io_keys_3_2_3(shreg_io_output_11[39:32]),
    .io_keys_3_3_0(shreg_io_output_11[31:24]),
    .io_keys_3_3_1(shreg_io_output_11[23:16]),
    .io_keys_3_3_2(shreg_io_output_11[15:8]),
    .io_keys_3_3_3(shreg_io_output_11[7:0]),
    .io_keys_4_0_0(shreg_io_output_10[127:120]),
    .io_keys_4_0_1(shreg_io_output_10[119:112]),
    .io_keys_4_0_2(shreg_io_output_10[111:104]),
    .io_keys_4_0_3(shreg_io_output_10[103:96]),
    .io_keys_4_1_0(shreg_io_output_10[95:88]),
    .io_keys_4_1_1(shreg_io_output_10[87:80]),
    .io_keys_4_1_2(shreg_io_output_10[79:72]),
    .io_keys_4_1_3(shreg_io_output_10[71:64]),
    .io_keys_4_2_0(shreg_io_output_10[63:56]),
    .io_keys_4_2_1(shreg_io_output_10[55:48]),
    .io_keys_4_2_2(shreg_io_output_10[47:40]),
    .io_keys_4_2_3(shreg_io_output_10[39:32]),
    .io_keys_4_3_0(shreg_io_output_10[31:24]),
    .io_keys_4_3_1(shreg_io_output_10[23:16]),
    .io_keys_4_3_2(shreg_io_output_10[15:8]),
    .io_keys_4_3_3(shreg_io_output_10[7:0]),
    .io_keys_5_0_0(shreg_io_output_9[127:120]),
    .io_keys_5_0_1(shreg_io_output_9[119:112]),
    .io_keys_5_0_2(shreg_io_output_9[111:104]),
    .io_keys_5_0_3(shreg_io_output_9[103:96]),
    .io_keys_5_1_0(shreg_io_output_9[95:88]),
    .io_keys_5_1_1(shreg_io_output_9[87:80]),
    .io_keys_5_1_2(shreg_io_output_9[79:72]),
    .io_keys_5_1_3(shreg_io_output_9[71:64]),
    .io_keys_5_2_0(shreg_io_output_9[63:56]),
    .io_keys_5_2_1(shreg_io_output_9[55:48]),
    .io_keys_5_2_2(shreg_io_output_9[47:40]),
    .io_keys_5_2_3(shreg_io_output_9[39:32]),
    .io_keys_5_3_0(shreg_io_output_9[31:24]),
    .io_keys_5_3_1(shreg_io_output_9[23:16]),
    .io_keys_5_3_2(shreg_io_output_9[15:8]),
    .io_keys_5_3_3(shreg_io_output_9[7:0]),
    .io_keys_6_0_0(shreg_io_output_8[127:120]),
    .io_keys_6_0_1(shreg_io_output_8[119:112]),
    .io_keys_6_0_2(shreg_io_output_8[111:104]),
    .io_keys_6_0_3(shreg_io_output_8[103:96]),
    .io_keys_6_1_0(shreg_io_output_8[95:88]),
    .io_keys_6_1_1(shreg_io_output_8[87:80]),
    .io_keys_6_1_2(shreg_io_output_8[79:72]),
    .io_keys_6_1_3(shreg_io_output_8[71:64]),
    .io_keys_6_2_0(shreg_io_output_8[63:56]),
    .io_keys_6_2_1(shreg_io_output_8[55:48]),
    .io_keys_6_2_2(shreg_io_output_8[47:40]),
    .io_keys_6_2_3(shreg_io_output_8[39:32]),
    .io_keys_6_3_0(shreg_io_output_8[31:24]),
    .io_keys_6_3_1(shreg_io_output_8[23:16]),
    .io_keys_6_3_2(shreg_io_output_8[15:8]),
    .io_keys_6_3_3(shreg_io_output_8[7:0]),
    .io_keys_7_0_0(shreg_io_output_7[127:120]),
    .io_keys_7_0_1(shreg_io_output_7[119:112]),
    .io_keys_7_0_2(shreg_io_output_7[111:104]),
    .io_keys_7_0_3(shreg_io_output_7[103:96]),
    .io_keys_7_1_0(shreg_io_output_7[95:88]),
    .io_keys_7_1_1(shreg_io_output_7[87:80]),
    .io_keys_7_1_2(shreg_io_output_7[79:72]),
    .io_keys_7_1_3(shreg_io_output_7[71:64]),
    .io_keys_7_2_0(shreg_io_output_7[63:56]),
    .io_keys_7_2_1(shreg_io_output_7[55:48]),
    .io_keys_7_2_2(shreg_io_output_7[47:40]),
    .io_keys_7_2_3(shreg_io_output_7[39:32]),
    .io_keys_7_3_0(shreg_io_output_7[31:24]),
    .io_keys_7_3_1(shreg_io_output_7[23:16]),
    .io_keys_7_3_2(shreg_io_output_7[15:8]),
    .io_keys_7_3_3(shreg_io_output_7[7:0]),
    .io_keys_8_0_0(shreg_io_output_6[127:120]),
    .io_keys_8_0_1(shreg_io_output_6[119:112]),
    .io_keys_8_0_2(shreg_io_output_6[111:104]),
    .io_keys_8_0_3(shreg_io_output_6[103:96]),
    .io_keys_8_1_0(shreg_io_output_6[95:88]),
    .io_keys_8_1_1(shreg_io_output_6[87:80]),
    .io_keys_8_1_2(shreg_io_output_6[79:72]),
    .io_keys_8_1_3(shreg_io_output_6[71:64]),
    .io_keys_8_2_0(shreg_io_output_6[63:56]),
    .io_keys_8_2_1(shreg_io_output_6[55:48]),
    .io_keys_8_2_2(shreg_io_output_6[47:40]),
    .io_keys_8_2_3(shreg_io_output_6[39:32]),
    .io_keys_8_3_0(shreg_io_output_6[31:24]),
    .io_keys_8_3_1(shreg_io_output_6[23:16]),
    .io_keys_8_3_2(shreg_io_output_6[15:8]),
    .io_keys_8_3_3(shreg_io_output_6[7:0]),
    .io_keys_9_0_0(shreg_io_output_5[127:120]),
    .io_keys_9_0_1(shreg_io_output_5[119:112]),
    .io_keys_9_0_2(shreg_io_output_5[111:104]),
    .io_keys_9_0_3(shreg_io_output_5[103:96]),
    .io_keys_9_1_0(shreg_io_output_5[95:88]),
    .io_keys_9_1_1(shreg_io_output_5[87:80]),
    .io_keys_9_1_2(shreg_io_output_5[79:72]),
    .io_keys_9_1_3(shreg_io_output_5[71:64]),
    .io_keys_9_2_0(shreg_io_output_5[63:56]),
    .io_keys_9_2_1(shreg_io_output_5[55:48]),
    .io_keys_9_2_2(shreg_io_output_5[47:40]),
    .io_keys_9_2_3(shreg_io_output_5[39:32]),
    .io_keys_9_3_0(shreg_io_output_5[31:24]),
    .io_keys_9_3_1(shreg_io_output_5[23:16]),
    .io_keys_9_3_2(shreg_io_output_5[15:8]),
    .io_keys_9_3_3(shreg_io_output_5[7:0]),
    .io_outputValid(dec_io_outputValid),
    .io_ready(dec_io_ready),
    .io_shift(dec_io_shift),
    .io_shiftCyc(dec_io_shiftCyc),
    .io_shiftRev(dec_io_shiftRev),
    .reset(reset)
  );
  (* src = "crypto_accelerator.v:7428" *)
  AesEncrypt enc (
    .clock(clock),
    .io_aes256(io_aes256),
    .io_dataIn(io_encDataIn),
    .io_dataOut(enc_io_dataOut),
    .io_dataValid(io_encDataValid),
    .io_ivIn(io_encIvIn),
    .io_ivOut(enc_io_ivOut),
    .io_keys_0_0_0(shreg_io_output_14[127:120]),
    .io_keys_0_0_1(shreg_io_output_14[119:112]),
    .io_keys_0_0_2(shreg_io_output_14[111:104]),
    .io_keys_0_0_3(shreg_io_output_14[103:96]),
    .io_keys_0_1_0(shreg_io_output_14[95:88]),
    .io_keys_0_1_1(shreg_io_output_14[87:80]),
    .io_keys_0_1_2(shreg_io_output_14[79:72]),
    .io_keys_0_1_3(shreg_io_output_14[71:64]),
    .io_keys_0_2_0(shreg_io_output_14[63:56]),
    .io_keys_0_2_1(shreg_io_output_14[55:48]),
    .io_keys_0_2_2(shreg_io_output_14[47:40]),
    .io_keys_0_2_3(shreg_io_output_14[39:32]),
    .io_keys_0_3_0(shreg_io_output_14[31:24]),
    .io_keys_0_3_1(shreg_io_output_14[23:16]),
    .io_keys_0_3_2(shreg_io_output_14[15:8]),
    .io_keys_0_3_3(shreg_io_output_14[7:0]),
    .io_outputValid(enc_io_outputValid),
    .io_ready(enc_io_ready),
    .io_shift(enc_io_shift),
    .io_shiftCyc(enc_io_shiftCyc),
    .reset(reset)
  );
  (* src = "crypto_accelerator.v:7405" *)
  ShiftRegister shreg (
    .clock(clock),
    .io_cyc(shreg_io_cyc),
    .io_enable(shreg_io_enable),
    .io_input(shreg_io_input),
    .io_output_0(shreg_io_output_0),
    .io_output_1(shreg_io_output_1),
    .io_output_10(shreg_io_output_10),
    .io_output_11(shreg_io_output_11),
    .io_output_12(shreg_io_output_12),
    .io_output_13(shreg_io_output_13),
    .io_output_14(shreg_io_output_14),
    .io_output_2(shreg_io_output_2),
    .io_output_3(shreg_io_output_3),
    .io_output_4(shreg_io_output_4),
    .io_output_5(shreg_io_output_5),
    .io_output_6(shreg_io_output_6),
    .io_output_7(shreg_io_output_7),
    .io_output_8(shreg_io_output_8),
    .io_output_9(shreg_io_output_9),
    .io_rev(dec_io_shiftRev),
    .io_tap(io_aes256)
  );
  assign _T_1128 = { _T_1094, _T_1121, _T_1096, _T_1099, _T_1100, _T_1117, _T_1114, _T_1106 };
  assign _T_1170 = { _T_1154, _T_1155, _T_1156, _T_1157, _T_1159, _T_1160, _T_1161, _T_1162 };
  assign _T_1178 = { _T_1141, _T_1143, _T_1145, _T_1147, _T_1149, _T_1150, _T_1151, _T_1152, _T_1154, _T_1155, _T_1156, _T_1157, _T_1159, _T_1160, _T_1161, _T_1162 };
  assign _T_321 = { _T_287, _T_314, _T_289, _T_292, _T_293, _T_310, _T_307, _T_299 };
  assign _T_5 = _GEN_42;
  assign _T_590 = { _T_556, _T_583, _T_558, _T_561, _T_562, _T_579, _T_576, _T_568 };
  assign _T_859 = { _T_825, _T_852, _T_827, _T_830, _T_831, _T_848, _T_845, _T_837 };
  assign dec_clock = clock;
  assign dec_io_aes256 = io_aes256;
  assign dec_io_dataIn = io_decDataIn;
  assign dec_io_dataValid = io_decDataValid;
  assign dec_io_ivIn = io_decIvIn;
  assign dec_io_keys_0_0_0 = shreg_io_output_14[127:120];
  assign dec_io_keys_0_0_1 = shreg_io_output_14[119:112];
  assign dec_io_keys_0_0_2 = shreg_io_output_14[111:104];
  assign dec_io_keys_0_0_3 = shreg_io_output_14[103:96];
  assign dec_io_keys_0_1_0 = shreg_io_output_14[95:88];
  assign dec_io_keys_0_1_1 = shreg_io_output_14[87:80];
  assign dec_io_keys_0_1_2 = shreg_io_output_14[79:72];
  assign dec_io_keys_0_1_3 = shreg_io_output_14[71:64];
  assign dec_io_keys_0_2_0 = shreg_io_output_14[63:56];
  assign dec_io_keys_0_2_1 = shreg_io_output_14[55:48];
  assign dec_io_keys_0_2_2 = shreg_io_output_14[47:40];
  assign dec_io_keys_0_2_3 = shreg_io_output_14[39:32];
  assign dec_io_keys_0_3_0 = shreg_io_output_14[31:24];
  assign dec_io_keys_0_3_1 = shreg_io_output_14[23:16];
  assign dec_io_keys_0_3_2 = shreg_io_output_14[15:8];
  assign dec_io_keys_0_3_3 = shreg_io_output_14[7:0];
  assign dec_io_keys_10_0_0 = shreg_io_output_4[127:120];
  assign dec_io_keys_10_0_1 = shreg_io_output_4[119:112];
  assign dec_io_keys_10_0_2 = shreg_io_output_4[111:104];
  assign dec_io_keys_10_0_3 = shreg_io_output_4[103:96];
  assign dec_io_keys_10_1_0 = shreg_io_output_4[95:88];
  assign dec_io_keys_10_1_1 = shreg_io_output_4[87:80];
  assign dec_io_keys_10_1_2 = shreg_io_output_4[79:72];
  assign dec_io_keys_10_1_3 = shreg_io_output_4[71:64];
  assign dec_io_keys_10_2_0 = shreg_io_output_4[63:56];
  assign dec_io_keys_10_2_1 = shreg_io_output_4[55:48];
  assign dec_io_keys_10_2_2 = shreg_io_output_4[47:40];
  assign dec_io_keys_10_2_3 = shreg_io_output_4[39:32];
  assign dec_io_keys_10_3_0 = shreg_io_output_4[31:24];
  assign dec_io_keys_10_3_1 = shreg_io_output_4[23:16];
  assign dec_io_keys_10_3_2 = shreg_io_output_4[15:8];
  assign dec_io_keys_10_3_3 = shreg_io_output_4[7:0];
  assign dec_io_keys_11_0_0 = shreg_io_output_3[127:120];
  assign dec_io_keys_11_0_1 = shreg_io_output_3[119:112];
  assign dec_io_keys_11_0_2 = shreg_io_output_3[111:104];
  assign dec_io_keys_11_0_3 = shreg_io_output_3[103:96];
  assign dec_io_keys_11_1_0 = shreg_io_output_3[95:88];
  assign dec_io_keys_11_1_1 = shreg_io_output_3[87:80];
  assign dec_io_keys_11_1_2 = shreg_io_output_3[79:72];
  assign dec_io_keys_11_1_3 = shreg_io_output_3[71:64];
  assign dec_io_keys_11_2_0 = shreg_io_output_3[63:56];
  assign dec_io_keys_11_2_1 = shreg_io_output_3[55:48];
  assign dec_io_keys_11_2_2 = shreg_io_output_3[47:40];
  assign dec_io_keys_11_2_3 = shreg_io_output_3[39:32];
  assign dec_io_keys_11_3_0 = shreg_io_output_3[31:24];
  assign dec_io_keys_11_3_1 = shreg_io_output_3[23:16];
  assign dec_io_keys_11_3_2 = shreg_io_output_3[15:8];
  assign dec_io_keys_11_3_3 = shreg_io_output_3[7:0];
  assign dec_io_keys_12_0_0 = shreg_io_output_2[127:120];
  assign dec_io_keys_12_0_1 = shreg_io_output_2[119:112];
  assign dec_io_keys_12_0_2 = shreg_io_output_2[111:104];
  assign dec_io_keys_12_0_3 = shreg_io_output_2[103:96];
  assign dec_io_keys_12_1_0 = shreg_io_output_2[95:88];
  assign dec_io_keys_12_1_1 = shreg_io_output_2[87:80];
  assign dec_io_keys_12_1_2 = shreg_io_output_2[79:72];
  assign dec_io_keys_12_1_3 = shreg_io_output_2[71:64];
  assign dec_io_keys_12_2_0 = shreg_io_output_2[63:56];
  assign dec_io_keys_12_2_1 = shreg_io_output_2[55:48];
  assign dec_io_keys_12_2_2 = shreg_io_output_2[47:40];
  assign dec_io_keys_12_2_3 = shreg_io_output_2[39:32];
  assign dec_io_keys_12_3_0 = shreg_io_output_2[31:24];
  assign dec_io_keys_12_3_1 = shreg_io_output_2[23:16];
  assign dec_io_keys_12_3_2 = shreg_io_output_2[15:8];
  assign dec_io_keys_12_3_3 = shreg_io_output_2[7:0];
  assign dec_io_keys_13_0_0 = shreg_io_output_1[127:120];
  assign dec_io_keys_13_0_1 = shreg_io_output_1[119:112];
  assign dec_io_keys_13_0_2 = shreg_io_output_1[111:104];
  assign dec_io_keys_13_0_3 = shreg_io_output_1[103:96];
  assign dec_io_keys_13_1_0 = shreg_io_output_1[95:88];
  assign dec_io_keys_13_1_1 = shreg_io_output_1[87:80];
  assign dec_io_keys_13_1_2 = shreg_io_output_1[79:72];
  assign dec_io_keys_13_1_3 = shreg_io_output_1[71:64];
  assign dec_io_keys_13_2_0 = shreg_io_output_1[63:56];
  assign dec_io_keys_13_2_1 = shreg_io_output_1[55:48];
  assign dec_io_keys_13_2_2 = shreg_io_output_1[47:40];
  assign dec_io_keys_13_2_3 = shreg_io_output_1[39:32];
  assign dec_io_keys_13_3_0 = shreg_io_output_1[31:24];
  assign dec_io_keys_13_3_1 = shreg_io_output_1[23:16];
  assign dec_io_keys_13_3_2 = shreg_io_output_1[15:8];
  assign dec_io_keys_13_3_3 = shreg_io_output_1[7:0];
  assign dec_io_keys_14_0_0 = shreg_io_output_0[127:120];
  assign dec_io_keys_14_0_1 = shreg_io_output_0[119:112];
  assign dec_io_keys_14_0_2 = shreg_io_output_0[111:104];
  assign dec_io_keys_14_0_3 = shreg_io_output_0[103:96];
  assign dec_io_keys_14_1_0 = shreg_io_output_0[95:88];
  assign dec_io_keys_14_1_1 = shreg_io_output_0[87:80];
  assign dec_io_keys_14_1_2 = shreg_io_output_0[79:72];
  assign dec_io_keys_14_1_3 = shreg_io_output_0[71:64];
  assign dec_io_keys_14_2_0 = shreg_io_output_0[63:56];
  assign dec_io_keys_14_2_1 = shreg_io_output_0[55:48];
  assign dec_io_keys_14_2_2 = shreg_io_output_0[47:40];
  assign dec_io_keys_14_2_3 = shreg_io_output_0[39:32];
  assign dec_io_keys_14_3_0 = shreg_io_output_0[31:24];
  assign dec_io_keys_14_3_1 = shreg_io_output_0[23:16];
  assign dec_io_keys_14_3_2 = shreg_io_output_0[15:8];
  assign dec_io_keys_14_3_3 = shreg_io_output_0[7:0];
  assign dec_io_keys_1_0_0 = shreg_io_output_13[127:120];
  assign dec_io_keys_1_0_1 = shreg_io_output_13[119:112];
  assign dec_io_keys_1_0_2 = shreg_io_output_13[111:104];
  assign dec_io_keys_1_0_3 = shreg_io_output_13[103:96];
  assign dec_io_keys_1_1_0 = shreg_io_output_13[95:88];
  assign dec_io_keys_1_1_1 = shreg_io_output_13[87:80];
  assign dec_io_keys_1_1_2 = shreg_io_output_13[79:72];
  assign dec_io_keys_1_1_3 = shreg_io_output_13[71:64];
  assign dec_io_keys_1_2_0 = shreg_io_output_13[63:56];
  assign dec_io_keys_1_2_1 = shreg_io_output_13[55:48];
  assign dec_io_keys_1_2_2 = shreg_io_output_13[47:40];
  assign dec_io_keys_1_2_3 = shreg_io_output_13[39:32];
  assign dec_io_keys_1_3_0 = shreg_io_output_13[31:24];
  assign dec_io_keys_1_3_1 = shreg_io_output_13[23:16];
  assign dec_io_keys_1_3_2 = shreg_io_output_13[15:8];
  assign dec_io_keys_1_3_3 = shreg_io_output_13[7:0];
  assign dec_io_keys_2_0_0 = shreg_io_output_12[127:120];
  assign dec_io_keys_2_0_1 = shreg_io_output_12[119:112];
  assign dec_io_keys_2_0_2 = shreg_io_output_12[111:104];
  assign dec_io_keys_2_0_3 = shreg_io_output_12[103:96];
  assign dec_io_keys_2_1_0 = shreg_io_output_12[95:88];
  assign dec_io_keys_2_1_1 = shreg_io_output_12[87:80];
  assign dec_io_keys_2_1_2 = shreg_io_output_12[79:72];
  assign dec_io_keys_2_1_3 = shreg_io_output_12[71:64];
  assign dec_io_keys_2_2_0 = shreg_io_output_12[63:56];
  assign dec_io_keys_2_2_1 = shreg_io_output_12[55:48];
  assign dec_io_keys_2_2_2 = shreg_io_output_12[47:40];
  assign dec_io_keys_2_2_3 = shreg_io_output_12[39:32];
  assign dec_io_keys_2_3_0 = shreg_io_output_12[31:24];
  assign dec_io_keys_2_3_1 = shreg_io_output_12[23:16];
  assign dec_io_keys_2_3_2 = shreg_io_output_12[15:8];
  assign dec_io_keys_2_3_3 = shreg_io_output_12[7:0];
  assign dec_io_keys_3_0_0 = shreg_io_output_11[127:120];
  assign dec_io_keys_3_0_1 = shreg_io_output_11[119:112];
  assign dec_io_keys_3_0_2 = shreg_io_output_11[111:104];
  assign dec_io_keys_3_0_3 = shreg_io_output_11[103:96];
  assign dec_io_keys_3_1_0 = shreg_io_output_11[95:88];
  assign dec_io_keys_3_1_1 = shreg_io_output_11[87:80];
  assign dec_io_keys_3_1_2 = shreg_io_output_11[79:72];
  assign dec_io_keys_3_1_3 = shreg_io_output_11[71:64];
  assign dec_io_keys_3_2_0 = shreg_io_output_11[63:56];
  assign dec_io_keys_3_2_1 = shreg_io_output_11[55:48];
  assign dec_io_keys_3_2_2 = shreg_io_output_11[47:40];
  assign dec_io_keys_3_2_3 = shreg_io_output_11[39:32];
  assign dec_io_keys_3_3_0 = shreg_io_output_11[31:24];
  assign dec_io_keys_3_3_1 = shreg_io_output_11[23:16];
  assign dec_io_keys_3_3_2 = shreg_io_output_11[15:8];
  assign dec_io_keys_3_3_3 = shreg_io_output_11[7:0];
  assign dec_io_keys_4_0_0 = shreg_io_output_10[127:120];
  assign dec_io_keys_4_0_1 = shreg_io_output_10[119:112];
  assign dec_io_keys_4_0_2 = shreg_io_output_10[111:104];
  assign dec_io_keys_4_0_3 = shreg_io_output_10[103:96];
  assign dec_io_keys_4_1_0 = shreg_io_output_10[95:88];
  assign dec_io_keys_4_1_1 = shreg_io_output_10[87:80];
  assign dec_io_keys_4_1_2 = shreg_io_output_10[79:72];
  assign dec_io_keys_4_1_3 = shreg_io_output_10[71:64];
  assign dec_io_keys_4_2_0 = shreg_io_output_10[63:56];
  assign dec_io_keys_4_2_1 = shreg_io_output_10[55:48];
  assign dec_io_keys_4_2_2 = shreg_io_output_10[47:40];
  assign dec_io_keys_4_2_3 = shreg_io_output_10[39:32];
  assign dec_io_keys_4_3_0 = shreg_io_output_10[31:24];
  assign dec_io_keys_4_3_1 = shreg_io_output_10[23:16];
  assign dec_io_keys_4_3_2 = shreg_io_output_10[15:8];
  assign dec_io_keys_4_3_3 = shreg_io_output_10[7:0];
  assign dec_io_keys_5_0_0 = shreg_io_output_9[127:120];
  assign dec_io_keys_5_0_1 = shreg_io_output_9[119:112];
  assign dec_io_keys_5_0_2 = shreg_io_output_9[111:104];
  assign dec_io_keys_5_0_3 = shreg_io_output_9[103:96];
  assign dec_io_keys_5_1_0 = shreg_io_output_9[95:88];
  assign dec_io_keys_5_1_1 = shreg_io_output_9[87:80];
  assign dec_io_keys_5_1_2 = shreg_io_output_9[79:72];
  assign dec_io_keys_5_1_3 = shreg_io_output_9[71:64];
  assign dec_io_keys_5_2_0 = shreg_io_output_9[63:56];
  assign dec_io_keys_5_2_1 = shreg_io_output_9[55:48];
  assign dec_io_keys_5_2_2 = shreg_io_output_9[47:40];
  assign dec_io_keys_5_2_3 = shreg_io_output_9[39:32];
  assign dec_io_keys_5_3_0 = shreg_io_output_9[31:24];
  assign dec_io_keys_5_3_1 = shreg_io_output_9[23:16];
  assign dec_io_keys_5_3_2 = shreg_io_output_9[15:8];
  assign dec_io_keys_5_3_3 = shreg_io_output_9[7:0];
  assign dec_io_keys_6_0_0 = shreg_io_output_8[127:120];
  assign dec_io_keys_6_0_1 = shreg_io_output_8[119:112];
  assign dec_io_keys_6_0_2 = shreg_io_output_8[111:104];
  assign dec_io_keys_6_0_3 = shreg_io_output_8[103:96];
  assign dec_io_keys_6_1_0 = shreg_io_output_8[95:88];
  assign dec_io_keys_6_1_1 = shreg_io_output_8[87:80];
  assign dec_io_keys_6_1_2 = shreg_io_output_8[79:72];
  assign dec_io_keys_6_1_3 = shreg_io_output_8[71:64];
  assign dec_io_keys_6_2_0 = shreg_io_output_8[63:56];
  assign dec_io_keys_6_2_1 = shreg_io_output_8[55:48];
  assign dec_io_keys_6_2_2 = shreg_io_output_8[47:40];
  assign dec_io_keys_6_2_3 = shreg_io_output_8[39:32];
  assign dec_io_keys_6_3_0 = shreg_io_output_8[31:24];
  assign dec_io_keys_6_3_1 = shreg_io_output_8[23:16];
  assign dec_io_keys_6_3_2 = shreg_io_output_8[15:8];
  assign dec_io_keys_6_3_3 = shreg_io_output_8[7:0];
  assign dec_io_keys_7_0_0 = shreg_io_output_7[127:120];
  assign dec_io_keys_7_0_1 = shreg_io_output_7[119:112];
  assign dec_io_keys_7_0_2 = shreg_io_output_7[111:104];
  assign dec_io_keys_7_0_3 = shreg_io_output_7[103:96];
  assign dec_io_keys_7_1_0 = shreg_io_output_7[95:88];
  assign dec_io_keys_7_1_1 = shreg_io_output_7[87:80];
  assign dec_io_keys_7_1_2 = shreg_io_output_7[79:72];
  assign dec_io_keys_7_1_3 = shreg_io_output_7[71:64];
  assign dec_io_keys_7_2_0 = shreg_io_output_7[63:56];
  assign dec_io_keys_7_2_1 = shreg_io_output_7[55:48];
  assign dec_io_keys_7_2_2 = shreg_io_output_7[47:40];
  assign dec_io_keys_7_2_3 = shreg_io_output_7[39:32];
  assign dec_io_keys_7_3_0 = shreg_io_output_7[31:24];
  assign dec_io_keys_7_3_1 = shreg_io_output_7[23:16];
  assign dec_io_keys_7_3_2 = shreg_io_output_7[15:8];
  assign dec_io_keys_7_3_3 = shreg_io_output_7[7:0];
  assign dec_io_keys_8_0_0 = shreg_io_output_6[127:120];
  assign dec_io_keys_8_0_1 = shreg_io_output_6[119:112];
  assign dec_io_keys_8_0_2 = shreg_io_output_6[111:104];
  assign dec_io_keys_8_0_3 = shreg_io_output_6[103:96];
  assign dec_io_keys_8_1_0 = shreg_io_output_6[95:88];
  assign dec_io_keys_8_1_1 = shreg_io_output_6[87:80];
  assign dec_io_keys_8_1_2 = shreg_io_output_6[79:72];
  assign dec_io_keys_8_1_3 = shreg_io_output_6[71:64];
  assign dec_io_keys_8_2_0 = shreg_io_output_6[63:56];
  assign dec_io_keys_8_2_1 = shreg_io_output_6[55:48];
  assign dec_io_keys_8_2_2 = shreg_io_output_6[47:40];
  assign dec_io_keys_8_2_3 = shreg_io_output_6[39:32];
  assign dec_io_keys_8_3_0 = shreg_io_output_6[31:24];
  assign dec_io_keys_8_3_1 = shreg_io_output_6[23:16];
  assign dec_io_keys_8_3_2 = shreg_io_output_6[15:8];
  assign dec_io_keys_8_3_3 = shreg_io_output_6[7:0];
  assign dec_io_keys_9_0_0 = shreg_io_output_5[127:120];
  assign dec_io_keys_9_0_1 = shreg_io_output_5[119:112];
  assign dec_io_keys_9_0_2 = shreg_io_output_5[111:104];
  assign dec_io_keys_9_0_3 = shreg_io_output_5[103:96];
  assign dec_io_keys_9_1_0 = shreg_io_output_5[95:88];
  assign dec_io_keys_9_1_1 = shreg_io_output_5[87:80];
  assign dec_io_keys_9_1_2 = shreg_io_output_5[79:72];
  assign dec_io_keys_9_1_3 = shreg_io_output_5[71:64];
  assign dec_io_keys_9_2_0 = shreg_io_output_5[63:56];
  assign dec_io_keys_9_2_1 = shreg_io_output_5[55:48];
  assign dec_io_keys_9_2_2 = shreg_io_output_5[47:40];
  assign dec_io_keys_9_2_3 = shreg_io_output_5[39:32];
  assign dec_io_keys_9_3_0 = shreg_io_output_5[31:24];
  assign dec_io_keys_9_3_1 = shreg_io_output_5[23:16];
  assign dec_io_keys_9_3_2 = shreg_io_output_5[15:8];
  assign dec_io_keys_9_3_3 = shreg_io_output_5[7:0];
  assign dec_reset = reset;
  assign enc_clock = clock;
  assign enc_io_aes256 = io_aes256;
  assign enc_io_dataIn = io_encDataIn;
  assign enc_io_dataValid = io_encDataValid;
  assign enc_io_ivIn = io_encIvIn;
  assign enc_io_keys_0_0_0 = shreg_io_output_14[127:120];
  assign enc_io_keys_0_0_1 = shreg_io_output_14[119:112];
  assign enc_io_keys_0_0_2 = shreg_io_output_14[111:104];
  assign enc_io_keys_0_0_3 = shreg_io_output_14[103:96];
  assign enc_io_keys_0_1_0 = shreg_io_output_14[95:88];
  assign enc_io_keys_0_1_1 = shreg_io_output_14[87:80];
  assign enc_io_keys_0_1_2 = shreg_io_output_14[79:72];
  assign enc_io_keys_0_1_3 = shreg_io_output_14[71:64];
  assign enc_io_keys_0_2_0 = shreg_io_output_14[63:56];
  assign enc_io_keys_0_2_1 = shreg_io_output_14[55:48];
  assign enc_io_keys_0_2_2 = shreg_io_output_14[47:40];
  assign enc_io_keys_0_2_3 = shreg_io_output_14[39:32];
  assign enc_io_keys_0_3_0 = shreg_io_output_14[31:24];
  assign enc_io_keys_0_3_1 = shreg_io_output_14[23:16];
  assign enc_io_keys_0_3_2 = shreg_io_output_14[15:8];
  assign enc_io_keys_0_3_3 = shreg_io_output_14[7:0];
  assign enc_reset = reset;
  assign io_decDataOut = dec_io_dataOut;
  assign io_decIvOut = dec_io_ivOut;
  assign io_decOutputValid = dec_io_outputValid;
  assign io_encDataOut = enc_io_dataOut;
  assign io_encIvOut = enc_io_ivOut;
  assign io_encOutputValid = enc_io_outputValid;
  assign shreg_clock = clock;
  assign shreg_io_rev = dec_io_shiftRev;
  assign shreg_io_tap = io_aes256;
endmodule
