module NV_NVDLA_CVIF_WRITE_cq(nvdla_core_clk, nvdla_core_rstn, cq_wr_prdy, cq_wr_pvld, cq_wr_thread_id, cq_wr_pd, cq_rd0_prdy, cq_rd0_pvld, cq_rd0_pd, cq_rd1_prdy, cq_rd1_pvld, cq_rd1_pd, cq_rd2_prdy, cq_rd2_pvld, cq_rd2_pd, cq_rd3_prdy, cq_rd3_pvld, cq_rd3_pd, cq_rd4_prdy, cq_rd4_pvld, cq_rd4_pd, pwrbus_ram_pd);
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2396" *)
  wire [8:0] _0000_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2396" *)
  wire _0001_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2492" *)
  wire [8:0] _0002_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2492" *)
  wire _0003_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2588" *)
  wire [8:0] _0004_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2588" *)
  wire _0005_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2684" *)
  wire [8:0] _0006_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2684" *)
  wire _0007_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2780" *)
  wire [8:0] _0008_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2780" *)
  wire _0009_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2065" *)
  wire [8:0] _0010_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2065" *)
  wire [8:0] _0011_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2065" *)
  wire [8:0] _0012_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2065" *)
  wire [8:0] _0013_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2065" *)
  wire [8:0] _0014_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1979" *)
  wire [4:0] _0015_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2828" *)
  wire [2:0] _0016_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:123" *)
  wire [8:0] _0017_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:176" *)
  wire [254:0] _0018_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0019_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0020_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0021_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0022_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0023_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2304" *)
  wire [7:0] _0024_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1979" *)
  wire _0025_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2336" *)
  wire [2:0] _0026_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2371" *)
  wire _0027_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2336" *)
  wire [2:0] _0028_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2371" *)
  wire _0029_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2336" *)
  wire [2:0] _0030_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2371" *)
  wire _0031_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2432" *)
  wire [2:0] _0032_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2467" *)
  wire _0033_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2432" *)
  wire [2:0] _0034_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2467" *)
  wire _0035_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2432" *)
  wire [2:0] _0036_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2467" *)
  wire _0037_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2528" *)
  wire [2:0] _0038_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2563" *)
  wire _0039_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2528" *)
  wire [2:0] _0040_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2563" *)
  wire _0041_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2528" *)
  wire [2:0] _0042_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2563" *)
  wire _0043_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2624" *)
  wire [2:0] _0044_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2659" *)
  wire _0045_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2624" *)
  wire [2:0] _0046_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2659" *)
  wire _0047_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2624" *)
  wire [2:0] _0048_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2659" *)
  wire _0049_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2720" *)
  wire [2:0] _0050_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2755" *)
  wire _0051_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2720" *)
  wire [2:0] _0052_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2755" *)
  wire _0053_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2720" *)
  wire [2:0] _0054_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2755" *)
  wire _0055_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2017" *)
  wire [4:0] _0056_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0057_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0058_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0059_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0060_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2142" *)
  wire [7:0] _0061_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2127" *)
  wire [4:0] _0062_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0063_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0064_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0065_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0066_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0067_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0068_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0069_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0070_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0071_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0072_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0073_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0074_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0075_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0076_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0077_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0078_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0079_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0080_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0081_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0082_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0083_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0084_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0085_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0086_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0087_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0088_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0089_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0090_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0091_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0092_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0093_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0094_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0095_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0096_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0097_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0098_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0099_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0100_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0101_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0102_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0103_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0104_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0105_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0106_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0107_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0108_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0109_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0110_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0111_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0112_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0113_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0114_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0115_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0116_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0117_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0118_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0119_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0120_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0121_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0122_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0123_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0124_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0125_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0126_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0127_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0128_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0129_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0130_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0131_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0132_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0133_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0134_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0135_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0136_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0137_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0138_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0139_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0140_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0141_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0142_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0143_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0144_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0145_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0146_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0147_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0148_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0149_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0150_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0151_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0152_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0153_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0154_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0155_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0156_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0157_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0158_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0159_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0160_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0161_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0162_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0163_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0164_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0165_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0166_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0167_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0168_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0169_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0170_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0171_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0172_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0173_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0174_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0175_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0176_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0177_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0178_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0179_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0180_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0181_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0182_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0183_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0184_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0185_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0186_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0187_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0188_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0189_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0190_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0191_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0192_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0193_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0194_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0195_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0196_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0197_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0198_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0199_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0200_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0201_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0202_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0203_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0204_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0205_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0206_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0207_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0208_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0209_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0210_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0211_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0212_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0213_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0214_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0215_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0216_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0217_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0218_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0219_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0220_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0221_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0222_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0223_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0224_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0225_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0226_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0227_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0228_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0229_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0230_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0231_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0232_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0233_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0234_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0235_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0236_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0237_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0238_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0239_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0240_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0241_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0242_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0243_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0244_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0245_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0246_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0247_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0248_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0249_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0250_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0251_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0252_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0253_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0254_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0255_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0256_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0257_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0258_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0259_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0260_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0261_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0262_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0263_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0264_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0265_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0266_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0267_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0268_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0269_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0270_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0271_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0272_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0273_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0274_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0275_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0276_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0277_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0278_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0279_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0280_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0281_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0282_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0283_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0284_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0285_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0286_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0287_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0288_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0289_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0290_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0291_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0292_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0293_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0294_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0295_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0296_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0297_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0298_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0299_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0300_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0301_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0302_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0303_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0304_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0305_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0306_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0307_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0308_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0309_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0310_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0311_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0312_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0313_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0314_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0315_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0316_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:191" *)
  wire _0317_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2051" *)
  wire [8:0] _0318_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2054" *)
  wire [8:0] _0319_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2057" *)
  wire [8:0] _0320_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2060" *)
  wire [8:0] _0321_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2063" *)
  wire [8:0] _0322_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:94" *)
  wire [8:0] _0323_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1000" *)
  wire _0324_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1003" *)
  wire _0325_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1005" *)
  wire _0326_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1008" *)
  wire _0327_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1010" *)
  wire _0328_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1013" *)
  wire _0329_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1015" *)
  wire _0330_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1018" *)
  wire _0331_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1020" *)
  wire _0332_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1023" *)
  wire _0333_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1025" *)
  wire _0334_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1028" *)
  wire _0335_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1030" *)
  wire _0336_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1033" *)
  wire _0337_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1035" *)
  wire _0338_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1038" *)
  wire _0339_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1040" *)
  wire _0340_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1043" *)
  wire _0341_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1045" *)
  wire _0342_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1048" *)
  wire _0343_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1050" *)
  wire _0344_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1053" *)
  wire _0345_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1055" *)
  wire _0346_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1058" *)
  wire _0347_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1060" *)
  wire _0348_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1063" *)
  wire _0349_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1065" *)
  wire _0350_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1068" *)
  wire _0351_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1070" *)
  wire _0352_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1073" *)
  wire _0353_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1075" *)
  wire _0354_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1078" *)
  wire _0355_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1080" *)
  wire _0356_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1083" *)
  wire _0357_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1085" *)
  wire _0358_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1088" *)
  wire _0359_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1090" *)
  wire _0360_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1093" *)
  wire _0361_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1095" *)
  wire _0362_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1098" *)
  wire _0363_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1100" *)
  wire _0364_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1103" *)
  wire _0365_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1105" *)
  wire _0366_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1108" *)
  wire _0367_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1110" *)
  wire _0368_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1113" *)
  wire _0369_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1115" *)
  wire _0370_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1118" *)
  wire _0371_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1120" *)
  wire _0372_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1123" *)
  wire _0373_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1125" *)
  wire _0374_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1128" *)
  wire _0375_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1130" *)
  wire _0376_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1133" *)
  wire _0377_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1135" *)
  wire _0378_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1138" *)
  wire _0379_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1140" *)
  wire _0380_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1143" *)
  wire _0381_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1145" *)
  wire _0382_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1148" *)
  wire _0383_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1150" *)
  wire _0384_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1153" *)
  wire _0385_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1155" *)
  wire _0386_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1158" *)
  wire _0387_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1160" *)
  wire _0388_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1163" *)
  wire _0389_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1165" *)
  wire _0390_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1168" *)
  wire _0391_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1170" *)
  wire _0392_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1173" *)
  wire _0393_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1175" *)
  wire _0394_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1178" *)
  wire _0395_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1180" *)
  wire _0396_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1183" *)
  wire _0397_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1185" *)
  wire _0398_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1188" *)
  wire _0399_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1190" *)
  wire _0400_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1193" *)
  wire _0401_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1195" *)
  wire _0402_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1198" *)
  wire _0403_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1200" *)
  wire _0404_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1203" *)
  wire _0405_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1205" *)
  wire _0406_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1208" *)
  wire _0407_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1210" *)
  wire _0408_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1213" *)
  wire _0409_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1215" *)
  wire _0410_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1218" *)
  wire _0411_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1220" *)
  wire _0412_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1223" *)
  wire _0413_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1225" *)
  wire _0414_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1228" *)
  wire _0415_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1230" *)
  wire _0416_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1233" *)
  wire _0417_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1235" *)
  wire _0418_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1238" *)
  wire _0419_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1240" *)
  wire _0420_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1243" *)
  wire _0421_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1245" *)
  wire _0422_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1248" *)
  wire _0423_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1250" *)
  wire _0424_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1253" *)
  wire _0425_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1255" *)
  wire _0426_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1258" *)
  wire _0427_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1260" *)
  wire _0428_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1263" *)
  wire _0429_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1265" *)
  wire _0430_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1268" *)
  wire _0431_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1270" *)
  wire _0432_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1273" *)
  wire _0433_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1275" *)
  wire _0434_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1278" *)
  wire _0435_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1280" *)
  wire _0436_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1283" *)
  wire _0437_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1285" *)
  wire _0438_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1288" *)
  wire _0439_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1290" *)
  wire _0440_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1293" *)
  wire _0441_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1295" *)
  wire _0442_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1298" *)
  wire _0443_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1300" *)
  wire _0444_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1303" *)
  wire _0445_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1305" *)
  wire _0446_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1308" *)
  wire _0447_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1310" *)
  wire _0448_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1313" *)
  wire _0449_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1315" *)
  wire _0450_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1318" *)
  wire _0451_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1320" *)
  wire _0452_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1323" *)
  wire _0453_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1325" *)
  wire _0454_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1328" *)
  wire _0455_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1330" *)
  wire _0456_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1333" *)
  wire _0457_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1335" *)
  wire _0458_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1338" *)
  wire _0459_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1340" *)
  wire _0460_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1343" *)
  wire _0461_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1345" *)
  wire _0462_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1348" *)
  wire _0463_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1350" *)
  wire _0464_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1353" *)
  wire _0465_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1355" *)
  wire _0466_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1358" *)
  wire _0467_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1360" *)
  wire _0468_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1363" *)
  wire _0469_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1365" *)
  wire _0470_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1368" *)
  wire _0471_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1370" *)
  wire _0472_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1373" *)
  wire _0473_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1375" *)
  wire _0474_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1378" *)
  wire _0475_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1380" *)
  wire _0476_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1383" *)
  wire _0477_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1385" *)
  wire _0478_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1388" *)
  wire _0479_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1390" *)
  wire _0480_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1393" *)
  wire _0481_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1395" *)
  wire _0482_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1398" *)
  wire _0483_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1400" *)
  wire _0484_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1403" *)
  wire _0485_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1405" *)
  wire _0486_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1408" *)
  wire _0487_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1410" *)
  wire _0488_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1413" *)
  wire _0489_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1415" *)
  wire _0490_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1418" *)
  wire _0491_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1420" *)
  wire _0492_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1423" *)
  wire _0493_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1425" *)
  wire _0494_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1428" *)
  wire _0495_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1430" *)
  wire _0496_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1433" *)
  wire _0497_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1435" *)
  wire _0498_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1438" *)
  wire _0499_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1440" *)
  wire _0500_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1443" *)
  wire _0501_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1445" *)
  wire _0502_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1448" *)
  wire _0503_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1450" *)
  wire _0504_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1453" *)
  wire _0505_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1455" *)
  wire _0506_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1458" *)
  wire _0507_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1460" *)
  wire _0508_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1463" *)
  wire _0509_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1465" *)
  wire _0510_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:193" *)
  wire _0511_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:195" *)
  wire _0512_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:198" *)
  wire _0513_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1985" *)
  wire _0514_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1986" *)
  wire _0515_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1987" *)
  wire _0516_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1988" *)
  wire _0517_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1989" *)
  wire _0518_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1999" *)
  wire _0519_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:200" *)
  wire _0520_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2000" *)
  wire _0521_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2001" *)
  wire _0522_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2002" *)
  wire _0523_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2003" *)
  wire _0524_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:203" *)
  wire _0525_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:205" *)
  wire _0526_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:208" *)
  wire _0527_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:210" *)
  wire _0528_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:213" *)
  wire _0529_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:215" *)
  wire _0530_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2152" *)
  wire _0531_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *)
  wire _0532_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2167" *)
  wire _0533_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *)
  wire _0534_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:218" *)
  wire _0535_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2182" *)
  wire _0536_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *)
  wire _0537_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2197" *)
  wire _0538_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *)
  wire _0539_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:220" *)
  wire _0540_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2212" *)
  wire _0541_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *)
  wire _0542_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:223" *)
  wire _0543_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:225" *)
  wire _0544_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:228" *)
  wire _0545_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:230" *)
  wire _0546_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:233" *)
  wire _0547_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:235" *)
  wire _0548_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:238" *)
  wire _0549_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *)
  wire _0550_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:240" *)
  wire _0551_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:243" *)
  wire _0552_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:245" *)
  wire _0553_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:248" *)
  wire _0554_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *)
  wire _0555_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:250" *)
  wire _0556_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:253" *)
  wire _0557_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:255" *)
  wire _0558_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:258" *)
  wire _0559_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *)
  wire _0560_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:260" *)
  wire _0561_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:263" *)
  wire _0562_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:265" *)
  wire _0563_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:268" *)
  wire _0564_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *)
  wire _0565_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:270" *)
  wire _0566_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:273" *)
  wire _0567_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:275" *)
  wire _0568_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *)
  wire _0569_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:278" *)
  wire _0570_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:280" *)
  wire _0571_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *)
  wire _0572_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *)
  wire _0573_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *)
  wire _0574_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *)
  wire _0575_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2806" *)
  wire _0576_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:283" *)
  wire _0577_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:285" *)
  wire _0578_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:288" *)
  wire _0579_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:290" *)
  wire _0580_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:293" *)
  wire _0581_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:295" *)
  wire _0582_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:298" *)
  wire _0583_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:300" *)
  wire _0584_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:303" *)
  wire _0585_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:305" *)
  wire _0586_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:308" *)
  wire _0587_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:310" *)
  wire _0588_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:313" *)
  wire _0589_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:315" *)
  wire _0590_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:318" *)
  wire _0591_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:320" *)
  wire _0592_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:323" *)
  wire _0593_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:325" *)
  wire _0594_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:328" *)
  wire _0595_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:330" *)
  wire _0596_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:333" *)
  wire _0597_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:335" *)
  wire _0598_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:338" *)
  wire _0599_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:340" *)
  wire _0600_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:343" *)
  wire _0601_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:345" *)
  wire _0602_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:348" *)
  wire _0603_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:350" *)
  wire _0604_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:353" *)
  wire _0605_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:355" *)
  wire _0606_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:358" *)
  wire _0607_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:360" *)
  wire _0608_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:363" *)
  wire _0609_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:365" *)
  wire _0610_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:368" *)
  wire _0611_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:370" *)
  wire _0612_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:373" *)
  wire _0613_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:375" *)
  wire _0614_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:378" *)
  wire _0615_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:380" *)
  wire _0616_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:383" *)
  wire _0617_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:385" *)
  wire _0618_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:388" *)
  wire _0619_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:390" *)
  wire _0620_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:393" *)
  wire _0621_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:395" *)
  wire _0622_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:398" *)
  wire _0623_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:400" *)
  wire _0624_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:403" *)
  wire _0625_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:405" *)
  wire _0626_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:408" *)
  wire _0627_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:410" *)
  wire _0628_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:413" *)
  wire _0629_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:415" *)
  wire _0630_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:418" *)
  wire _0631_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:420" *)
  wire _0632_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:423" *)
  wire _0633_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:425" *)
  wire _0634_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:428" *)
  wire _0635_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:430" *)
  wire _0636_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:433" *)
  wire _0637_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:435" *)
  wire _0638_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:438" *)
  wire _0639_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:440" *)
  wire _0640_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:443" *)
  wire _0641_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:445" *)
  wire _0642_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:448" *)
  wire _0643_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:450" *)
  wire _0644_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:453" *)
  wire _0645_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:455" *)
  wire _0646_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:458" *)
  wire _0647_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:460" *)
  wire _0648_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:463" *)
  wire _0649_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:465" *)
  wire _0650_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:468" *)
  wire _0651_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:470" *)
  wire _0652_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:473" *)
  wire _0653_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:475" *)
  wire _0654_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:478" *)
  wire _0655_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:480" *)
  wire _0656_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:483" *)
  wire _0657_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:485" *)
  wire _0658_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:488" *)
  wire _0659_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:490" *)
  wire _0660_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:493" *)
  wire _0661_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:495" *)
  wire _0662_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:498" *)
  wire _0663_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:500" *)
  wire _0664_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:503" *)
  wire _0665_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:505" *)
  wire _0666_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:508" *)
  wire _0667_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:510" *)
  wire _0668_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:513" *)
  wire _0669_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:515" *)
  wire _0670_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:518" *)
  wire _0671_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:520" *)
  wire _0672_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:523" *)
  wire _0673_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:525" *)
  wire _0674_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:528" *)
  wire _0675_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:530" *)
  wire _0676_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:533" *)
  wire _0677_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:535" *)
  wire _0678_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:538" *)
  wire _0679_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:540" *)
  wire _0680_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:543" *)
  wire _0681_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:545" *)
  wire _0682_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:548" *)
  wire _0683_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:550" *)
  wire _0684_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:553" *)
  wire _0685_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:555" *)
  wire _0686_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:558" *)
  wire _0687_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:560" *)
  wire _0688_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:563" *)
  wire _0689_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:565" *)
  wire _0690_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:568" *)
  wire _0691_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:570" *)
  wire _0692_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:573" *)
  wire _0693_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:575" *)
  wire _0694_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:578" *)
  wire _0695_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:580" *)
  wire _0696_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:583" *)
  wire _0697_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:585" *)
  wire _0698_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:588" *)
  wire _0699_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:590" *)
  wire _0700_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:593" *)
  wire _0701_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:595" *)
  wire _0702_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:598" *)
  wire _0703_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:600" *)
  wire _0704_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:603" *)
  wire _0705_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:605" *)
  wire _0706_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:608" *)
  wire _0707_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:610" *)
  wire _0708_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:613" *)
  wire _0709_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:615" *)
  wire _0710_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:618" *)
  wire _0711_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:620" *)
  wire _0712_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:623" *)
  wire _0713_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:625" *)
  wire _0714_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:628" *)
  wire _0715_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:630" *)
  wire _0716_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:633" *)
  wire _0717_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:635" *)
  wire _0718_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:638" *)
  wire _0719_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:640" *)
  wire _0720_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:643" *)
  wire _0721_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:645" *)
  wire _0722_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:648" *)
  wire _0723_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:650" *)
  wire _0724_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:653" *)
  wire _0725_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:655" *)
  wire _0726_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:658" *)
  wire _0727_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:660" *)
  wire _0728_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:663" *)
  wire _0729_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:665" *)
  wire _0730_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:668" *)
  wire _0731_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:670" *)
  wire _0732_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:673" *)
  wire _0733_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:675" *)
  wire _0734_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:678" *)
  wire _0735_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:680" *)
  wire _0736_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:683" *)
  wire _0737_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:685" *)
  wire _0738_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:688" *)
  wire _0739_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:690" *)
  wire _0740_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:693" *)
  wire _0741_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:695" *)
  wire _0742_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:698" *)
  wire _0743_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:700" *)
  wire _0744_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:703" *)
  wire _0745_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:705" *)
  wire _0746_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:708" *)
  wire _0747_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:710" *)
  wire _0748_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:713" *)
  wire _0749_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:715" *)
  wire _0750_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:718" *)
  wire _0751_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:720" *)
  wire _0752_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:723" *)
  wire _0753_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:725" *)
  wire _0754_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:728" *)
  wire _0755_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:730" *)
  wire _0756_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:733" *)
  wire _0757_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:735" *)
  wire _0758_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:738" *)
  wire _0759_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:740" *)
  wire _0760_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:743" *)
  wire _0761_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:745" *)
  wire _0762_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:748" *)
  wire _0763_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:750" *)
  wire _0764_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:753" *)
  wire _0765_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:755" *)
  wire _0766_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:758" *)
  wire _0767_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:760" *)
  wire _0768_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:763" *)
  wire _0769_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:765" *)
  wire _0770_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:768" *)
  wire _0771_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:770" *)
  wire _0772_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:773" *)
  wire _0773_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:775" *)
  wire _0774_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:778" *)
  wire _0775_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:780" *)
  wire _0776_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:783" *)
  wire _0777_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:785" *)
  wire _0778_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:788" *)
  wire _0779_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:790" *)
  wire _0780_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:793" *)
  wire _0781_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:795" *)
  wire _0782_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:798" *)
  wire _0783_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:800" *)
  wire _0784_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:803" *)
  wire _0785_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:805" *)
  wire _0786_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:808" *)
  wire _0787_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:810" *)
  wire _0788_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:813" *)
  wire _0789_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:815" *)
  wire _0790_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:818" *)
  wire _0791_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:820" *)
  wire _0792_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:823" *)
  wire _0793_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:825" *)
  wire _0794_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:828" *)
  wire _0795_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:830" *)
  wire _0796_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:833" *)
  wire _0797_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:835" *)
  wire _0798_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:838" *)
  wire _0799_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:840" *)
  wire _0800_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:843" *)
  wire _0801_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:845" *)
  wire _0802_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:848" *)
  wire _0803_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:850" *)
  wire _0804_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:853" *)
  wire _0805_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:855" *)
  wire _0806_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:858" *)
  wire _0807_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:860" *)
  wire _0808_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:863" *)
  wire _0809_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:865" *)
  wire _0810_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:868" *)
  wire _0811_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:870" *)
  wire _0812_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:873" *)
  wire _0813_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:875" *)
  wire _0814_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:878" *)
  wire _0815_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:880" *)
  wire _0816_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:883" *)
  wire _0817_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:885" *)
  wire _0818_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:888" *)
  wire _0819_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:890" *)
  wire _0820_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:893" *)
  wire _0821_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:895" *)
  wire _0822_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:898" *)
  wire _0823_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:900" *)
  wire _0824_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:903" *)
  wire _0825_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:905" *)
  wire _0826_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:908" *)
  wire _0827_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:910" *)
  wire _0828_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:913" *)
  wire _0829_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:915" *)
  wire _0830_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:918" *)
  wire _0831_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:920" *)
  wire _0832_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:923" *)
  wire _0833_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:925" *)
  wire _0834_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:928" *)
  wire _0835_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:930" *)
  wire _0836_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:933" *)
  wire _0837_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:935" *)
  wire _0838_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:938" *)
  wire _0839_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:940" *)
  wire _0840_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:943" *)
  wire _0841_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:945" *)
  wire _0842_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:948" *)
  wire _0843_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:950" *)
  wire _0844_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:953" *)
  wire _0845_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:955" *)
  wire _0846_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:958" *)
  wire _0847_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:960" *)
  wire _0848_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:963" *)
  wire _0849_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:965" *)
  wire _0850_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:968" *)
  wire _0851_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:970" *)
  wire _0852_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:973" *)
  wire _0853_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:975" *)
  wire _0854_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:978" *)
  wire _0855_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:980" *)
  wire _0856_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:983" *)
  wire _0857_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:985" *)
  wire _0858_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:988" *)
  wire _0859_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:990" *)
  wire _0860_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:993" *)
  wire _0861_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:995" *)
  wire _0862_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:998" *)
  wire _0863_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2122" *)
  wire _0864_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2123" *)
  wire _0865_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2124" *)
  wire _0866_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2125" *)
  wire _0867_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2126" *)
  wire _0868_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1000" *)
  wire _0869_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1003" *)
  wire _0870_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1005" *)
  wire _0871_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1008" *)
  wire _0872_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1010" *)
  wire _0873_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1013" *)
  wire _0874_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1015" *)
  wire _0875_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1018" *)
  wire _0876_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1020" *)
  wire _0877_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1023" *)
  wire _0878_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1025" *)
  wire _0879_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1028" *)
  wire _0880_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1030" *)
  wire _0881_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1033" *)
  wire _0882_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1035" *)
  wire _0883_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1038" *)
  wire _0884_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1040" *)
  wire _0885_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1043" *)
  wire _0886_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1045" *)
  wire _0887_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1048" *)
  wire _0888_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1050" *)
  wire _0889_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1053" *)
  wire _0890_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1055" *)
  wire _0891_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1058" *)
  wire _0892_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1060" *)
  wire _0893_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1063" *)
  wire _0894_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1065" *)
  wire _0895_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1068" *)
  wire _0896_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1070" *)
  wire _0897_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1073" *)
  wire _0898_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1075" *)
  wire _0899_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1078" *)
  wire _0900_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1080" *)
  wire _0901_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1083" *)
  wire _0902_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1085" *)
  wire _0903_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1088" *)
  wire _0904_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1090" *)
  wire _0905_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1093" *)
  wire _0906_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1095" *)
  wire _0907_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1098" *)
  wire _0908_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1100" *)
  wire _0909_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1103" *)
  wire _0910_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1105" *)
  wire _0911_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1108" *)
  wire _0912_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1110" *)
  wire _0913_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1113" *)
  wire _0914_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1115" *)
  wire _0915_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1118" *)
  wire _0916_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1120" *)
  wire _0917_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1123" *)
  wire _0918_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1125" *)
  wire _0919_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1128" *)
  wire _0920_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1130" *)
  wire _0921_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1133" *)
  wire _0922_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1135" *)
  wire _0923_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1138" *)
  wire _0924_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1140" *)
  wire _0925_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1143" *)
  wire _0926_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1145" *)
  wire _0927_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1148" *)
  wire _0928_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1150" *)
  wire _0929_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1153" *)
  wire _0930_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1155" *)
  wire _0931_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1158" *)
  wire _0932_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1160" *)
  wire _0933_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1163" *)
  wire _0934_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1165" *)
  wire _0935_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1168" *)
  wire _0936_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1170" *)
  wire _0937_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1173" *)
  wire _0938_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1175" *)
  wire _0939_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1178" *)
  wire _0940_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1180" *)
  wire _0941_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1183" *)
  wire _0942_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1185" *)
  wire _0943_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1188" *)
  wire _0944_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1190" *)
  wire _0945_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1193" *)
  wire _0946_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1195" *)
  wire _0947_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1198" *)
  wire _0948_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1200" *)
  wire _0949_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1203" *)
  wire _0950_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1205" *)
  wire _0951_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1208" *)
  wire _0952_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1210" *)
  wire _0953_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1213" *)
  wire _0954_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1215" *)
  wire _0955_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1218" *)
  wire _0956_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1220" *)
  wire _0957_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1223" *)
  wire _0958_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1225" *)
  wire _0959_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1228" *)
  wire _0960_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1230" *)
  wire _0961_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1233" *)
  wire _0962_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1235" *)
  wire _0963_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1238" *)
  wire _0964_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1240" *)
  wire _0965_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1243" *)
  wire _0966_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1245" *)
  wire _0967_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1248" *)
  wire _0968_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1250" *)
  wire _0969_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1253" *)
  wire _0970_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1255" *)
  wire _0971_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1258" *)
  wire _0972_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1260" *)
  wire _0973_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1263" *)
  wire _0974_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1265" *)
  wire _0975_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1268" *)
  wire _0976_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1270" *)
  wire _0977_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1273" *)
  wire _0978_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1275" *)
  wire _0979_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1278" *)
  wire _0980_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1280" *)
  wire _0981_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1283" *)
  wire _0982_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1285" *)
  wire _0983_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1288" *)
  wire _0984_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1290" *)
  wire _0985_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1293" *)
  wire _0986_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1295" *)
  wire _0987_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1298" *)
  wire _0988_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1300" *)
  wire _0989_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1303" *)
  wire _0990_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1305" *)
  wire _0991_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1308" *)
  wire _0992_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1310" *)
  wire _0993_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1313" *)
  wire _0994_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1315" *)
  wire _0995_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1318" *)
  wire _0996_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1320" *)
  wire _0997_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1323" *)
  wire _0998_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1325" *)
  wire _0999_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1328" *)
  wire _1000_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1330" *)
  wire _1001_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1333" *)
  wire _1002_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1335" *)
  wire _1003_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1338" *)
  wire _1004_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1340" *)
  wire _1005_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1343" *)
  wire _1006_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1345" *)
  wire _1007_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1348" *)
  wire _1008_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1350" *)
  wire _1009_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1353" *)
  wire _1010_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1355" *)
  wire _1011_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1358" *)
  wire _1012_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1360" *)
  wire _1013_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1363" *)
  wire _1014_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1365" *)
  wire _1015_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1368" *)
  wire _1016_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1370" *)
  wire _1017_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1373" *)
  wire _1018_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1375" *)
  wire _1019_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1378" *)
  wire _1020_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1380" *)
  wire _1021_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1383" *)
  wire _1022_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1385" *)
  wire _1023_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1388" *)
  wire _1024_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1390" *)
  wire _1025_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1393" *)
  wire _1026_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1395" *)
  wire _1027_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1398" *)
  wire _1028_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1400" *)
  wire _1029_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1403" *)
  wire _1030_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1405" *)
  wire _1031_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1408" *)
  wire _1032_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1410" *)
  wire _1033_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1413" *)
  wire _1034_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1415" *)
  wire _1035_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1418" *)
  wire _1036_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1420" *)
  wire _1037_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1423" *)
  wire _1038_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1425" *)
  wire _1039_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1428" *)
  wire _1040_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1430" *)
  wire _1041_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1433" *)
  wire _1042_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1435" *)
  wire _1043_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1438" *)
  wire _1044_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1440" *)
  wire _1045_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1443" *)
  wire _1046_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1445" *)
  wire _1047_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1448" *)
  wire _1048_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1450" *)
  wire _1049_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1453" *)
  wire _1050_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1455" *)
  wire _1051_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1458" *)
  wire _1052_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1460" *)
  wire _1053_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1463" *)
  wire _1054_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1465" *)
  wire _1055_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:193" *)
  wire _1056_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:195" *)
  wire _1057_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:198" *)
  wire _1058_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:200" *)
  wire _1059_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:203" *)
  wire _1060_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:205" *)
  wire _1061_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:208" *)
  wire _1062_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:210" *)
  wire _1063_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:213" *)
  wire _1064_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:215" *)
  wire _1065_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2152" *)
  wire _1066_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *)
  wire _1067_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *)
  wire _1068_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2167" *)
  wire _1069_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *)
  wire _1070_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *)
  wire _1071_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:218" *)
  wire _1072_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2182" *)
  wire _1073_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *)
  wire _1074_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *)
  wire _1075_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2197" *)
  wire _1076_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *)
  wire _1077_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *)
  wire _1078_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:220" *)
  wire _1079_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2212" *)
  wire _1080_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *)
  wire _1081_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *)
  wire _1082_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:223" *)
  wire _1083_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2244" *)
  wire _1084_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2245" *)
  wire _1085_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2246" *)
  wire _1086_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2247" *)
  wire _1087_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2248" *)
  wire _1088_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:225" *)
  wire _1089_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2256" *)
  wire _1090_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2257" *)
  wire _1091_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2258" *)
  wire _1092_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2259" *)
  wire _1093_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2260" *)
  wire _1094_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2268" *)
  wire _1095_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2269" *)
  wire _1096_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2270" *)
  wire _1097_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2271" *)
  wire _1098_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2272" *)
  wire _1099_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:228" *)
  wire _1100_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:230" *)
  wire _1101_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:233" *)
  wire _1102_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1103_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1104_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1105_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2339" *)
  wire _1106_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *)
  wire _1107_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *)
  wire _1108_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:235" *)
  wire _1109_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2351" *)
  wire _1110_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *)
  wire _1111_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *)
  wire _1112_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *)
  wire _1113_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *)
  wire _1114_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *)
  wire _1115_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:238" *)
  wire _1116_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2380" *)
  wire _1117_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *)
  wire _1118_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *)
  wire _1119_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *)
  wire _1120_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *)
  wire _1121_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1122_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1123_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1124_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:240" *)
  wire _1125_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:243" *)
  wire _1126_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1127_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1128_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1129_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2435" *)
  wire _1130_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *)
  wire _1131_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *)
  wire _1132_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2447" *)
  wire _1133_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:245" *)
  wire _1134_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *)
  wire _1135_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *)
  wire _1136_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *)
  wire _1137_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *)
  wire _1138_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *)
  wire _1139_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2476" *)
  wire _1140_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:248" *)
  wire _1141_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *)
  wire _1142_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *)
  wire _1143_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *)
  wire _1144_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *)
  wire _1145_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1146_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1147_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1148_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:250" *)
  wire _1149_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1150_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1151_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1152_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:253" *)
  wire _1153_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2531" *)
  wire _1154_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *)
  wire _1155_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *)
  wire _1156_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2543" *)
  wire _1157_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:255" *)
  wire _1158_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *)
  wire _1159_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *)
  wire _1160_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *)
  wire _1161_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *)
  wire _1162_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *)
  wire _1163_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2572" *)
  wire _1164_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:258" *)
  wire _1165_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *)
  wire _1166_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *)
  wire _1167_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *)
  wire _1168_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *)
  wire _1169_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1170_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1171_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1172_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:260" *)
  wire _1173_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1174_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1175_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1176_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2627" *)
  wire _1177_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:263" *)
  wire _1178_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *)
  wire _1179_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *)
  wire _1180_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2639" *)
  wire _1181_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *)
  wire _1182_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *)
  wire _1183_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *)
  wire _1184_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:265" *)
  wire _1185_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *)
  wire _1186_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *)
  wire _1187_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2668" *)
  wire _1188_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:268" *)
  wire _1189_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *)
  wire _1190_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *)
  wire _1191_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *)
  wire _1192_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *)
  wire _1193_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1194_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1195_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1196_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:270" *)
  wire _1197_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1198_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1199_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1200_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2723" *)
  wire _1201_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:273" *)
  wire _1202_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *)
  wire _1203_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *)
  wire _1204_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2735" *)
  wire _1205_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *)
  wire _1206_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *)
  wire _1207_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *)
  wire _1208_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:275" *)
  wire _1209_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *)
  wire _1210_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *)
  wire _1211_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2764" *)
  wire _1212_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *)
  wire _1213_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *)
  wire _1214_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *)
  wire _1215_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *)
  wire _1216_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1217_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1218_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1219_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:278" *)
  wire _1220_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:280" *)
  wire _1221_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *)
  wire _1222_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *)
  wire _1223_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *)
  wire _1224_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *)
  wire _1225_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *)
  wire _1226_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *)
  wire _1227_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *)
  wire _1228_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *)
  wire _1229_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *)
  wire _1230_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *)
  wire _1231_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *)
  wire _1232_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *)
  wire _1233_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *)
  wire _1234_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *)
  wire _1235_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *)
  wire _1236_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *)
  wire _1237_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *)
  wire _1238_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *)
  wire _1239_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *)
  wire _1240_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2812" *)
  wire _1241_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *)
  wire _1242_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *)
  wire _1243_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *)
  wire _1244_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *)
  wire _1245_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *)
  wire _1246_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *)
  wire _1247_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *)
  wire _1248_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2817" *)
  wire _1249_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2818" *)
  wire _1250_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2818" *)
  wire _1251_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *)
  wire _1252_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *)
  wire _1253_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *)
  wire _1254_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *)
  wire _1255_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2822" *)
  wire _1256_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2823" *)
  wire _1257_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2823" *)
  wire _1258_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *)
  wire _1259_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *)
  wire _1260_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *)
  wire _1261_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:283" *)
  wire _1262_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:285" *)
  wire _1263_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:288" *)
  wire _1264_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:290" *)
  wire _1265_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:293" *)
  wire _1266_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:295" *)
  wire _1267_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:298" *)
  wire _1268_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:300" *)
  wire _1269_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:303" *)
  wire _1270_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:305" *)
  wire _1271_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:308" *)
  wire _1272_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:310" *)
  wire _1273_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:313" *)
  wire _1274_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:315" *)
  wire _1275_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:318" *)
  wire _1276_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:320" *)
  wire _1277_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:323" *)
  wire _1278_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:325" *)
  wire _1279_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:328" *)
  wire _1280_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:330" *)
  wire _1281_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:333" *)
  wire _1282_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:335" *)
  wire _1283_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:338" *)
  wire _1284_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:340" *)
  wire _1285_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:343" *)
  wire _1286_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:345" *)
  wire _1287_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:348" *)
  wire _1288_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:350" *)
  wire _1289_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:353" *)
  wire _1290_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:355" *)
  wire _1291_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:358" *)
  wire _1292_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:360" *)
  wire _1293_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:363" *)
  wire _1294_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:365" *)
  wire _1295_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:368" *)
  wire _1296_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:370" *)
  wire _1297_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:373" *)
  wire _1298_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:375" *)
  wire _1299_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:378" *)
  wire _1300_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:380" *)
  wire _1301_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:383" *)
  wire _1302_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:385" *)
  wire _1303_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:388" *)
  wire _1304_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:390" *)
  wire _1305_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:393" *)
  wire _1306_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:395" *)
  wire _1307_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:398" *)
  wire _1308_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:400" *)
  wire _1309_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:403" *)
  wire _1310_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:405" *)
  wire _1311_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:408" *)
  wire _1312_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:410" *)
  wire _1313_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:413" *)
  wire _1314_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:415" *)
  wire _1315_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:418" *)
  wire _1316_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:420" *)
  wire _1317_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:423" *)
  wire _1318_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:425" *)
  wire _1319_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:428" *)
  wire _1320_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:430" *)
  wire _1321_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:433" *)
  wire _1322_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:435" *)
  wire _1323_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:438" *)
  wire _1324_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:440" *)
  wire _1325_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:443" *)
  wire _1326_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:445" *)
  wire _1327_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:448" *)
  wire _1328_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:450" *)
  wire _1329_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:453" *)
  wire _1330_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:455" *)
  wire _1331_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:458" *)
  wire _1332_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:460" *)
  wire _1333_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:463" *)
  wire _1334_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:465" *)
  wire _1335_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:468" *)
  wire _1336_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:470" *)
  wire _1337_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:473" *)
  wire _1338_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:475" *)
  wire _1339_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:478" *)
  wire _1340_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:480" *)
  wire _1341_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:483" *)
  wire _1342_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:485" *)
  wire _1343_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:488" *)
  wire _1344_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:490" *)
  wire _1345_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:493" *)
  wire _1346_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:495" *)
  wire _1347_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:498" *)
  wire _1348_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:500" *)
  wire _1349_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:503" *)
  wire _1350_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:505" *)
  wire _1351_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:508" *)
  wire _1352_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:510" *)
  wire _1353_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:513" *)
  wire _1354_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:515" *)
  wire _1355_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:518" *)
  wire _1356_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:520" *)
  wire _1357_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:523" *)
  wire _1358_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:525" *)
  wire _1359_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:528" *)
  wire _1360_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:530" *)
  wire _1361_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:533" *)
  wire _1362_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:535" *)
  wire _1363_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:538" *)
  wire _1364_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:540" *)
  wire _1365_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:543" *)
  wire _1366_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:545" *)
  wire _1367_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:548" *)
  wire _1368_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:550" *)
  wire _1369_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:553" *)
  wire _1370_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:555" *)
  wire _1371_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:558" *)
  wire _1372_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:560" *)
  wire _1373_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:563" *)
  wire _1374_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:565" *)
  wire _1375_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:568" *)
  wire _1376_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:570" *)
  wire _1377_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:573" *)
  wire _1378_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:575" *)
  wire _1379_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:578" *)
  wire _1380_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:580" *)
  wire _1381_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:583" *)
  wire _1382_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:585" *)
  wire _1383_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:588" *)
  wire _1384_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:590" *)
  wire _1385_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:593" *)
  wire _1386_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:595" *)
  wire _1387_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:598" *)
  wire _1388_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:600" *)
  wire _1389_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:603" *)
  wire _1390_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:605" *)
  wire _1391_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:608" *)
  wire _1392_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:610" *)
  wire _1393_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:613" *)
  wire _1394_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:615" *)
  wire _1395_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:618" *)
  wire _1396_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:620" *)
  wire _1397_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:623" *)
  wire _1398_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:625" *)
  wire _1399_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:628" *)
  wire _1400_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:630" *)
  wire _1401_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:633" *)
  wire _1402_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:635" *)
  wire _1403_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:638" *)
  wire _1404_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:640" *)
  wire _1405_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:643" *)
  wire _1406_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:645" *)
  wire _1407_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:648" *)
  wire _1408_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:650" *)
  wire _1409_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:653" *)
  wire _1410_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:655" *)
  wire _1411_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:658" *)
  wire _1412_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:660" *)
  wire _1413_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:663" *)
  wire _1414_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:665" *)
  wire _1415_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:668" *)
  wire _1416_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:670" *)
  wire _1417_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:673" *)
  wire _1418_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:675" *)
  wire _1419_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:678" *)
  wire _1420_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:680" *)
  wire _1421_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:683" *)
  wire _1422_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:685" *)
  wire _1423_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:688" *)
  wire _1424_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:690" *)
  wire _1425_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:693" *)
  wire _1426_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:695" *)
  wire _1427_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:698" *)
  wire _1428_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:700" *)
  wire _1429_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:703" *)
  wire _1430_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:705" *)
  wire _1431_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:708" *)
  wire _1432_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:710" *)
  wire _1433_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:713" *)
  wire _1434_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:715" *)
  wire _1435_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:718" *)
  wire _1436_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:720" *)
  wire _1437_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:723" *)
  wire _1438_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:725" *)
  wire _1439_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:728" *)
  wire _1440_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:730" *)
  wire _1441_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:733" *)
  wire _1442_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:735" *)
  wire _1443_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:738" *)
  wire _1444_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:740" *)
  wire _1445_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:743" *)
  wire _1446_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:745" *)
  wire _1447_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:748" *)
  wire _1448_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:750" *)
  wire _1449_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:753" *)
  wire _1450_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:755" *)
  wire _1451_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:758" *)
  wire _1452_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:760" *)
  wire _1453_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:763" *)
  wire _1454_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:765" *)
  wire _1455_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:768" *)
  wire _1456_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:770" *)
  wire _1457_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:773" *)
  wire _1458_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:775" *)
  wire _1459_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:778" *)
  wire _1460_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:780" *)
  wire _1461_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:783" *)
  wire _1462_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:785" *)
  wire _1463_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:788" *)
  wire _1464_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:790" *)
  wire _1465_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:793" *)
  wire _1466_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:795" *)
  wire _1467_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:798" *)
  wire _1468_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:800" *)
  wire _1469_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:803" *)
  wire _1470_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:805" *)
  wire _1471_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:808" *)
  wire _1472_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:810" *)
  wire _1473_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:813" *)
  wire _1474_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:815" *)
  wire _1475_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:818" *)
  wire _1476_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:820" *)
  wire _1477_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:823" *)
  wire _1478_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:825" *)
  wire _1479_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:828" *)
  wire _1480_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:830" *)
  wire _1481_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:833" *)
  wire _1482_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:835" *)
  wire _1483_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:838" *)
  wire _1484_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:840" *)
  wire _1485_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:843" *)
  wire _1486_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:845" *)
  wire _1487_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:848" *)
  wire _1488_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:850" *)
  wire _1489_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:853" *)
  wire _1490_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:855" *)
  wire _1491_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:858" *)
  wire _1492_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:860" *)
  wire _1493_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:863" *)
  wire _1494_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:865" *)
  wire _1495_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:868" *)
  wire _1496_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:870" *)
  wire _1497_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:873" *)
  wire _1498_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:875" *)
  wire _1499_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:878" *)
  wire _1500_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:880" *)
  wire _1501_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:883" *)
  wire _1502_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:885" *)
  wire _1503_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:888" *)
  wire _1504_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:890" *)
  wire _1505_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:893" *)
  wire _1506_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:895" *)
  wire _1507_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:898" *)
  wire _1508_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:900" *)
  wire _1509_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:903" *)
  wire _1510_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:905" *)
  wire _1511_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:908" *)
  wire _1512_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:910" *)
  wire _1513_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:913" *)
  wire _1514_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:915" *)
  wire _1515_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:918" *)
  wire _1516_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:920" *)
  wire _1517_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:923" *)
  wire _1518_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:925" *)
  wire _1519_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:928" *)
  wire _1520_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:930" *)
  wire _1521_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:933" *)
  wire _1522_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:935" *)
  wire _1523_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:938" *)
  wire _1524_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:940" *)
  wire _1525_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:943" *)
  wire _1526_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:945" *)
  wire _1527_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:948" *)
  wire _1528_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:950" *)
  wire _1529_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:953" *)
  wire _1530_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:955" *)
  wire _1531_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:958" *)
  wire _1532_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:960" *)
  wire _1533_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:963" *)
  wire _1534_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:965" *)
  wire _1535_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:968" *)
  wire _1536_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:970" *)
  wire _1537_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:973" *)
  wire _1538_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:975" *)
  wire _1539_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:978" *)
  wire _1540_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:980" *)
  wire _1541_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:983" *)
  wire _1542_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:985" *)
  wire _1543_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:988" *)
  wire _1544_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:990" *)
  wire _1545_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:993" *)
  wire _1546_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:995" *)
  wire _1547_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:998" *)
  wire _1548_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:140" *)
  wire _1549_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1550_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1551_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *)
  wire _1552_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *)
  wire _1553_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *)
  wire _1554_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *)
  wire _1555_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1556_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1557_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1558_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1559_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *)
  wire _1560_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *)
  wire _1561_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *)
  wire _1562_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *)
  wire _1563_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1564_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1565_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1566_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1567_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *)
  wire _1568_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *)
  wire _1569_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *)
  wire _1570_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *)
  wire _1571_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1572_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1573_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1574_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1575_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *)
  wire _1576_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *)
  wire _1577_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *)
  wire _1578_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *)
  wire _1579_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1580_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1581_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1582_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1583_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *)
  wire _1584_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *)
  wire _1585_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *)
  wire _1586_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *)
  wire _1587_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1588_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1589_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *)
  wire _1590_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *)
  wire _1591_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *)
  wire _1592_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *)
  wire _1593_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *)
  wire _1594_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:180" *)
  wire _1595_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *)
  wire _1596_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2131" *)
  wire _1597_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *)
  wire _1598_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *)
  wire _1599_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *)
  wire _1600_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *)
  wire _1601_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *)
  wire _1602_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1603_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *)
  wire _1604_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *)
  wire _1605_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *)
  wire _1606_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *)
  wire _1607_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *)
  wire _1608_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *)
  wire _1609_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *)
  wire _1610_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *)
  wire _1611_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *)
  wire _1612_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *)
  wire _1613_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *)
  wire _1614_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *)
  wire _1615_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *)
  wire _1616_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *)
  wire _1617_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1618_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *)
  wire _1619_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1620_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *)
  wire _1621_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *)
  wire _1622_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *)
  wire _1623_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *)
  wire _1624_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *)
  wire _1625_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *)
  wire _1626_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *)
  wire _1627_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *)
  wire _1628_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *)
  wire _1629_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *)
  wire _1630_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *)
  wire _1631_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *)
  wire _1632_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *)
  wire _1633_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *)
  wire _1634_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1635_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *)
  wire _1636_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1637_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *)
  wire _1638_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *)
  wire _1639_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *)
  wire _1640_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *)
  wire _1641_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *)
  wire _1642_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *)
  wire _1643_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *)
  wire _1644_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *)
  wire _1645_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *)
  wire _1646_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *)
  wire _1647_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *)
  wire _1648_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *)
  wire _1649_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *)
  wire _1650_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *)
  wire _1651_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1652_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *)
  wire _1653_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1654_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *)
  wire _1655_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *)
  wire _1656_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *)
  wire _1657_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *)
  wire _1658_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *)
  wire _1659_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *)
  wire _1660_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *)
  wire _1661_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *)
  wire _1662_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *)
  wire _1663_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *)
  wire _1664_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *)
  wire _1665_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *)
  wire _1666_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *)
  wire _1667_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *)
  wire _1668_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1669_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *)
  wire _1670_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1671_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *)
  wire _1672_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *)
  wire _1673_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *)
  wire _1674_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *)
  wire _1675_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *)
  wire _1676_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *)
  wire _1677_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *)
  wire _1678_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *)
  wire _1679_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *)
  wire _1680_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *)
  wire _1681_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *)
  wire _1682_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *)
  wire _1683_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *)
  wire _1684_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *)
  wire _1685_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1686_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *)
  wire _1687_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *)
  wire _1688_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *)
  wire _1689_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *)
  wire _1690_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1691_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1692_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1693_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1694_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1695_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1696_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1697_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1698_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1699_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1700_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1701_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1702_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1703_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1704_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1705_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *)
  wire _1706_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2244" *)
  wire _1707_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2245" *)
  wire _1708_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2246" *)
  wire _1709_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2247" *)
  wire _1710_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2248" *)
  wire _1711_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2403" *)
  wire _1712_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2403" *)
  wire _1713_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2499" *)
  wire _1714_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2499" *)
  wire _1715_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2595" *)
  wire _1716_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2595" *)
  wire _1717_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2691" *)
  wire _1718_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2691" *)
  wire _1719_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2787" *)
  wire _1720_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2787" *)
  wire _1721_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1722_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *)
  wire _1723_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2401" *)
  wire _1724_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2497" *)
  wire _1725_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2593" *)
  wire _1726_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2689" *)
  wire _1727_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2785" *)
  wire _1728_;
  wire [2:0] _1729_;
  wire [2:0] _1730_;
  wire [2:0] _1731_;
  wire [2:0] _1732_;
  wire [2:0] _1733_;
  wire [2:0] _1734_;
  wire [2:0] _1735_;
  wire [2:0] _1736_;
  wire [2:0] _1737_;
  wire [2:0] _1738_;
  wire [7:0] _1739_;
  wire [7:0] _1740_;
  wire [7:0] _1741_;
  wire [7:0] _1742_;
  wire [7:0] _1743_;
  wire _1744_;
  wire _1745_;
  wire _1746_;
  wire _1747_;
  wire _1748_;
  wire _1749_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2052" *)
  wire [8:0] _1750_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2055" *)
  wire [8:0] _1751_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2058" *)
  wire [8:0] _1752_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2061" *)
  wire [8:0] _1753_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2064" *)
  wire [8:0] _1754_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:93" *)
  wire [8:0] _1755_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2051" *)
  wire [8:0] _1756_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2052" *)
  wire [8:0] _1757_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2054" *)
  wire [8:0] _1758_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2055" *)
  wire [8:0] _1759_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2057" *)
  wire [8:0] _1760_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2058" *)
  wire [8:0] _1761_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2060" *)
  wire [8:0] _1762_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2061" *)
  wire [8:0] _1763_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2063" *)
  wire [8:0] _1764_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2064" *)
  wire [8:0] _1765_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2268" *)
  wire [7:0] _1766_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2269" *)
  wire [7:0] _1767_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2270" *)
  wire [7:0] _1768_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2271" *)
  wire [7:0] _1769_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2272" *)
  wire [7:0] _1770_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2338" *)
  wire [2:0] _1771_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2350" *)
  wire [2:0] _1772_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2403" *)
  wire _1773_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2434" *)
  wire [2:0] _1774_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2446" *)
  wire [2:0] _1775_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2499" *)
  wire _1776_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2530" *)
  wire [2:0] _1777_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2542" *)
  wire [2:0] _1778_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2595" *)
  wire _1779_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2626" *)
  wire [2:0] _1780_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2638" *)
  wire [2:0] _1781_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2691" *)
  wire _1782_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2722" *)
  wire [2:0] _1783_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2734" *)
  wire [2:0] _1784_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2787" *)
  wire _1785_;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2037" *)
  wire [7:0] adr_ram_rd_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2038" *)
  wire [7:0] adr_ram_rd_data;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2039" *)
  wire adr_ram_rd_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2034" *)
  wire [7:0] adr_ram_wr_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2035" *)
  wire [7:0] adr_ram_wr_data;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2036" *)
  wire adr_ram_wr_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2385" *)
  reg [8:0] cq_rd0_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2386" *)
  reg cq_rd0_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2389" *)
  wire [8:0] cq_rd0_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2387" *)
  wire [8:0] cq_rd0_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2388" *)
  wire [8:0] cq_rd0_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:50" *)
  output [2:0] cq_rd0_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:48" *)
  input cq_rd0_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2326" *)
  reg cq_rd0_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:49" *)
  output cq_rd0_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2481" *)
  reg [8:0] cq_rd1_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2482" *)
  reg cq_rd1_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2485" *)
  wire [8:0] cq_rd1_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2483" *)
  wire [8:0] cq_rd1_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2484" *)
  wire [8:0] cq_rd1_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:53" *)
  output [2:0] cq_rd1_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:51" *)
  input cq_rd1_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2422" *)
  reg cq_rd1_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:52" *)
  output cq_rd1_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2577" *)
  reg [8:0] cq_rd2_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2578" *)
  reg cq_rd2_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2581" *)
  wire [8:0] cq_rd2_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2579" *)
  wire [8:0] cq_rd2_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2580" *)
  wire [8:0] cq_rd2_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:56" *)
  output [2:0] cq_rd2_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:54" *)
  input cq_rd2_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2518" *)
  reg cq_rd2_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:55" *)
  output cq_rd2_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2673" *)
  reg [8:0] cq_rd3_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2674" *)
  reg cq_rd3_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2677" *)
  wire [8:0] cq_rd3_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2675" *)
  wire [8:0] cq_rd3_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2676" *)
  wire [8:0] cq_rd3_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:59" *)
  output [2:0] cq_rd3_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:57" *)
  input cq_rd3_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2614" *)
  reg cq_rd3_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:58" *)
  output cq_rd3_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2769" *)
  reg [8:0] cq_rd4_credits;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2770" *)
  reg cq_rd4_credits_ne0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2773" *)
  wire [8:0] cq_rd4_credits_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2771" *)
  wire [8:0] cq_rd4_credits_w_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2772" *)
  wire [8:0] cq_rd4_credits_wo_take_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:62" *)
  output [2:0] cq_rd4_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:60" *)
  input cq_rd4_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2710" *)
  reg cq_rd4_prdy_d;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:61" *)
  output cq_rd4_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:147" *)
  wire [7:0] cq_rd_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:148" *)
  wire [7:0] cq_rd_adr_p;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2040" *)
  reg [8:0] cq_rd_count0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2042" *)
  reg [8:0] cq_rd_count1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2044" *)
  reg [8:0] cq_rd_count2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2046" *)
  reg [8:0] cq_rd_count3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2048" *)
  reg [8:0] cq_rd_count4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1977" *)
  reg [4:0] cq_rd_credit;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:66" *)
  wire [2:0] cq_rd_pd_p;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:65" *)
  wire cq_rd_take;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2317" *)
  wire [4:0] cq_rd_take_elig;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:67" *)
  wire [2:0] cq_rd_take_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2801" *)
  wire [4:0] cq_rd_take_thread_id_is_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2807" *)
  wire [4:0] cq_rd_take_thread_id_is_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2813" *)
  wire [4:0] cq_rd_take_thread_id_is_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2819" *)
  wire [4:0] cq_rd_take_thread_id_is_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2800" *)
  reg [2:0] cq_rd_take_thread_id_last;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:146" *)
  wire [7:0] cq_wr_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:87" *)
  reg cq_wr_busy_int;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:110" *)
  wire cq_wr_busy_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:91" *)
  reg [8:0] cq_wr_count;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:47" *)
  input [2:0] cq_wr_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:41" *)
  output cq_wr_prdy;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:42" *)
  input cq_wr_pvld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:43" *)
  input [2:0] cq_wr_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1469" *)
  wire flag_l0_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1470" *)
  wire flag_l0_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1479" *)
  wire flag_l0_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1569" *)
  wire flag_l0_100;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1570" *)
  wire flag_l0_101;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1571" *)
  wire flag_l0_102;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1572" *)
  wire flag_l0_103;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1573" *)
  wire flag_l0_104;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1574" *)
  wire flag_l0_105;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1575" *)
  wire flag_l0_106;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1576" *)
  wire flag_l0_107;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1577" *)
  wire flag_l0_108;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1578" *)
  wire flag_l0_109;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1480" *)
  wire flag_l0_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1579" *)
  wire flag_l0_110;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1580" *)
  wire flag_l0_111;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1581" *)
  wire flag_l0_112;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1582" *)
  wire flag_l0_113;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1583" *)
  wire flag_l0_114;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1584" *)
  wire flag_l0_115;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1585" *)
  wire flag_l0_116;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1586" *)
  wire flag_l0_117;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1587" *)
  wire flag_l0_118;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1588" *)
  wire flag_l0_119;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1481" *)
  wire flag_l0_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1589" *)
  wire flag_l0_120;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1590" *)
  wire flag_l0_121;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1591" *)
  wire flag_l0_122;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1592" *)
  wire flag_l0_123;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1593" *)
  wire flag_l0_124;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1594" *)
  wire flag_l0_125;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1595" *)
  wire flag_l0_126;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1482" *)
  wire flag_l0_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1483" *)
  wire flag_l0_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1484" *)
  wire flag_l0_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1485" *)
  wire flag_l0_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1486" *)
  wire flag_l0_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1487" *)
  wire flag_l0_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1488" *)
  wire flag_l0_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1471" *)
  wire flag_l0_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1489" *)
  wire flag_l0_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1490" *)
  wire flag_l0_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1491" *)
  wire flag_l0_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1492" *)
  wire flag_l0_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1493" *)
  wire flag_l0_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1494" *)
  wire flag_l0_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1495" *)
  wire flag_l0_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1496" *)
  wire flag_l0_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1497" *)
  wire flag_l0_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1498" *)
  wire flag_l0_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1472" *)
  wire flag_l0_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1499" *)
  wire flag_l0_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1500" *)
  wire flag_l0_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1501" *)
  wire flag_l0_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1502" *)
  wire flag_l0_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1503" *)
  wire flag_l0_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1504" *)
  wire flag_l0_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1505" *)
  wire flag_l0_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1506" *)
  wire flag_l0_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1507" *)
  wire flag_l0_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1508" *)
  wire flag_l0_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1473" *)
  wire flag_l0_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1509" *)
  wire flag_l0_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1510" *)
  wire flag_l0_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1511" *)
  wire flag_l0_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1512" *)
  wire flag_l0_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1513" *)
  wire flag_l0_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1514" *)
  wire flag_l0_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1515" *)
  wire flag_l0_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1516" *)
  wire flag_l0_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1517" *)
  wire flag_l0_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1518" *)
  wire flag_l0_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1474" *)
  wire flag_l0_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1519" *)
  wire flag_l0_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1520" *)
  wire flag_l0_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1521" *)
  wire flag_l0_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1522" *)
  wire flag_l0_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1523" *)
  wire flag_l0_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1524" *)
  wire flag_l0_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1525" *)
  wire flag_l0_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1526" *)
  wire flag_l0_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1527" *)
  wire flag_l0_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1528" *)
  wire flag_l0_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1475" *)
  wire flag_l0_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1529" *)
  wire flag_l0_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1530" *)
  wire flag_l0_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1531" *)
  wire flag_l0_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1532" *)
  wire flag_l0_63;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1533" *)
  wire flag_l0_64;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1534" *)
  wire flag_l0_65;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1535" *)
  wire flag_l0_66;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1536" *)
  wire flag_l0_67;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1537" *)
  wire flag_l0_68;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1538" *)
  wire flag_l0_69;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1476" *)
  wire flag_l0_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1539" *)
  wire flag_l0_70;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1540" *)
  wire flag_l0_71;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1541" *)
  wire flag_l0_72;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1542" *)
  wire flag_l0_73;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1543" *)
  wire flag_l0_74;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1544" *)
  wire flag_l0_75;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1545" *)
  wire flag_l0_76;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1546" *)
  wire flag_l0_77;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1547" *)
  wire flag_l0_78;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1548" *)
  wire flag_l0_79;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1477" *)
  wire flag_l0_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1549" *)
  wire flag_l0_80;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1550" *)
  wire flag_l0_81;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1551" *)
  wire flag_l0_82;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1552" *)
  wire flag_l0_83;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1553" *)
  wire flag_l0_84;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1554" *)
  wire flag_l0_85;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1555" *)
  wire flag_l0_86;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1556" *)
  wire flag_l0_87;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1557" *)
  wire flag_l0_88;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1558" *)
  wire flag_l0_89;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1478" *)
  wire flag_l0_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1559" *)
  wire flag_l0_90;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1560" *)
  wire flag_l0_91;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1561" *)
  wire flag_l0_92;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1562" *)
  wire flag_l0_93;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1563" *)
  wire flag_l0_94;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1564" *)
  wire flag_l0_95;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1565" *)
  wire flag_l0_96;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1566" *)
  wire flag_l0_97;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1567" *)
  wire flag_l0_98;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1568" *)
  wire flag_l0_99;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1596" *)
  wire flag_l1_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1597" *)
  wire flag_l1_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1606" *)
  wire flag_l1_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1607" *)
  wire flag_l1_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1608" *)
  wire flag_l1_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1609" *)
  wire flag_l1_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1610" *)
  wire flag_l1_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1611" *)
  wire flag_l1_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1612" *)
  wire flag_l1_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1613" *)
  wire flag_l1_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1614" *)
  wire flag_l1_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1615" *)
  wire flag_l1_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1598" *)
  wire flag_l1_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1616" *)
  wire flag_l1_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1617" *)
  wire flag_l1_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1618" *)
  wire flag_l1_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1619" *)
  wire flag_l1_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1620" *)
  wire flag_l1_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1621" *)
  wire flag_l1_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1622" *)
  wire flag_l1_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1623" *)
  wire flag_l1_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1624" *)
  wire flag_l1_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1625" *)
  wire flag_l1_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1599" *)
  wire flag_l1_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1626" *)
  wire flag_l1_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1627" *)
  wire flag_l1_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1628" *)
  wire flag_l1_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1629" *)
  wire flag_l1_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1630" *)
  wire flag_l1_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1631" *)
  wire flag_l1_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1632" *)
  wire flag_l1_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1633" *)
  wire flag_l1_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1634" *)
  wire flag_l1_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1635" *)
  wire flag_l1_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1600" *)
  wire flag_l1_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1636" *)
  wire flag_l1_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1637" *)
  wire flag_l1_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1638" *)
  wire flag_l1_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1639" *)
  wire flag_l1_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1640" *)
  wire flag_l1_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1641" *)
  wire flag_l1_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1642" *)
  wire flag_l1_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1643" *)
  wire flag_l1_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1644" *)
  wire flag_l1_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1645" *)
  wire flag_l1_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1601" *)
  wire flag_l1_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1646" *)
  wire flag_l1_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1647" *)
  wire flag_l1_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1648" *)
  wire flag_l1_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1649" *)
  wire flag_l1_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1650" *)
  wire flag_l1_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1651" *)
  wire flag_l1_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1652" *)
  wire flag_l1_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1653" *)
  wire flag_l1_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1654" *)
  wire flag_l1_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1655" *)
  wire flag_l1_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1602" *)
  wire flag_l1_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1656" *)
  wire flag_l1_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1657" *)
  wire flag_l1_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1658" *)
  wire flag_l1_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1603" *)
  wire flag_l1_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1604" *)
  wire flag_l1_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1605" *)
  wire flag_l1_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1659" *)
  wire flag_l2_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1660" *)
  wire flag_l2_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1669" *)
  wire flag_l2_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1670" *)
  wire flag_l2_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1671" *)
  wire flag_l2_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1672" *)
  wire flag_l2_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1673" *)
  wire flag_l2_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1674" *)
  wire flag_l2_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1675" *)
  wire flag_l2_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1676" *)
  wire flag_l2_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1677" *)
  wire flag_l2_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1678" *)
  wire flag_l2_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1661" *)
  wire flag_l2_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1679" *)
  wire flag_l2_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1680" *)
  wire flag_l2_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1681" *)
  wire flag_l2_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1682" *)
  wire flag_l2_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1683" *)
  wire flag_l2_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1684" *)
  wire flag_l2_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1685" *)
  wire flag_l2_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1686" *)
  wire flag_l2_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1687" *)
  wire flag_l2_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1688" *)
  wire flag_l2_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1662" *)
  wire flag_l2_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1689" *)
  wire flag_l2_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1663" *)
  wire flag_l2_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1664" *)
  wire flag_l2_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1665" *)
  wire flag_l2_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1666" *)
  wire flag_l2_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1667" *)
  wire flag_l2_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1668" *)
  wire flag_l2_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1690" *)
  wire flag_l3_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1691" *)
  wire flag_l3_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1700" *)
  wire flag_l3_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1701" *)
  wire flag_l3_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1702" *)
  wire flag_l3_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1703" *)
  wire flag_l3_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1704" *)
  wire flag_l3_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1692" *)
  wire flag_l3_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1693" *)
  wire flag_l3_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1694" *)
  wire flag_l3_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1695" *)
  wire flag_l3_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1696" *)
  wire flag_l3_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1697" *)
  wire flag_l3_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1698" *)
  wire flag_l3_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1699" *)
  wire flag_l3_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1705" *)
  wire flag_l4_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1706" *)
  wire flag_l4_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1707" *)
  wire flag_l4_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1708" *)
  wire flag_l4_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1709" *)
  wire flag_l4_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1710" *)
  wire flag_l4_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1711" *)
  wire flag_l4_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1712" *)
  wire flag_l5_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1713" *)
  wire flag_l5_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1714" *)
  wire flag_l5_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1715" *)
  wire flag_l6_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:172" *)
  wire [7:0] free_adr_index;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:174" *)
  reg [254:0] free_adr_mask;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:173" *)
  wire [254:0] free_adr_mask_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2004" *)
  reg [7:0] head0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2006" *)
  reg [7:0] head1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2008" *)
  reg [7:0] head2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2010" *)
  reg [7:0] head3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2012" *)
  reg [7:0] head4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1716" *)
  wire index_l0_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1717" *)
  wire index_l0_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1726" *)
  wire index_l0_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1816" *)
  wire index_l0_100;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1817" *)
  wire index_l0_101;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1818" *)
  wire index_l0_102;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1819" *)
  wire index_l0_103;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1820" *)
  wire index_l0_104;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1821" *)
  wire index_l0_105;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1822" *)
  wire index_l0_106;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1823" *)
  wire index_l0_107;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1824" *)
  wire index_l0_108;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1825" *)
  wire index_l0_109;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1727" *)
  wire index_l0_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1826" *)
  wire index_l0_110;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1827" *)
  wire index_l0_111;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1828" *)
  wire index_l0_112;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1829" *)
  wire index_l0_113;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1830" *)
  wire index_l0_114;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1831" *)
  wire index_l0_115;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1832" *)
  wire index_l0_116;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1833" *)
  wire index_l0_117;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1834" *)
  wire index_l0_118;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1835" *)
  wire index_l0_119;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1728" *)
  wire index_l0_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1836" *)
  wire index_l0_120;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1837" *)
  wire index_l0_121;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1838" *)
  wire index_l0_122;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1839" *)
  wire index_l0_123;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1840" *)
  wire index_l0_124;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1841" *)
  wire index_l0_125;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1842" *)
  wire index_l0_126;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1843" *)
  wire index_l0_127;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1729" *)
  wire index_l0_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1730" *)
  wire index_l0_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1731" *)
  wire index_l0_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1732" *)
  wire index_l0_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1733" *)
  wire index_l0_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1734" *)
  wire index_l0_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1735" *)
  wire index_l0_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1718" *)
  wire index_l0_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1736" *)
  wire index_l0_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1737" *)
  wire index_l0_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1738" *)
  wire index_l0_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1739" *)
  wire index_l0_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1740" *)
  wire index_l0_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1741" *)
  wire index_l0_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1742" *)
  wire index_l0_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1743" *)
  wire index_l0_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1744" *)
  wire index_l0_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1745" *)
  wire index_l0_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1719" *)
  wire index_l0_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1746" *)
  wire index_l0_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1747" *)
  wire index_l0_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1748" *)
  wire index_l0_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1749" *)
  wire index_l0_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1750" *)
  wire index_l0_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1751" *)
  wire index_l0_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1752" *)
  wire index_l0_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1753" *)
  wire index_l0_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1754" *)
  wire index_l0_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1755" *)
  wire index_l0_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1720" *)
  wire index_l0_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1756" *)
  wire index_l0_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1757" *)
  wire index_l0_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1758" *)
  wire index_l0_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1759" *)
  wire index_l0_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1760" *)
  wire index_l0_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1761" *)
  wire index_l0_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1762" *)
  wire index_l0_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1763" *)
  wire index_l0_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1764" *)
  wire index_l0_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1765" *)
  wire index_l0_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1721" *)
  wire index_l0_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1766" *)
  wire index_l0_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1767" *)
  wire index_l0_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1768" *)
  wire index_l0_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1769" *)
  wire index_l0_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1770" *)
  wire index_l0_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1771" *)
  wire index_l0_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1772" *)
  wire index_l0_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1773" *)
  wire index_l0_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1774" *)
  wire index_l0_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1775" *)
  wire index_l0_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1722" *)
  wire index_l0_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1776" *)
  wire index_l0_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1777" *)
  wire index_l0_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1778" *)
  wire index_l0_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1779" *)
  wire index_l0_63;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1780" *)
  wire index_l0_64;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1781" *)
  wire index_l0_65;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1782" *)
  wire index_l0_66;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1783" *)
  wire index_l0_67;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1784" *)
  wire index_l0_68;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1785" *)
  wire index_l0_69;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1723" *)
  wire index_l0_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1786" *)
  wire index_l0_70;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1787" *)
  wire index_l0_71;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1788" *)
  wire index_l0_72;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1789" *)
  wire index_l0_73;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1790" *)
  wire index_l0_74;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1791" *)
  wire index_l0_75;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1792" *)
  wire index_l0_76;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1793" *)
  wire index_l0_77;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1794" *)
  wire index_l0_78;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1795" *)
  wire index_l0_79;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1724" *)
  wire index_l0_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1796" *)
  wire index_l0_80;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1797" *)
  wire index_l0_81;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1798" *)
  wire index_l0_82;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1799" *)
  wire index_l0_83;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1800" *)
  wire index_l0_84;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1801" *)
  wire index_l0_85;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1802" *)
  wire index_l0_86;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1803" *)
  wire index_l0_87;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1804" *)
  wire index_l0_88;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1805" *)
  wire index_l0_89;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1725" *)
  wire index_l0_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1806" *)
  wire index_l0_90;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1807" *)
  wire index_l0_91;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1808" *)
  wire index_l0_92;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1809" *)
  wire index_l0_93;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1810" *)
  wire index_l0_94;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1811" *)
  wire index_l0_95;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1812" *)
  wire index_l0_96;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1813" *)
  wire index_l0_97;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1814" *)
  wire index_l0_98;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1815" *)
  wire index_l0_99;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1844" *)
  wire [1:0] index_l1_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1845" *)
  wire [1:0] index_l1_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1854" *)
  wire [1:0] index_l1_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1855" *)
  wire [1:0] index_l1_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1856" *)
  wire [1:0] index_l1_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1857" *)
  wire [1:0] index_l1_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1858" *)
  wire [1:0] index_l1_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1859" *)
  wire [1:0] index_l1_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1860" *)
  wire [1:0] index_l1_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1861" *)
  wire [1:0] index_l1_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1862" *)
  wire [1:0] index_l1_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1863" *)
  wire [1:0] index_l1_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1846" *)
  wire [1:0] index_l1_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1864" *)
  wire [1:0] index_l1_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1865" *)
  wire [1:0] index_l1_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1866" *)
  wire [1:0] index_l1_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1867" *)
  wire [1:0] index_l1_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1868" *)
  wire [1:0] index_l1_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1869" *)
  wire [1:0] index_l1_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1870" *)
  wire [1:0] index_l1_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1871" *)
  wire [1:0] index_l1_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1872" *)
  wire [1:0] index_l1_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1873" *)
  wire [1:0] index_l1_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1847" *)
  wire [1:0] index_l1_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1874" *)
  wire [1:0] index_l1_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1875" *)
  wire [1:0] index_l1_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1876" *)
  wire [1:0] index_l1_32;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1877" *)
  wire [1:0] index_l1_33;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1878" *)
  wire [1:0] index_l1_34;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1879" *)
  wire [1:0] index_l1_35;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1880" *)
  wire [1:0] index_l1_36;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1881" *)
  wire [1:0] index_l1_37;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1882" *)
  wire [1:0] index_l1_38;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1883" *)
  wire [1:0] index_l1_39;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1848" *)
  wire [1:0] index_l1_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1884" *)
  wire [1:0] index_l1_40;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1885" *)
  wire [1:0] index_l1_41;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1886" *)
  wire [1:0] index_l1_42;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1887" *)
  wire [1:0] index_l1_43;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1888" *)
  wire [1:0] index_l1_44;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1889" *)
  wire [1:0] index_l1_45;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1890" *)
  wire [1:0] index_l1_46;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1891" *)
  wire [1:0] index_l1_47;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1892" *)
  wire [1:0] index_l1_48;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1893" *)
  wire [1:0] index_l1_49;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1849" *)
  wire [1:0] index_l1_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1894" *)
  wire [1:0] index_l1_50;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1895" *)
  wire [1:0] index_l1_51;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1896" *)
  wire [1:0] index_l1_52;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1897" *)
  wire [1:0] index_l1_53;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1898" *)
  wire [1:0] index_l1_54;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1899" *)
  wire [1:0] index_l1_55;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1900" *)
  wire [1:0] index_l1_56;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1901" *)
  wire [1:0] index_l1_57;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1902" *)
  wire [1:0] index_l1_58;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1903" *)
  wire [1:0] index_l1_59;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1850" *)
  wire [1:0] index_l1_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1904" *)
  wire [1:0] index_l1_60;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1905" *)
  wire [1:0] index_l1_61;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1906" *)
  wire [1:0] index_l1_62;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1907" *)
  wire [1:0] index_l1_63;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1851" *)
  wire [1:0] index_l1_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1852" *)
  wire [1:0] index_l1_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1853" *)
  wire [1:0] index_l1_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1908" *)
  wire [2:0] index_l2_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1909" *)
  wire [2:0] index_l2_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1918" *)
  wire [2:0] index_l2_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1919" *)
  wire [2:0] index_l2_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1920" *)
  wire [2:0] index_l2_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1921" *)
  wire [2:0] index_l2_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1922" *)
  wire [2:0] index_l2_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1923" *)
  wire [2:0] index_l2_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1924" *)
  wire [2:0] index_l2_16;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1925" *)
  wire [2:0] index_l2_17;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1926" *)
  wire [2:0] index_l2_18;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1927" *)
  wire [2:0] index_l2_19;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1910" *)
  wire [2:0] index_l2_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1928" *)
  wire [2:0] index_l2_20;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1929" *)
  wire [2:0] index_l2_21;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1930" *)
  wire [2:0] index_l2_22;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1931" *)
  wire [2:0] index_l2_23;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1932" *)
  wire [2:0] index_l2_24;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1933" *)
  wire [2:0] index_l2_25;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1934" *)
  wire [2:0] index_l2_26;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1935" *)
  wire [2:0] index_l2_27;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1936" *)
  wire [2:0] index_l2_28;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1937" *)
  wire [2:0] index_l2_29;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1911" *)
  wire [2:0] index_l2_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1938" *)
  wire [2:0] index_l2_30;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1939" *)
  wire [2:0] index_l2_31;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1912" *)
  wire [2:0] index_l2_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1913" *)
  wire [2:0] index_l2_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1914" *)
  wire [2:0] index_l2_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1915" *)
  wire [2:0] index_l2_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1916" *)
  wire [2:0] index_l2_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1917" *)
  wire [2:0] index_l2_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1940" *)
  wire [3:0] index_l3_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1941" *)
  wire [3:0] index_l3_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1950" *)
  wire [3:0] index_l3_10;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1951" *)
  wire [3:0] index_l3_11;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1952" *)
  wire [3:0] index_l3_12;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1953" *)
  wire [3:0] index_l3_13;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1954" *)
  wire [3:0] index_l3_14;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1955" *)
  wire [3:0] index_l3_15;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1942" *)
  wire [3:0] index_l3_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1943" *)
  wire [3:0] index_l3_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1944" *)
  wire [3:0] index_l3_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1945" *)
  wire [3:0] index_l3_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1946" *)
  wire [3:0] index_l3_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1947" *)
  wire [3:0] index_l3_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1948" *)
  wire [3:0] index_l3_8;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1949" *)
  wire [3:0] index_l3_9;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1956" *)
  wire [4:0] index_l4_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1957" *)
  wire [4:0] index_l4_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1958" *)
  wire [4:0] index_l4_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1959" *)
  wire [4:0] index_l4_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1960" *)
  wire [4:0] index_l4_4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1961" *)
  wire [4:0] index_l4_5;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1962" *)
  wire [4:0] index_l4_6;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1963" *)
  wire [4:0] index_l4_7;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1964" *)
  wire [5:0] index_l5_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1965" *)
  wire [5:0] index_l5_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1966" *)
  wire [5:0] index_l5_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1967" *)
  wire [5:0] index_l5_3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1968" *)
  wire [6:0] index_l6_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1969" *)
  wire [6:0] index_l6_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1970" *)
  wire [7:0] index_l7_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:39" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:75" *)
  wire nvdla_core_clk_mgated;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:74" *)
  wire nvdla_core_clk_mgated_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:71" *)
  wire nvdla_core_clk_mgated_skid;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:72" *)
  wire nvdla_core_clk_mgated_skid_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:40" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:63" *)
  input [31:0] pwrbus_ram_pd;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2294" *)
  reg [7:0] rd_adr_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2319" *)
  wire rd_bypassing0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2415" *)
  wire rd_bypassing1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2511" *)
  wire rd_bypassing2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2607" *)
  wire rd_bypassing3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2703" *)
  wire rd_bypassing4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2041" *)
  wire [8:0] rd_count0_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2043" *)
  wire [8:0] rd_count1_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2045" *)
  wire [8:0] rd_count2_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2047" *)
  wire [8:0] rd_count3_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2049" *)
  wire [8:0] rd_count4_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:149" *)
  wire rd_enable;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:161" *)
  wire rd_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:171" *)
  wire [7:0] rd_popping_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2318" *)
  wire rd_pre_bypassing0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2414" *)
  wire rd_pre_bypassing1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2510" *)
  wire rd_pre_bypassing2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2606" *)
  wire rd_pre_bypassing3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2702" *)
  wire rd_pre_bypassing4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:164" *)
  wire rd_pushing;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1994" *)
  wire rd_pushing0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1995" *)
  wire rd_pushing1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1996" *)
  wire rd_pushing2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1997" *)
  wire rd_pushing3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1998" *)
  wire rd_pushing4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:166" *)
  wire [7:0] rd_pushing_adr;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1978" *)
  reg rd_pushing_q;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:165" *)
  wire [2:0] rd_pushing_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2320" *)
  reg [2:0] rd_skid0_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2323" *)
  reg rd_skid0_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2321" *)
  reg [2:0] rd_skid0_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2324" *)
  reg rd_skid0_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2322" *)
  reg [2:0] rd_skid0_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2325" *)
  reg rd_skid0_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2416" *)
  reg [2:0] rd_skid1_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2419" *)
  reg rd_skid1_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2417" *)
  reg [2:0] rd_skid1_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2420" *)
  reg rd_skid1_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2418" *)
  reg [2:0] rd_skid1_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2421" *)
  reg rd_skid1_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2512" *)
  reg [2:0] rd_skid2_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2515" *)
  reg rd_skid2_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2513" *)
  reg [2:0] rd_skid2_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2516" *)
  reg rd_skid2_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2514" *)
  reg [2:0] rd_skid2_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2517" *)
  reg rd_skid2_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2608" *)
  reg [2:0] rd_skid3_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2611" *)
  reg rd_skid3_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2609" *)
  reg [2:0] rd_skid3_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2612" *)
  reg rd_skid3_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2610" *)
  reg [2:0] rd_skid3_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2613" *)
  reg rd_skid3_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2704" *)
  reg [2:0] rd_skid4_0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2707" *)
  reg rd_skid4_0_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2705" *)
  reg [2:0] rd_skid4_1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2708" *)
  reg rd_skid4_1_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2706" *)
  reg [2:0] rd_skid4_2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2709" *)
  reg rd_skid4_2_vld;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1999" *)
  wire rd_take0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2000" *)
  wire rd_take1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2001" *)
  wire rd_take2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2002" *)
  wire rd_take3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2003" *)
  wire rd_take4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2292" *)
  reg rd_take_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2015" *)
  wire rd_take_dly_cg;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2014" *)
  reg [4:0] rd_take_n_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2005" *)
  reg [7:0] tail0;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2007" *)
  reg [7:0] tail1;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2009" *)
  reg [7:0] tail2;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2011" *)
  reg [7:0] tail3;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2013" *)
  reg [7:0] tail4;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2120" *)
  reg [4:0] update_head;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2121" *)
  wire [4:0] update_head_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2016" *)
  wire update_rd_take_n_dly;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:145" *)
  wire wr_adr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:69" *)
  wire wr_bypassing;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:95" *)
  wire [8:0] wr_count_next;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:98" *)
  wire wr_count_next_is_256;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:94" *)
  wire [8:0] wr_count_next_no_wr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:97" *)
  wire wr_count_next_no_wr_popping_is_256;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:93" *)
  wire [8:0] wr_count_next_wr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:100" *)
  wire [8:0] wr_limit_muxed;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:101" *)
  wire [8:0] wr_limit_reg;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:90" *)
  wire wr_popping;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:140" *)
  wire wr_pushing;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:141" *)
  wire [2:0] wr_pushing_thread_id;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:86" *)
  wire wr_reserving;
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:92" *)
  wire wr_reserving_and_not_bypassing;
  assign _0318_ = cq_rd_count0 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2051" *) 1'b1;
  assign _0319_ = cq_rd_count1 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2054" *) 1'b1;
  assign _0320_ = cq_rd_count2 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2057" *) 1'b1;
  assign _0321_ = cq_rd_count3 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2060" *) 1'b1;
  assign _0322_ = cq_rd_count4 + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2063" *) 1'b1;
  assign cq_rd0_credits_wo_take_next = cq_rd0_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2387" *) cq_rd_credit[0];
  assign cq_rd1_credits_wo_take_next = cq_rd1_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2483" *) cq_rd_credit[1];
  assign cq_rd2_credits_wo_take_next = cq_rd2_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2579" *) cq_rd_credit[2];
  assign cq_rd3_credits_wo_take_next = cq_rd3_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2675" *) cq_rd_credit[3];
  assign cq_rd4_credits_wo_take_next = cq_rd4_credits + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2771" *) cq_rd_credit[4];
  assign _0323_ = cq_wr_count + (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:94" *) 1'b1;
  assign _0324_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1000" *) 8'b10100001;
  assign _0325_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1003" *) 8'b10100010;
  assign _0326_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1005" *) 8'b10100010;
  assign _0327_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1008" *) 8'b10100011;
  assign _0328_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1010" *) 8'b10100011;
  assign _0329_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1013" *) 8'b10100100;
  assign _0330_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1015" *) 8'b10100100;
  assign _0331_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1018" *) 8'b10100101;
  assign _0332_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1020" *) 8'b10100101;
  assign _0333_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1023" *) 8'b10100110;
  assign _0334_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1025" *) 8'b10100110;
  assign _0335_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1028" *) 8'b10100111;
  assign _0336_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1030" *) 8'b10100111;
  assign _0337_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1033" *) 8'b10101000;
  assign _0338_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1035" *) 8'b10101000;
  assign _0339_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1038" *) 8'b10101001;
  assign _0340_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1040" *) 8'b10101001;
  assign _0341_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1043" *) 8'b10101010;
  assign _0342_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1045" *) 8'b10101010;
  assign _0343_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1048" *) 8'b10101011;
  assign _0344_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1050" *) 8'b10101011;
  assign _0345_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1053" *) 8'b10101100;
  assign _0346_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1055" *) 8'b10101100;
  assign _0347_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1058" *) 8'b10101101;
  assign _0348_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1060" *) 8'b10101101;
  assign _0349_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1063" *) 8'b10101110;
  assign _0350_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1065" *) 8'b10101110;
  assign _0351_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1068" *) 8'b10101111;
  assign _0352_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1070" *) 8'b10101111;
  assign _0353_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1073" *) 8'b10110000;
  assign _0354_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1075" *) 8'b10110000;
  assign _0355_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1078" *) 8'b10110001;
  assign _0356_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1080" *) 8'b10110001;
  assign _0357_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1083" *) 8'b10110010;
  assign _0358_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1085" *) 8'b10110010;
  assign _0359_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1088" *) 8'b10110011;
  assign _0360_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1090" *) 8'b10110011;
  assign _0361_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1093" *) 8'b10110100;
  assign _0362_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1095" *) 8'b10110100;
  assign _0363_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1098" *) 8'b10110101;
  assign _0364_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1100" *) 8'b10110101;
  assign _0365_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1103" *) 8'b10110110;
  assign _0366_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1105" *) 8'b10110110;
  assign _0367_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1108" *) 8'b10110111;
  assign _0368_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1110" *) 8'b10110111;
  assign _0369_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1113" *) 8'b10111000;
  assign _0370_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1115" *) 8'b10111000;
  assign _0371_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1118" *) 8'b10111001;
  assign _0372_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1120" *) 8'b10111001;
  assign _0373_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1123" *) 8'b10111010;
  assign _0374_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1125" *) 8'b10111010;
  assign _0375_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1128" *) 8'b10111011;
  assign _0376_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1130" *) 8'b10111011;
  assign _0377_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1133" *) 8'b10111100;
  assign _0378_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1135" *) 8'b10111100;
  assign _0379_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1138" *) 8'b10111101;
  assign _0380_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1140" *) 8'b10111101;
  assign _0381_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1143" *) 8'b10111110;
  assign _0382_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1145" *) 8'b10111110;
  assign _0383_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1148" *) 8'b10111111;
  assign _0384_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1150" *) 8'b10111111;
  assign _0385_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1153" *) 8'b11000000;
  assign _0386_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1155" *) 8'b11000000;
  assign _0387_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1158" *) 8'b11000001;
  assign _0388_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1160" *) 8'b11000001;
  assign _0389_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1163" *) 8'b11000010;
  assign _0390_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1165" *) 8'b11000010;
  assign _0391_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1168" *) 8'b11000011;
  assign _0392_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1170" *) 8'b11000011;
  assign _0393_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1173" *) 8'b11000100;
  assign _0394_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1175" *) 8'b11000100;
  assign _0395_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1178" *) 8'b11000101;
  assign _0396_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1180" *) 8'b11000101;
  assign _0397_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1183" *) 8'b11000110;
  assign _0398_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1185" *) 8'b11000110;
  assign _0399_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1188" *) 8'b11000111;
  assign _0400_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1190" *) 8'b11000111;
  assign _0401_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1193" *) 8'b11001000;
  assign _0402_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1195" *) 8'b11001000;
  assign _0403_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1198" *) 8'b11001001;
  assign _0404_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1200" *) 8'b11001001;
  assign _0405_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1203" *) 8'b11001010;
  assign _0406_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1205" *) 8'b11001010;
  assign _0407_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1208" *) 8'b11001011;
  assign _0408_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1210" *) 8'b11001011;
  assign _0409_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1213" *) 8'b11001100;
  assign _0410_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1215" *) 8'b11001100;
  assign _0411_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1218" *) 8'b11001101;
  assign _0412_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1220" *) 8'b11001101;
  assign _0413_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1223" *) 8'b11001110;
  assign _0414_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1225" *) 8'b11001110;
  assign _0415_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1228" *) 8'b11001111;
  assign _0416_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1230" *) 8'b11001111;
  assign _0417_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1233" *) 8'b11010000;
  assign _0418_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1235" *) 8'b11010000;
  assign _0419_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1238" *) 8'b11010001;
  assign _0420_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1240" *) 8'b11010001;
  assign _0421_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1243" *) 8'b11010010;
  assign _0422_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1245" *) 8'b11010010;
  assign _0423_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1248" *) 8'b11010011;
  assign _0424_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1250" *) 8'b11010011;
  assign _0425_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1253" *) 8'b11010100;
  assign _0426_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1255" *) 8'b11010100;
  assign _0427_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1258" *) 8'b11010101;
  assign _0428_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1260" *) 8'b11010101;
  assign _0429_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1263" *) 8'b11010110;
  assign _0430_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1265" *) 8'b11010110;
  assign _0431_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1268" *) 8'b11010111;
  assign _0432_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1270" *) 8'b11010111;
  assign _0433_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1273" *) 8'b11011000;
  assign _0434_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1275" *) 8'b11011000;
  assign _0435_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1278" *) 8'b11011001;
  assign _0436_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1280" *) 8'b11011001;
  assign _0437_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1283" *) 8'b11011010;
  assign _0438_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1285" *) 8'b11011010;
  assign _0439_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1288" *) 8'b11011011;
  assign _0440_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1290" *) 8'b11011011;
  assign _0441_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1293" *) 8'b11011100;
  assign _0442_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1295" *) 8'b11011100;
  assign _0443_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1298" *) 8'b11011101;
  assign _0444_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1300" *) 8'b11011101;
  assign _0445_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1303" *) 8'b11011110;
  assign _0446_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1305" *) 8'b11011110;
  assign _0447_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1308" *) 8'b11011111;
  assign _0448_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1310" *) 8'b11011111;
  assign _0449_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1313" *) 8'b11100000;
  assign _0450_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1315" *) 8'b11100000;
  assign _0451_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1318" *) 8'b11100001;
  assign _0452_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1320" *) 8'b11100001;
  assign _0453_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1323" *) 8'b11100010;
  assign _0454_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1325" *) 8'b11100010;
  assign _0455_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1328" *) 8'b11100011;
  assign _0456_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1330" *) 8'b11100011;
  assign _0457_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1333" *) 8'b11100100;
  assign _0458_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1335" *) 8'b11100100;
  assign _0459_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1338" *) 8'b11100101;
  assign _0460_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1340" *) 8'b11100101;
  assign _0461_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1343" *) 8'b11100110;
  assign _0462_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1345" *) 8'b11100110;
  assign _0463_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1348" *) 8'b11100111;
  assign _0464_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1350" *) 8'b11100111;
  assign _0465_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1353" *) 8'b11101000;
  assign _0466_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1355" *) 8'b11101000;
  assign _0467_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1358" *) 8'b11101001;
  assign _0468_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1360" *) 8'b11101001;
  assign _0469_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1363" *) 8'b11101010;
  assign _0470_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1365" *) 8'b11101010;
  assign _0471_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1368" *) 8'b11101011;
  assign _0472_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1370" *) 8'b11101011;
  assign _0473_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1373" *) 8'b11101100;
  assign _0474_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1375" *) 8'b11101100;
  assign _0475_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1378" *) 8'b11101101;
  assign _0476_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1380" *) 8'b11101101;
  assign _0477_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1383" *) 8'b11101110;
  assign _0478_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1385" *) 8'b11101110;
  assign _0479_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1388" *) 8'b11101111;
  assign _0480_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1390" *) 8'b11101111;
  assign _0481_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1393" *) 8'b11110000;
  assign _0482_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1395" *) 8'b11110000;
  assign _0483_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1398" *) 8'b11110001;
  assign _0484_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1400" *) 8'b11110001;
  assign _0485_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1403" *) 8'b11110010;
  assign _0486_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1405" *) 8'b11110010;
  assign _0487_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1408" *) 8'b11110011;
  assign _0488_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1410" *) 8'b11110011;
  assign _0489_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1413" *) 8'b11110100;
  assign _0490_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1415" *) 8'b11110100;
  assign _0491_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1418" *) 8'b11110101;
  assign _0492_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1420" *) 8'b11110101;
  assign _0493_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1423" *) 8'b11110110;
  assign _0494_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1425" *) 8'b11110110;
  assign _0495_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1428" *) 8'b11110111;
  assign _0496_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1430" *) 8'b11110111;
  assign _0497_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1433" *) 8'b11111000;
  assign _0498_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1435" *) 8'b11111000;
  assign _0499_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1438" *) 8'b11111001;
  assign _0500_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1440" *) 8'b11111001;
  assign _0501_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1443" *) 8'b11111010;
  assign _0502_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1445" *) 8'b11111010;
  assign _0503_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1448" *) 8'b11111011;
  assign _0504_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1450" *) 8'b11111011;
  assign _0505_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1453" *) 8'b11111100;
  assign _0506_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1455" *) 8'b11111100;
  assign _0507_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1458" *) 8'b11111101;
  assign _0508_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1460" *) 8'b11111101;
  assign _0509_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1463" *) 8'b11111110;
  assign _0510_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1465" *) 8'b11111110;
  assign _0511_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:193" *) rd_adr_dly;
  assign _0512_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:195" *) adr_ram_wr_data;
  assign _0513_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:198" *) 1'b1;
  assign _0514_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1985" *) cq_wr_thread_id;
  assign _0515_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1986" *) 1'b1;
  assign _0516_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1987" *) 2'b10;
  assign _0517_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1988" *) 2'b11;
  assign _0518_ = cq_wr_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1989" *) 3'b100;
  assign _0519_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1999" *) cq_rd_take_thread_id;
  assign _0520_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:200" *) 1'b1;
  assign _0521_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2000" *) 1'b1;
  assign _0522_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2001" *) 2'b10;
  assign _0523_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2002" *) 2'b11;
  assign _0524_ = cq_rd_take_thread_id == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2003" *) 3'b100;
  assign _0525_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:203" *) 2'b10;
  assign _0526_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:205" *) 2'b10;
  assign _0527_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:208" *) 2'b11;
  assign _0528_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:210" *) 2'b11;
  assign _0529_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:213" *) 3'b100;
  assign _0530_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:215" *) 3'b100;
  assign _0531_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2152" *) cq_rd_count0;
  assign _0532_ = cq_rd_count0 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *) 1'b1;
  assign _0533_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2167" *) cq_rd_count1;
  assign _0534_ = cq_rd_count1 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *) 1'b1;
  assign _0535_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:218" *) 3'b101;
  assign _0536_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2182" *) cq_rd_count2;
  assign _0537_ = cq_rd_count2 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *) 1'b1;
  assign _0538_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2197" *) cq_rd_count3;
  assign _0539_ = cq_rd_count3 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *) 1'b1;
  assign _0540_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:220" *) 3'b101;
  assign _0541_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2212" *) cq_rd_count4;
  assign _0542_ = cq_rd_count4 == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *) 1'b1;
  assign _0543_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:223" *) 3'b110;
  assign _0544_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:225" *) 3'b110;
  assign _0545_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:228" *) 3'b111;
  assign _0546_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:230" *) 3'b111;
  assign _0547_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:233" *) 4'b1000;
  assign _0548_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:235" *) 4'b1000;
  assign _0549_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:238" *) 4'b1001;
  assign _0550_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) cq_rd0_credits;
  assign _0551_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:240" *) 4'b1001;
  assign _0552_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:243" *) 4'b1010;
  assign _0553_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:245" *) 4'b1010;
  assign _0554_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:248" *) 4'b1011;
  assign _0555_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) cq_rd1_credits;
  assign _0556_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:250" *) 4'b1011;
  assign _0557_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:253" *) 4'b1100;
  assign _0558_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:255" *) 4'b1100;
  assign _0559_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:258" *) 4'b1101;
  assign _0560_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) cq_rd2_credits;
  assign _0561_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:260" *) 4'b1101;
  assign _0562_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:263" *) 4'b1110;
  assign _0563_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:265" *) 4'b1110;
  assign _0564_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:268" *) 4'b1111;
  assign _0565_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) cq_rd3_credits;
  assign _0566_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:270" *) 4'b1111;
  assign _0567_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:273" *) 5'b10000;
  assign _0568_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:275" *) 5'b10000;
  assign _0569_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) cq_rd4_credits;
  assign _0570_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:278" *) 5'b10001;
  assign _0571_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:280" *) 5'b10001;
  assign _0572_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *) 3'b100;
  assign _0573_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *) 2'b11;
  assign _0574_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *) 2'b10;
  assign _0575_ = cq_rd_take_thread_id_last == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) 1'b1;
  assign _0576_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2806" *) cq_rd_take_thread_id_last;
  assign _0577_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:283" *) 5'b10010;
  assign _0578_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:285" *) 5'b10010;
  assign _0579_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:288" *) 5'b10011;
  assign _0580_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:290" *) 5'b10011;
  assign _0581_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:293" *) 5'b10100;
  assign _0582_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:295" *) 5'b10100;
  assign _0583_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:298" *) 5'b10101;
  assign _0584_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:300" *) 5'b10101;
  assign _0585_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:303" *) 5'b10110;
  assign _0586_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:305" *) 5'b10110;
  assign _0587_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:308" *) 5'b10111;
  assign _0588_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:310" *) 5'b10111;
  assign _0589_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:313" *) 5'b11000;
  assign _0590_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:315" *) 5'b11000;
  assign _0591_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:318" *) 5'b11001;
  assign _0592_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:320" *) 5'b11001;
  assign _0593_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:323" *) 5'b11010;
  assign _0594_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:325" *) 5'b11010;
  assign _0595_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:328" *) 5'b11011;
  assign _0596_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:330" *) 5'b11011;
  assign _0597_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:333" *) 5'b11100;
  assign _0598_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:335" *) 5'b11100;
  assign _0599_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:338" *) 5'b11101;
  assign _0600_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:340" *) 5'b11101;
  assign _0601_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:343" *) 5'b11110;
  assign _0602_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:345" *) 5'b11110;
  assign _0603_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:348" *) 5'b11111;
  assign _0604_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:350" *) 5'b11111;
  assign _0605_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:353" *) 6'b100000;
  assign _0606_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:355" *) 6'b100000;
  assign _0607_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:358" *) 6'b100001;
  assign _0608_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:360" *) 6'b100001;
  assign _0609_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:363" *) 6'b100010;
  assign _0610_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:365" *) 6'b100010;
  assign _0611_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:368" *) 6'b100011;
  assign _0612_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:370" *) 6'b100011;
  assign _0613_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:373" *) 6'b100100;
  assign _0614_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:375" *) 6'b100100;
  assign _0615_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:378" *) 6'b100101;
  assign _0616_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:380" *) 6'b100101;
  assign _0617_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:383" *) 6'b100110;
  assign _0618_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:385" *) 6'b100110;
  assign _0619_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:388" *) 6'b100111;
  assign _0620_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:390" *) 6'b100111;
  assign _0621_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:393" *) 6'b101000;
  assign _0622_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:395" *) 6'b101000;
  assign _0623_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:398" *) 6'b101001;
  assign _0624_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:400" *) 6'b101001;
  assign _0625_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:403" *) 6'b101010;
  assign _0626_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:405" *) 6'b101010;
  assign _0627_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:408" *) 6'b101011;
  assign _0628_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:410" *) 6'b101011;
  assign _0629_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:413" *) 6'b101100;
  assign _0630_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:415" *) 6'b101100;
  assign _0631_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:418" *) 6'b101101;
  assign _0632_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:420" *) 6'b101101;
  assign _0633_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:423" *) 6'b101110;
  assign _0634_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:425" *) 6'b101110;
  assign _0635_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:428" *) 6'b101111;
  assign _0636_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:430" *) 6'b101111;
  assign _0637_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:433" *) 6'b110000;
  assign _0638_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:435" *) 6'b110000;
  assign _0639_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:438" *) 6'b110001;
  assign _0640_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:440" *) 6'b110001;
  assign _0641_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:443" *) 6'b110010;
  assign _0642_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:445" *) 6'b110010;
  assign _0643_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:448" *) 6'b110011;
  assign _0644_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:450" *) 6'b110011;
  assign _0645_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:453" *) 6'b110100;
  assign _0646_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:455" *) 6'b110100;
  assign _0647_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:458" *) 6'b110101;
  assign _0648_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:460" *) 6'b110101;
  assign _0649_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:463" *) 6'b110110;
  assign _0650_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:465" *) 6'b110110;
  assign _0651_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:468" *) 6'b110111;
  assign _0652_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:470" *) 6'b110111;
  assign _0653_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:473" *) 6'b111000;
  assign _0654_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:475" *) 6'b111000;
  assign _0655_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:478" *) 6'b111001;
  assign _0656_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:480" *) 6'b111001;
  assign _0657_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:483" *) 6'b111010;
  assign _0658_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:485" *) 6'b111010;
  assign _0659_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:488" *) 6'b111011;
  assign _0660_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:490" *) 6'b111011;
  assign _0661_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:493" *) 6'b111100;
  assign _0662_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:495" *) 6'b111100;
  assign _0663_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:498" *) 6'b111101;
  assign _0664_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:500" *) 6'b111101;
  assign _0665_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:503" *) 6'b111110;
  assign _0666_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:505" *) 6'b111110;
  assign _0667_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:508" *) 6'b111111;
  assign _0668_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:510" *) 6'b111111;
  assign _0669_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:513" *) 7'b1000000;
  assign _0670_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:515" *) 7'b1000000;
  assign _0671_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:518" *) 7'b1000001;
  assign _0672_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:520" *) 7'b1000001;
  assign _0673_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:523" *) 7'b1000010;
  assign _0674_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:525" *) 7'b1000010;
  assign _0675_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:528" *) 7'b1000011;
  assign _0676_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:530" *) 7'b1000011;
  assign _0677_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:533" *) 7'b1000100;
  assign _0678_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:535" *) 7'b1000100;
  assign _0679_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:538" *) 7'b1000101;
  assign _0680_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:540" *) 7'b1000101;
  assign _0681_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:543" *) 7'b1000110;
  assign _0682_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:545" *) 7'b1000110;
  assign _0683_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:548" *) 7'b1000111;
  assign _0684_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:550" *) 7'b1000111;
  assign _0685_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:553" *) 7'b1001000;
  assign _0686_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:555" *) 7'b1001000;
  assign _0687_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:558" *) 7'b1001001;
  assign _0688_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:560" *) 7'b1001001;
  assign _0689_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:563" *) 7'b1001010;
  assign _0690_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:565" *) 7'b1001010;
  assign _0691_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:568" *) 7'b1001011;
  assign _0692_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:570" *) 7'b1001011;
  assign _0693_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:573" *) 7'b1001100;
  assign _0694_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:575" *) 7'b1001100;
  assign _0695_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:578" *) 7'b1001101;
  assign _0696_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:580" *) 7'b1001101;
  assign _0697_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:583" *) 7'b1001110;
  assign _0698_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:585" *) 7'b1001110;
  assign _0699_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:588" *) 7'b1001111;
  assign _0700_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:590" *) 7'b1001111;
  assign _0701_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:593" *) 7'b1010000;
  assign _0702_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:595" *) 7'b1010000;
  assign _0703_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:598" *) 7'b1010001;
  assign _0704_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:600" *) 7'b1010001;
  assign _0705_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:603" *) 7'b1010010;
  assign _0706_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:605" *) 7'b1010010;
  assign _0707_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:608" *) 7'b1010011;
  assign _0708_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:610" *) 7'b1010011;
  assign _0709_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:613" *) 7'b1010100;
  assign _0710_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:615" *) 7'b1010100;
  assign _0711_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:618" *) 7'b1010101;
  assign _0712_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:620" *) 7'b1010101;
  assign _0713_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:623" *) 7'b1010110;
  assign _0714_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:625" *) 7'b1010110;
  assign _0715_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:628" *) 7'b1010111;
  assign _0716_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:630" *) 7'b1010111;
  assign _0717_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:633" *) 7'b1011000;
  assign _0718_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:635" *) 7'b1011000;
  assign _0719_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:638" *) 7'b1011001;
  assign _0720_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:640" *) 7'b1011001;
  assign _0721_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:643" *) 7'b1011010;
  assign _0722_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:645" *) 7'b1011010;
  assign _0723_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:648" *) 7'b1011011;
  assign _0724_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:650" *) 7'b1011011;
  assign _0725_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:653" *) 7'b1011100;
  assign _0726_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:655" *) 7'b1011100;
  assign _0727_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:658" *) 7'b1011101;
  assign _0728_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:660" *) 7'b1011101;
  assign _0729_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:663" *) 7'b1011110;
  assign _0730_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:665" *) 7'b1011110;
  assign _0731_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:668" *) 7'b1011111;
  assign _0732_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:670" *) 7'b1011111;
  assign _0733_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:673" *) 7'b1100000;
  assign _0734_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:675" *) 7'b1100000;
  assign _0735_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:678" *) 7'b1100001;
  assign _0736_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:680" *) 7'b1100001;
  assign _0737_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:683" *) 7'b1100010;
  assign _0738_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:685" *) 7'b1100010;
  assign _0739_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:688" *) 7'b1100011;
  assign _0740_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:690" *) 7'b1100011;
  assign _0741_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:693" *) 7'b1100100;
  assign _0742_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:695" *) 7'b1100100;
  assign _0743_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:698" *) 7'b1100101;
  assign _0744_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:700" *) 7'b1100101;
  assign _0745_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:703" *) 7'b1100110;
  assign _0746_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:705" *) 7'b1100110;
  assign _0747_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:708" *) 7'b1100111;
  assign _0748_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:710" *) 7'b1100111;
  assign _0749_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:713" *) 7'b1101000;
  assign _0750_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:715" *) 7'b1101000;
  assign _0751_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:718" *) 7'b1101001;
  assign _0752_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:720" *) 7'b1101001;
  assign _0753_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:723" *) 7'b1101010;
  assign _0754_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:725" *) 7'b1101010;
  assign _0755_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:728" *) 7'b1101011;
  assign _0756_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:730" *) 7'b1101011;
  assign _0757_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:733" *) 7'b1101100;
  assign _0758_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:735" *) 7'b1101100;
  assign _0759_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:738" *) 7'b1101101;
  assign _0760_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:740" *) 7'b1101101;
  assign _0761_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:743" *) 7'b1101110;
  assign _0762_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:745" *) 7'b1101110;
  assign _0763_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:748" *) 7'b1101111;
  assign _0764_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:750" *) 7'b1101111;
  assign _0765_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:753" *) 7'b1110000;
  assign _0766_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:755" *) 7'b1110000;
  assign _0767_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:758" *) 7'b1110001;
  assign _0768_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:760" *) 7'b1110001;
  assign _0769_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:763" *) 7'b1110010;
  assign _0770_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:765" *) 7'b1110010;
  assign _0771_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:768" *) 7'b1110011;
  assign _0772_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:770" *) 7'b1110011;
  assign _0773_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:773" *) 7'b1110100;
  assign _0774_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:775" *) 7'b1110100;
  assign _0775_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:778" *) 7'b1110101;
  assign _0776_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:780" *) 7'b1110101;
  assign _0777_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:783" *) 7'b1110110;
  assign _0778_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:785" *) 7'b1110110;
  assign _0779_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:788" *) 7'b1110111;
  assign _0780_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:790" *) 7'b1110111;
  assign _0781_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:793" *) 7'b1111000;
  assign _0782_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:795" *) 7'b1111000;
  assign _0783_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:798" *) 7'b1111001;
  assign _0784_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:800" *) 7'b1111001;
  assign _0785_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:803" *) 7'b1111010;
  assign _0786_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:805" *) 7'b1111010;
  assign _0787_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:808" *) 7'b1111011;
  assign _0788_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:810" *) 7'b1111011;
  assign _0789_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:813" *) 7'b1111100;
  assign _0790_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:815" *) 7'b1111100;
  assign _0791_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:818" *) 7'b1111101;
  assign _0792_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:820" *) 7'b1111101;
  assign _0793_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:823" *) 7'b1111110;
  assign _0794_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:825" *) 7'b1111110;
  assign _0795_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:828" *) 7'b1111111;
  assign _0796_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:830" *) 7'b1111111;
  assign _0797_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:833" *) 8'b10000000;
  assign _0798_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:835" *) 8'b10000000;
  assign _0799_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:838" *) 8'b10000001;
  assign _0800_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:840" *) 8'b10000001;
  assign _0801_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:843" *) 8'b10000010;
  assign _0802_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:845" *) 8'b10000010;
  assign _0803_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:848" *) 8'b10000011;
  assign _0804_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:850" *) 8'b10000011;
  assign _0805_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:853" *) 8'b10000100;
  assign _0806_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:855" *) 8'b10000100;
  assign _0807_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:858" *) 8'b10000101;
  assign _0808_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:860" *) 8'b10000101;
  assign _0809_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:863" *) 8'b10000110;
  assign _0810_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:865" *) 8'b10000110;
  assign _0811_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:868" *) 8'b10000111;
  assign _0812_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:870" *) 8'b10000111;
  assign _0813_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:873" *) 8'b10001000;
  assign _0814_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:875" *) 8'b10001000;
  assign _0815_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:878" *) 8'b10001001;
  assign _0816_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:880" *) 8'b10001001;
  assign _0817_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:883" *) 8'b10001010;
  assign _0818_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:885" *) 8'b10001010;
  assign _0819_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:888" *) 8'b10001011;
  assign _0820_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:890" *) 8'b10001011;
  assign _0821_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:893" *) 8'b10001100;
  assign _0822_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:895" *) 8'b10001100;
  assign _0823_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:898" *) 8'b10001101;
  assign _0824_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:900" *) 8'b10001101;
  assign _0825_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:903" *) 8'b10001110;
  assign _0826_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:905" *) 8'b10001110;
  assign _0827_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:908" *) 8'b10001111;
  assign _0828_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:910" *) 8'b10001111;
  assign _0829_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:913" *) 8'b10010000;
  assign _0830_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:915" *) 8'b10010000;
  assign _0831_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:918" *) 8'b10010001;
  assign _0832_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:920" *) 8'b10010001;
  assign _0833_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:923" *) 8'b10010010;
  assign _0834_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:925" *) 8'b10010010;
  assign _0835_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:928" *) 8'b10010011;
  assign _0836_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:930" *) 8'b10010011;
  assign _0837_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:933" *) 8'b10010100;
  assign _0838_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:935" *) 8'b10010100;
  assign _0839_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:938" *) 8'b10010101;
  assign _0840_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:940" *) 8'b10010101;
  assign _0841_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:943" *) 8'b10010110;
  assign _0842_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:945" *) 8'b10010110;
  assign _0843_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:948" *) 8'b10010111;
  assign _0844_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:950" *) 8'b10010111;
  assign _0845_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:953" *) 8'b10011000;
  assign _0846_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:955" *) 8'b10011000;
  assign _0847_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:958" *) 8'b10011001;
  assign _0848_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:960" *) 8'b10011001;
  assign _0849_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:963" *) 8'b10011010;
  assign _0850_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:965" *) 8'b10011010;
  assign _0851_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:968" *) 8'b10011011;
  assign wr_count_next_no_wr_popping_is_256 = wr_count_next_no_wr_popping == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:97" *) 9'b100000000;
  assign _0852_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:970" *) 8'b10011011;
  assign _0853_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:973" *) 8'b10011100;
  assign _0854_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:975" *) 8'b10011100;
  assign _0855_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:978" *) 8'b10011101;
  assign _0856_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:980" *) 8'b10011101;
  assign _0857_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:983" *) 8'b10011110;
  assign _0858_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:985" *) 8'b10011110;
  assign _0859_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:988" *) 8'b10011111;
  assign _0860_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:990" *) 8'b10011111;
  assign _0861_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:993" *) 8'b10100000;
  assign _0862_ = adr_ram_wr_data == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:995" *) 8'b10100000;
  assign _0863_ = rd_adr_dly == (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:998" *) 8'b10100001;
  assign _0864_ = cq_rd_count0 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2122" *) 1'b1;
  assign _0865_ = cq_rd_count1 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2123" *) 1'b1;
  assign _0866_ = cq_rd_count2 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2124" *) 1'b1;
  assign _0867_ = cq_rd_count3 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2125" *) 1'b1;
  assign _0868_ = cq_rd_count4 > (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2126" *) 1'b1;
  assign _0869_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1000" *) _0324_;
  assign _0870_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1003" *) _0325_;
  assign _0871_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1005" *) _0326_;
  assign _0872_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1008" *) _0327_;
  assign _0873_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1010" *) _0328_;
  assign _0874_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1013" *) _0329_;
  assign _0875_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1015" *) _0330_;
  assign _0876_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1018" *) _0331_;
  assign _0877_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1020" *) _0332_;
  assign _0878_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1023" *) _0333_;
  assign _0879_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1025" *) _0334_;
  assign _0880_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1028" *) _0335_;
  assign _0881_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1030" *) _0336_;
  assign _0882_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1033" *) _0337_;
  assign _0883_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1035" *) _0338_;
  assign _0884_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1038" *) _0339_;
  assign _0885_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1040" *) _0340_;
  assign _0886_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1043" *) _0341_;
  assign _0887_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1045" *) _0342_;
  assign _0888_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1048" *) _0343_;
  assign _0889_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1050" *) _0344_;
  assign _0890_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1053" *) _0345_;
  assign _0891_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1055" *) _0346_;
  assign _0892_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1058" *) _0347_;
  assign _0893_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1060" *) _0348_;
  assign _0894_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1063" *) _0349_;
  assign _0895_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1065" *) _0350_;
  assign _0896_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1068" *) _0351_;
  assign _0897_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1070" *) _0352_;
  assign _0898_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1073" *) _0353_;
  assign _0899_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1075" *) _0354_;
  assign _0900_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1078" *) _0355_;
  assign _0901_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1080" *) _0356_;
  assign _0902_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1083" *) _0357_;
  assign _0903_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1085" *) _0358_;
  assign _0904_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1088" *) _0359_;
  assign _0905_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1090" *) _0360_;
  assign _0906_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1093" *) _0361_;
  assign _0907_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1095" *) _0362_;
  assign _0908_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1098" *) _0363_;
  assign _0909_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1100" *) _0364_;
  assign _0910_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1103" *) _0365_;
  assign _0911_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1105" *) _0366_;
  assign _0912_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1108" *) _0367_;
  assign _0913_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1110" *) _0368_;
  assign _0914_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1113" *) _0369_;
  assign _0915_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1115" *) _0370_;
  assign _0916_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1118" *) _0371_;
  assign _0917_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1120" *) _0372_;
  assign _0918_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1123" *) _0373_;
  assign _0919_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1125" *) _0374_;
  assign _0920_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1128" *) _0375_;
  assign _0921_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1130" *) _0376_;
  assign _0922_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1133" *) _0377_;
  assign _0923_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1135" *) _0378_;
  assign _0924_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1138" *) _0379_;
  assign _0925_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1140" *) _0380_;
  assign _0926_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1143" *) _0381_;
  assign _0927_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1145" *) _0382_;
  assign _0928_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1148" *) _0383_;
  assign _0929_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1150" *) _0384_;
  assign _0930_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1153" *) _0385_;
  assign _0931_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1155" *) _0386_;
  assign _0932_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1158" *) _0387_;
  assign _0933_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1160" *) _0388_;
  assign _0934_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1163" *) _0389_;
  assign _0935_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1165" *) _0390_;
  assign _0936_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1168" *) _0391_;
  assign _0937_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1170" *) _0392_;
  assign _0938_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1173" *) _0393_;
  assign _0939_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1175" *) _0394_;
  assign _0940_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1178" *) _0395_;
  assign _0941_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1180" *) _0396_;
  assign _0942_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1183" *) _0397_;
  assign _0943_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1185" *) _0398_;
  assign _0944_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1188" *) _0399_;
  assign _0945_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1190" *) _0400_;
  assign _0946_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1193" *) _0401_;
  assign _0947_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1195" *) _0402_;
  assign _0948_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1198" *) _0403_;
  assign _0949_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1200" *) _0404_;
  assign _0950_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1203" *) _0405_;
  assign _0951_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1205" *) _0406_;
  assign _0952_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1208" *) _0407_;
  assign _0953_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1210" *) _0408_;
  assign _0954_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1213" *) _0409_;
  assign _0955_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1215" *) _0410_;
  assign _0956_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1218" *) _0411_;
  assign _0957_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1220" *) _0412_;
  assign _0958_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1223" *) _0413_;
  assign _0959_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1225" *) _0414_;
  assign _0960_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1228" *) _0415_;
  assign _0961_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1230" *) _0416_;
  assign _0962_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1233" *) _0417_;
  assign _0963_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1235" *) _0418_;
  assign _0964_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1238" *) _0419_;
  assign _0965_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1240" *) _0420_;
  assign _0966_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1243" *) _0421_;
  assign _0967_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1245" *) _0422_;
  assign _0968_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1248" *) _0423_;
  assign _0969_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1250" *) _0424_;
  assign _0970_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1253" *) _0425_;
  assign _0971_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1255" *) _0426_;
  assign _0972_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1258" *) _0427_;
  assign _0973_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1260" *) _0428_;
  assign _0974_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1263" *) _0429_;
  assign _0975_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1265" *) _0430_;
  assign _0976_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1268" *) _0431_;
  assign _0977_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1270" *) _0432_;
  assign _0978_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1273" *) _0433_;
  assign _0979_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1275" *) _0434_;
  assign _0980_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1278" *) _0435_;
  assign _0981_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1280" *) _0436_;
  assign _0982_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1283" *) _0437_;
  assign _0983_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1285" *) _0438_;
  assign _0984_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1288" *) _0439_;
  assign _0985_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1290" *) _0440_;
  assign _0986_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1293" *) _0441_;
  assign _0987_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1295" *) _0442_;
  assign _0988_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1298" *) _0443_;
  assign _0989_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1300" *) _0444_;
  assign _0990_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1303" *) _0445_;
  assign _0991_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1305" *) _0446_;
  assign _0992_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1308" *) _0447_;
  assign _0993_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1310" *) _0448_;
  assign _0994_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1313" *) _0449_;
  assign _0995_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1315" *) _0450_;
  assign _0996_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1318" *) _0451_;
  assign _0997_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1320" *) _0452_;
  assign _0998_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1323" *) _0453_;
  assign _0999_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1325" *) _0454_;
  assign _1000_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1328" *) _0455_;
  assign _1001_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1330" *) _0456_;
  assign _1002_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1333" *) _0457_;
  assign _1003_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1335" *) _0458_;
  assign _1004_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1338" *) _0459_;
  assign _1005_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1340" *) _0460_;
  assign _1006_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1343" *) _0461_;
  assign _1007_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1345" *) _0462_;
  assign _1008_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1348" *) _0463_;
  assign _1009_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1350" *) _0464_;
  assign _1010_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1353" *) _0465_;
  assign _1011_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1355" *) _0466_;
  assign _1012_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1358" *) _0467_;
  assign _1013_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1360" *) _0468_;
  assign _1014_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1363" *) _0469_;
  assign _1015_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1365" *) _0470_;
  assign _1016_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1368" *) _0471_;
  assign _1017_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1370" *) _0472_;
  assign _1018_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1373" *) _0473_;
  assign _1019_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1375" *) _0474_;
  assign _1020_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1378" *) _0475_;
  assign _1021_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1380" *) _0476_;
  assign _1022_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1383" *) _0477_;
  assign _1023_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1385" *) _0478_;
  assign _1024_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1388" *) _0479_;
  assign _1025_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1390" *) _0480_;
  assign _1026_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1393" *) _0481_;
  assign _1027_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1395" *) _0482_;
  assign _1028_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1398" *) _0483_;
  assign rd_pushing = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:140" *) _1549_;
  assign _1029_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1400" *) _0484_;
  assign _1030_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1403" *) _0485_;
  assign _1031_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1405" *) _0486_;
  assign _1032_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1408" *) _0487_;
  assign _1033_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1410" *) _0488_;
  assign _1034_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1413" *) _0489_;
  assign _1035_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1415" *) _0490_;
  assign _1036_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1418" *) _0491_;
  assign _1037_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1420" *) _0492_;
  assign _1038_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1423" *) _0493_;
  assign _1039_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1425" *) _0494_;
  assign _1040_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1428" *) _0495_;
  assign _1041_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1430" *) _0496_;
  assign _1042_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1433" *) _0497_;
  assign _1043_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1435" *) _0498_;
  assign _1044_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1438" *) _0499_;
  assign _1045_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1440" *) _0500_;
  assign _1046_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1443" *) _0501_;
  assign _1047_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1445" *) _0502_;
  assign _1048_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1448" *) _0503_;
  assign _1049_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1450" *) _0504_;
  assign _1050_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1453" *) _0505_;
  assign _1051_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1455" *) _0506_;
  assign _1052_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1458" *) _0507_;
  assign _1053_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1460" *) _0508_;
  assign _1054_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1463" *) _0509_;
  assign _1055_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1465" *) _0510_;
  assign _1056_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:193" *) _0511_;
  assign _1057_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:195" *) _0512_;
  assign _1058_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:198" *) _0513_;
  assign rd_pushing0 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1985" *) _0514_;
  assign rd_pushing1 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1986" *) _0515_;
  assign rd_pushing2 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1987" *) _0516_;
  assign rd_pushing3 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1988" *) _0517_;
  assign rd_pushing4 = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1989" *) _0518_;
  assign rd_take0 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1999" *) _0519_;
  assign _1059_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:200" *) _0520_;
  assign rd_take1 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2000" *) _0521_;
  assign rd_take2 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2001" *) _0522_;
  assign rd_take3 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2002" *) _0523_;
  assign rd_take4 = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2003" *) _0524_;
  assign _1060_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:203" *) _0525_;
  assign _1061_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:205" *) _0526_;
  assign _1062_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:208" *) _0527_;
  assign _1063_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:210" *) _0528_;
  assign update_head_next[0] = rd_take0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2122" *) _0864_;
  assign update_head_next[1] = rd_take1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2123" *) _0865_;
  assign update_head_next[2] = rd_take2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2124" *) _0866_;
  assign update_head_next[3] = rd_take3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2125" *) _0867_;
  assign update_head_next[4] = rd_take4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2126" *) _0868_;
  assign _1064_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:213" *) _0529_;
  assign _1065_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:215" *) _0530_;
  assign _1066_ = rd_pushing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2152" *) _0531_;
  assign _1067_ = rd_pushing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *) rd_take0;
  assign _1068_ = _1067_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *) _0532_;
  assign _1069_ = rd_pushing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2167" *) _0533_;
  assign _1070_ = rd_pushing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *) rd_take1;
  assign _1071_ = _1070_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *) _0534_;
  assign _1072_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:218" *) _0535_;
  assign _1073_ = rd_pushing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2182" *) _0536_;
  assign _1074_ = rd_pushing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *) rd_take2;
  assign _1075_ = _1074_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *) _0537_;
  assign _1076_ = rd_pushing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2197" *) _0538_;
  assign _1077_ = rd_pushing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *) rd_take3;
  assign _1078_ = _1077_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *) _0539_;
  assign _1079_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:220" *) _0540_;
  assign _1080_ = rd_pushing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2212" *) _0541_;
  assign _1081_ = rd_pushing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *) rd_take4;
  assign _1082_ = _1081_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *) _0542_;
  assign _1083_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:223" *) _0543_;
  assign _1084_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2244" *) _1707_;
  assign _1085_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2245" *) _1708_;
  assign _1086_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2246" *) _1709_;
  assign _1087_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2247" *) _1710_;
  assign _1088_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2248" *) _1711_;
  assign _1089_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:225" *) _0544_;
  assign _1090_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2256" *) _1707_;
  assign _1091_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2257" *) _1708_;
  assign _1092_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2258" *) _1709_;
  assign _1093_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2259" *) _1710_;
  assign _1094_ = cq_rd_take && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2260" *) _1711_;
  assign _1095_ = rd_take_n_dly[0] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2268" *) update_head[0];
  assign _1096_ = rd_take_n_dly[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2269" *) update_head[1];
  assign _1097_ = rd_take_n_dly[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2270" *) update_head[2];
  assign _1098_ = rd_take_n_dly[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2271" *) update_head[3];
  assign _1099_ = rd_take_n_dly[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2272" *) update_head[4];
  assign _1100_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:228" *) _0545_;
  assign _1101_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:230" *) _0546_;
  assign _1102_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:233" *) _0547_;
  assign _1103_ = cq_rd0_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) cq_rd0_prdy;
  assign _1104_ = _1103_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) _1551_;
  assign _1105_ = _1603_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) _1604_;
  assign _1106_ = _1103_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2339" *) rd_skid0_1_vld;
  assign _1107_ = _1103_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *) _1552_;
  assign _1108_ = _1603_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *) _1605_;
  assign _1109_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:235" *) _0548_;
  assign _1110_ = _1103_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2351" *) rd_skid0_2_vld;
  assign _1111_ = _1603_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *) rd_skid0_0_vld;
  assign _1112_ = _1111_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *) rd_skid0_1_vld;
  assign _1113_ = _1112_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *) _1606_;
  assign _1114_ = rd_bypassing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *) rd_skid0_0_vld;
  assign _1115_ = rd_skid0_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *) _1603_;
  assign _1116_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:238" *) _0549_;
  assign _1117_ = rd_skid0_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2380" *) _1603_;
  assign _1118_ = _1552_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) _1554_;
  assign cq_rd_take_elig[0] = _1615_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) _1616_;
  assign wr_reserving = cq_wr_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) cq_wr_prdy;
  assign _1119_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) _0514_;
  assign _1120_ = _1119_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) _0550_;
  assign _1121_ = _1120_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) _1555_;
  assign rd_pre_bypassing0 = _1121_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) _1617_;
  assign _1122_ = _1556_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) rd_skid0_0_vld;
  assign _1123_ = _1122_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) rd_skid0_1_vld;
  assign _1124_ = rd_pre_bypassing0 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) _1619_;
  assign rd_bypassing0 = _1124_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) _1554_;
  assign _1125_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:240" *) _0551_;
  assign _1126_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:243" *) _0552_;
  assign _1127_ = cq_rd1_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) cq_rd1_prdy;
  assign _1128_ = _1127_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) _1559_;
  assign _1129_ = _1620_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) _1621_;
  assign _1130_ = _1127_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2435" *) rd_skid1_1_vld;
  assign _1131_ = _1127_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *) _1560_;
  assign _1132_ = _1620_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *) _1622_;
  assign _1133_ = _1127_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2447" *) rd_skid1_2_vld;
  assign _1134_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:245" *) _0553_;
  assign _1135_ = _1620_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *) rd_skid1_0_vld;
  assign _1136_ = _1135_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *) rd_skid1_1_vld;
  assign _1137_ = _1136_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *) _1623_;
  assign _1138_ = rd_bypassing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *) rd_skid1_0_vld;
  assign _1139_ = rd_skid1_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *) _1620_;
  assign _1140_ = rd_skid1_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2476" *) _1620_;
  assign _1141_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:248" *) _0554_;
  assign _1142_ = _1560_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) _1562_;
  assign cq_rd_take_elig[1] = _1632_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) _1633_;
  assign _1143_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) _0515_;
  assign _1144_ = _1143_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) _0555_;
  assign _1145_ = _1144_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) _1563_;
  assign rd_pre_bypassing1 = _1145_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) _1634_;
  assign _1146_ = _1564_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) rd_skid1_0_vld;
  assign _1147_ = _1146_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) rd_skid1_1_vld;
  assign _1148_ = rd_pre_bypassing1 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) _1636_;
  assign rd_bypassing1 = _1148_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) _1562_;
  assign _1149_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:250" *) _0556_;
  assign _1150_ = cq_rd2_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) cq_rd2_prdy;
  assign _1151_ = _1150_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) _1567_;
  assign _1152_ = _1637_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) _1638_;
  assign _1153_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:253" *) _0557_;
  assign _1154_ = _1150_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2531" *) rd_skid2_1_vld;
  assign _1155_ = _1150_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *) _1568_;
  assign _1156_ = _1637_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *) _1639_;
  assign _1157_ = _1150_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2543" *) rd_skid2_2_vld;
  assign _1158_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:255" *) _0558_;
  assign _1159_ = _1637_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *) rd_skid2_0_vld;
  assign _1160_ = _1159_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *) rd_skid2_1_vld;
  assign _1161_ = _1160_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *) _1640_;
  assign _1162_ = rd_bypassing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *) rd_skid2_0_vld;
  assign _1163_ = rd_skid2_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *) _1637_;
  assign _1164_ = rd_skid2_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2572" *) _1637_;
  assign _1165_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:258" *) _0559_;
  assign _1166_ = _1568_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) _1570_;
  assign cq_rd_take_elig[2] = _1649_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) _1650_;
  assign _1167_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) _0516_;
  assign _1168_ = _1167_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) _0560_;
  assign _1169_ = _1168_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) _1571_;
  assign rd_pre_bypassing2 = _1169_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) _1651_;
  assign _1170_ = _1572_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) rd_skid2_0_vld;
  assign _1171_ = _1170_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) rd_skid2_1_vld;
  assign _1172_ = rd_pre_bypassing2 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) _1653_;
  assign rd_bypassing2 = _1172_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) _1570_;
  assign _1173_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:260" *) _0561_;
  assign _1174_ = cq_rd3_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) cq_rd3_prdy;
  assign _1175_ = _1174_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) _1575_;
  assign _1176_ = _1654_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) _1655_;
  assign _1177_ = _1174_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2627" *) rd_skid3_1_vld;
  assign _1178_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:263" *) _0562_;
  assign _1179_ = _1174_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *) _1576_;
  assign _1180_ = _1654_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *) _1656_;
  assign _1181_ = _1174_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2639" *) rd_skid3_2_vld;
  assign _1182_ = _1654_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *) rd_skid3_0_vld;
  assign _1183_ = _1182_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *) rd_skid3_1_vld;
  assign _1184_ = _1183_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *) _1657_;
  assign _1185_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:265" *) _0563_;
  assign _1186_ = rd_bypassing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *) rd_skid3_0_vld;
  assign _1187_ = rd_skid3_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *) _1654_;
  assign _1188_ = rd_skid3_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2668" *) _1654_;
  assign _1189_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:268" *) _0564_;
  assign _1190_ = _1576_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) _1578_;
  assign cq_rd_take_elig[3] = _1666_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) _1667_;
  assign _1191_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) _0517_;
  assign _1192_ = _1191_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) _0565_;
  assign _1193_ = _1192_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) _1579_;
  assign rd_pre_bypassing3 = _1193_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) _1668_;
  assign _1194_ = _1580_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) rd_skid3_0_vld;
  assign _1195_ = _1194_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) rd_skid3_1_vld;
  assign _1196_ = rd_pre_bypassing3 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) _1670_;
  assign rd_bypassing3 = _1196_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) _1578_;
  assign _1197_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:270" *) _0566_;
  assign _1198_ = cq_rd4_pvld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) cq_rd4_prdy;
  assign _1199_ = _1198_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) _1583_;
  assign _1200_ = _1671_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) _1672_;
  assign _1201_ = _1198_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2723" *) rd_skid4_1_vld;
  assign _1202_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:273" *) _0567_;
  assign _1203_ = _1198_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *) _1584_;
  assign _1204_ = _1671_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *) _1673_;
  assign _1205_ = _1198_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2735" *) rd_skid4_2_vld;
  assign _1206_ = _1671_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *) rd_skid4_0_vld;
  assign _1207_ = _1206_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *) rd_skid4_1_vld;
  assign _1208_ = _1207_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *) _1674_;
  assign _1209_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:275" *) _0568_;
  assign _1210_ = rd_bypassing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *) rd_skid4_0_vld;
  assign _1211_ = rd_skid4_1_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *) _1671_;
  assign _1212_ = rd_skid4_2_vld && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2764" *) _1671_;
  assign _1213_ = _1584_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) _1586_;
  assign cq_rd_take_elig[4] = _1683_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) _1684_;
  assign _1214_ = wr_reserving && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) _0518_;
  assign _1215_ = _1214_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) _0569_;
  assign _1216_ = _1215_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) _1587_;
  assign rd_pre_bypassing4 = _1216_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) _1685_;
  assign _1217_ = _1588_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) rd_skid4_0_vld;
  assign _1218_ = _1217_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) rd_skid4_1_vld;
  assign _1219_ = rd_pre_bypassing4 && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) _1687_;
  assign rd_bypassing4 = _1219_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) _1586_;
  assign _1220_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:278" *) _0570_;
  assign _1221_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:280" *) _0571_;
  assign _1222_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *) _0572_;
  assign cq_rd_take_thread_id_is_1[4] = _1222_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *) _1590_;
  assign _1223_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *) _0573_;
  assign _1224_ = _1223_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *) _1591_;
  assign cq_rd_take_thread_id_is_1[3] = _1224_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *) _1590_;
  assign _1225_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *) _0574_;
  assign _1226_ = _1225_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *) _1592_;
  assign _1227_ = _1226_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *) _1591_;
  assign cq_rd_take_thread_id_is_1[2] = _1227_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *) _1590_;
  assign _1228_ = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) _0575_;
  assign _1229_ = _1228_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) _1593_;
  assign _1230_ = _1229_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) _1592_;
  assign _1231_ = _1230_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) _1591_;
  assign cq_rd_take_thread_id_is_1[1] = _1231_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) _1590_;
  assign cq_rd_take_thread_id_is_1[0] = cq_rd_take_elig[1] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2806" *) _0576_;
  assign _1232_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *) _0572_;
  assign _1233_ = _1232_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *) _1590_;
  assign cq_rd_take_thread_id_is_2[4] = _1233_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *) _1594_;
  assign _1234_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *) _0573_;
  assign _1235_ = _1234_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *) _1591_;
  assign _1236_ = _1235_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *) _1590_;
  assign cq_rd_take_thread_id_is_2[3] = _1236_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2809" *) _1594_;
  assign _1237_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *) _0574_;
  assign _1238_ = _1237_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *) _1592_;
  assign _1239_ = _1238_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *) _1591_;
  assign _1240_ = _1239_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *) _1590_;
  assign cq_rd_take_thread_id_is_2[2] = _1240_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2810" *) _1594_;
  assign cq_rd_take_thread_id_is_2[1] = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2811" *) _0575_;
  assign _1241_ = cq_rd_take_elig[2] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2812" *) _0576_;
  assign cq_rd_take_thread_id_is_2[0] = _1241_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2812" *) _1594_;
  assign _1242_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *) _0572_;
  assign _1243_ = _1242_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *) _1590_;
  assign _1244_ = _1243_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *) _1594_;
  assign cq_rd_take_thread_id_is_3[4] = _1244_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2814" *) _1593_;
  assign _1245_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *) _0573_;
  assign _1246_ = _1245_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *) _1591_;
  assign _1247_ = _1246_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *) _1590_;
  assign _1248_ = _1247_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *) _1594_;
  assign cq_rd_take_thread_id_is_3[3] = _1248_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2815" *) _1593_;
  assign cq_rd_take_thread_id_is_3[2] = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2816" *) _0574_;
  assign _1249_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2817" *) _0575_;
  assign cq_rd_take_thread_id_is_3[1] = _1249_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2817" *) _1593_;
  assign _1250_ = cq_rd_take_elig[3] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2818" *) _0576_;
  assign _1251_ = _1250_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2818" *) _1594_;
  assign cq_rd_take_thread_id_is_3[0] = _1251_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2818" *) _1593_;
  assign _1252_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *) _0572_;
  assign _1253_ = _1252_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *) _1590_;
  assign _1254_ = _1253_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *) _1594_;
  assign _1255_ = _1254_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *) _1593_;
  assign cq_rd_take_thread_id_is_4[4] = _1255_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2820" *) _1592_;
  assign cq_rd_take_thread_id_is_4[3] = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2821" *) _0573_;
  assign _1256_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2822" *) _0574_;
  assign cq_rd_take_thread_id_is_4[2] = _1256_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2822" *) _1592_;
  assign _1257_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2823" *) _0575_;
  assign _1258_ = _1257_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2823" *) _1593_;
  assign cq_rd_take_thread_id_is_4[1] = _1258_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2823" *) _1592_;
  assign _1259_ = cq_rd_take_elig[4] && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *) _0576_;
  assign _1260_ = _1259_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *) _1594_;
  assign _1261_ = _1260_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *) _1593_;
  assign cq_rd_take_thread_id_is_4[0] = _1261_ && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2824" *) _1592_;
  assign _1262_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:283" *) _0577_;
  assign _1263_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:285" *) _0578_;
  assign _1264_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:288" *) _0579_;
  assign _1265_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:290" *) _0580_;
  assign _1266_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:293" *) _0581_;
  assign _1267_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:295" *) _0582_;
  assign _1268_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:298" *) _0583_;
  assign _1269_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:300" *) _0584_;
  assign _1270_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:303" *) _0585_;
  assign _1271_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:305" *) _0586_;
  assign _1272_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:308" *) _0587_;
  assign _1273_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:310" *) _0588_;
  assign _1274_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:313" *) _0589_;
  assign _1275_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:315" *) _0590_;
  assign _1276_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:318" *) _0591_;
  assign _1277_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:320" *) _0592_;
  assign _1278_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:323" *) _0593_;
  assign _1279_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:325" *) _0594_;
  assign _1280_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:328" *) _0595_;
  assign _1281_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:330" *) _0596_;
  assign _1282_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:333" *) _0597_;
  assign _1283_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:335" *) _0598_;
  assign _1284_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:338" *) _0599_;
  assign _1285_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:340" *) _0600_;
  assign _1286_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:343" *) _0601_;
  assign _1287_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:345" *) _0602_;
  assign _1288_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:348" *) _0603_;
  assign _1289_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:350" *) _0604_;
  assign _1290_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:353" *) _0605_;
  assign _1291_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:355" *) _0606_;
  assign _1292_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:358" *) _0607_;
  assign _1293_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:360" *) _0608_;
  assign _1294_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:363" *) _0609_;
  assign _1295_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:365" *) _0610_;
  assign _1296_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:368" *) _0611_;
  assign _1297_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:370" *) _0612_;
  assign _1298_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:373" *) _0613_;
  assign _1299_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:375" *) _0614_;
  assign _1300_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:378" *) _0615_;
  assign _1301_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:380" *) _0616_;
  assign _1302_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:383" *) _0617_;
  assign _1303_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:385" *) _0618_;
  assign _1304_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:388" *) _0619_;
  assign _1305_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:390" *) _0620_;
  assign _1306_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:393" *) _0621_;
  assign _1307_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:395" *) _0622_;
  assign _1308_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:398" *) _0623_;
  assign _1309_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:400" *) _0624_;
  assign _1310_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:403" *) _0625_;
  assign _1311_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:405" *) _0626_;
  assign _1312_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:408" *) _0627_;
  assign _1313_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:410" *) _0628_;
  assign _1314_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:413" *) _0629_;
  assign _1315_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:415" *) _0630_;
  assign _1316_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:418" *) _0631_;
  assign _1317_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:420" *) _0632_;
  assign _1318_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:423" *) _0633_;
  assign _1319_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:425" *) _0634_;
  assign _1320_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:428" *) _0635_;
  assign _1321_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:430" *) _0636_;
  assign _1322_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:433" *) _0637_;
  assign _1323_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:435" *) _0638_;
  assign _1324_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:438" *) _0639_;
  assign _1325_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:440" *) _0640_;
  assign _1326_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:443" *) _0641_;
  assign _1327_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:445" *) _0642_;
  assign _1328_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:448" *) _0643_;
  assign _1329_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:450" *) _0644_;
  assign _1330_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:453" *) _0645_;
  assign _1331_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:455" *) _0646_;
  assign _1332_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:458" *) _0647_;
  assign _1333_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:460" *) _0648_;
  assign _1334_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:463" *) _0649_;
  assign _1335_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:465" *) _0650_;
  assign _1336_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:468" *) _0651_;
  assign _1337_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:470" *) _0652_;
  assign _1338_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:473" *) _0653_;
  assign _1339_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:475" *) _0654_;
  assign _1340_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:478" *) _0655_;
  assign _1341_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:480" *) _0656_;
  assign _1342_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:483" *) _0657_;
  assign _1343_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:485" *) _0658_;
  assign _1344_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:488" *) _0659_;
  assign _1345_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:490" *) _0660_;
  assign _1346_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:493" *) _0661_;
  assign _1347_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:495" *) _0662_;
  assign _1348_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:498" *) _0663_;
  assign _1349_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:500" *) _0664_;
  assign _1350_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:503" *) _0665_;
  assign _1351_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:505" *) _0666_;
  assign _1352_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:508" *) _0667_;
  assign _1353_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:510" *) _0668_;
  assign _1354_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:513" *) _0669_;
  assign _1355_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:515" *) _0670_;
  assign _1356_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:518" *) _0671_;
  assign _1357_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:520" *) _0672_;
  assign _1358_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:523" *) _0673_;
  assign _1359_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:525" *) _0674_;
  assign _1360_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:528" *) _0675_;
  assign _1361_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:530" *) _0676_;
  assign _1362_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:533" *) _0677_;
  assign _1363_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:535" *) _0678_;
  assign _1364_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:538" *) _0679_;
  assign _1365_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:540" *) _0680_;
  assign _1366_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:543" *) _0681_;
  assign _1367_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:545" *) _0682_;
  assign _1368_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:548" *) _0683_;
  assign _1369_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:550" *) _0684_;
  assign _1370_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:553" *) _0685_;
  assign _1371_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:555" *) _0686_;
  assign _1372_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:558" *) _0687_;
  assign _1373_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:560" *) _0688_;
  assign _1374_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:563" *) _0689_;
  assign _1375_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:565" *) _0690_;
  assign _1376_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:568" *) _0691_;
  assign _1377_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:570" *) _0692_;
  assign _1378_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:573" *) _0693_;
  assign _1379_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:575" *) _0694_;
  assign _1380_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:578" *) _0695_;
  assign _1381_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:580" *) _0696_;
  assign _1382_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:583" *) _0697_;
  assign _1383_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:585" *) _0698_;
  assign _1384_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:588" *) _0699_;
  assign _1385_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:590" *) _0700_;
  assign _1386_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:593" *) _0701_;
  assign _1387_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:595" *) _0702_;
  assign _1388_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:598" *) _0703_;
  assign _1389_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:600" *) _0704_;
  assign _1390_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:603" *) _0705_;
  assign _1391_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:605" *) _0706_;
  assign _1392_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:608" *) _0707_;
  assign _1393_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:610" *) _0708_;
  assign _1394_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:613" *) _0709_;
  assign _1395_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:615" *) _0710_;
  assign _1396_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:618" *) _0711_;
  assign _1397_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:620" *) _0712_;
  assign _1398_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:623" *) _0713_;
  assign _1399_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:625" *) _0714_;
  assign _1400_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:628" *) _0715_;
  assign _1401_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:630" *) _0716_;
  assign _1402_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:633" *) _0717_;
  assign _1403_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:635" *) _0718_;
  assign _1404_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:638" *) _0719_;
  assign _1405_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:640" *) _0720_;
  assign _1406_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:643" *) _0721_;
  assign _1407_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:645" *) _0722_;
  assign _1408_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:648" *) _0723_;
  assign _1409_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:650" *) _0724_;
  assign _1410_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:653" *) _0725_;
  assign _1411_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:655" *) _0726_;
  assign _1412_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:658" *) _0727_;
  assign _1413_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:660" *) _0728_;
  assign _1414_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:663" *) _0729_;
  assign _1415_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:665" *) _0730_;
  assign _1416_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:668" *) _0731_;
  assign _1417_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:670" *) _0732_;
  assign _1418_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:673" *) _0733_;
  assign _1419_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:675" *) _0734_;
  assign _1420_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:678" *) _0735_;
  assign _1421_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:680" *) _0736_;
  assign _1422_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:683" *) _0737_;
  assign _1423_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:685" *) _0738_;
  assign _1424_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:688" *) _0739_;
  assign _1425_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:690" *) _0740_;
  assign _1426_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:693" *) _0741_;
  assign _1427_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:695" *) _0742_;
  assign _1428_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:698" *) _0743_;
  assign _1429_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:700" *) _0744_;
  assign _1430_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:703" *) _0745_;
  assign _1431_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:705" *) _0746_;
  assign _1432_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:708" *) _0747_;
  assign _1433_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:710" *) _0748_;
  assign _1434_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:713" *) _0749_;
  assign _1435_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:715" *) _0750_;
  assign _1436_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:718" *) _0751_;
  assign _1437_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:720" *) _0752_;
  assign _1438_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:723" *) _0753_;
  assign _1439_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:725" *) _0754_;
  assign _1440_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:728" *) _0755_;
  assign _1441_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:730" *) _0756_;
  assign _1442_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:733" *) _0757_;
  assign _1443_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:735" *) _0758_;
  assign _1444_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:738" *) _0759_;
  assign _1445_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:740" *) _0760_;
  assign _1446_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:743" *) _0761_;
  assign _1447_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:745" *) _0762_;
  assign _1448_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:748" *) _0763_;
  assign _1449_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:750" *) _0764_;
  assign _1450_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:753" *) _0765_;
  assign _1451_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:755" *) _0766_;
  assign _1452_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:758" *) _0767_;
  assign _1453_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:760" *) _0768_;
  assign _1454_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:763" *) _0769_;
  assign _1455_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:765" *) _0770_;
  assign _1456_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:768" *) _0771_;
  assign _1457_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:770" *) _0772_;
  assign _1458_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:773" *) _0773_;
  assign _1459_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:775" *) _0774_;
  assign _1460_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:778" *) _0775_;
  assign _1461_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:780" *) _0776_;
  assign _1462_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:783" *) _0777_;
  assign _1463_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:785" *) _0778_;
  assign _1464_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:788" *) _0779_;
  assign _1465_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:790" *) _0780_;
  assign _1466_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:793" *) _0781_;
  assign _1467_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:795" *) _0782_;
  assign _1468_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:798" *) _0783_;
  assign _1469_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:800" *) _0784_;
  assign _1470_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:803" *) _0785_;
  assign _1471_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:805" *) _0786_;
  assign _1472_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:808" *) _0787_;
  assign _1473_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:810" *) _0788_;
  assign _1474_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:813" *) _0789_;
  assign _1475_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:815" *) _0790_;
  assign _1476_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:818" *) _0791_;
  assign _1477_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:820" *) _0792_;
  assign _1478_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:823" *) _0793_;
  assign _1479_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:825" *) _0794_;
  assign _1480_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:828" *) _0795_;
  assign _1481_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:830" *) _0796_;
  assign _1482_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:833" *) _0797_;
  assign _1483_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:835" *) _0798_;
  assign _1484_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:838" *) _0799_;
  assign _1485_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:840" *) _0800_;
  assign _1486_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:843" *) _0801_;
  assign _1487_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:845" *) _0802_;
  assign _1488_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:848" *) _0803_;
  assign _1489_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:850" *) _0804_;
  assign _1490_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:853" *) _0805_;
  assign _1491_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:855" *) _0806_;
  assign _1492_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:858" *) _0807_;
  assign _1493_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:860" *) _0808_;
  assign _1494_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:863" *) _0809_;
  assign _1495_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:865" *) _0810_;
  assign _1496_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:868" *) _0811_;
  assign _1497_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:870" *) _0812_;
  assign _1498_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:873" *) _0813_;
  assign _1499_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:875" *) _0814_;
  assign _1500_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:878" *) _0815_;
  assign _1501_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:880" *) _0816_;
  assign _1502_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:883" *) _0817_;
  assign _1503_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:885" *) _0818_;
  assign _1504_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:888" *) _0819_;
  assign _1505_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:890" *) _0820_;
  assign _1506_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:893" *) _0821_;
  assign _1507_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:895" *) _0822_;
  assign _1508_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:898" *) _0823_;
  assign _1509_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:900" *) _0824_;
  assign _1510_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:903" *) _0825_;
  assign _1511_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:905" *) _0826_;
  assign _1512_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:908" *) _0827_;
  assign _1513_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:910" *) _0828_;
  assign _1514_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:913" *) _0829_;
  assign _1515_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:915" *) _0830_;
  assign _1516_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:918" *) _0831_;
  assign _1517_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:920" *) _0832_;
  assign _1518_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:923" *) _0833_;
  assign _1519_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:925" *) _0834_;
  assign _1520_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:928" *) _0835_;
  assign _1521_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:930" *) _0836_;
  assign _1522_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:933" *) _0837_;
  assign _1523_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:935" *) _0838_;
  assign _1524_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:938" *) _0839_;
  assign _1525_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:940" *) _0840_;
  assign _1526_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:943" *) _0841_;
  assign _1527_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:945" *) _0842_;
  assign _1528_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:948" *) _0843_;
  assign _1529_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:950" *) _0844_;
  assign _1530_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:953" *) _0845_;
  assign _1531_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:955" *) _0846_;
  assign _1532_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:958" *) _0847_;
  assign _1533_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:960" *) _0848_;
  assign _1534_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:963" *) _0849_;
  assign _1535_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:965" *) _0850_;
  assign _1536_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:968" *) _0851_;
  assign _1537_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:970" *) _0852_;
  assign _1538_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:973" *) _0853_;
  assign _1539_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:975" *) _0854_;
  assign _1540_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:978" *) _0855_;
  assign _1541_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:980" *) _0856_;
  assign _1542_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:983" *) _0857_;
  assign _1543_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:985" *) _0858_;
  assign _1544_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:988" *) _0859_;
  assign _1545_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:990" *) _0860_;
  assign _1546_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:993" *) _0861_;
  assign _1547_ = rd_pushing && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:995" *) _0862_;
  assign _1548_ = rd_take_dly && (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:998" *) _0863_;
  assign _1549_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:140" *) wr_bypassing;
  assign index_l0_0 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1716" *) free_adr_mask[0];
  assign index_l0_1 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1717" *) free_adr_mask[2];
  assign index_l0_2 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1718" *) free_adr_mask[4];
  assign index_l0_3 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1719" *) free_adr_mask[6];
  assign index_l0_4 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1720" *) free_adr_mask[8];
  assign index_l0_5 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1721" *) free_adr_mask[10];
  assign index_l0_6 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1722" *) free_adr_mask[12];
  assign index_l0_7 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1723" *) free_adr_mask[14];
  assign index_l0_8 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1724" *) free_adr_mask[16];
  assign index_l0_9 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1725" *) free_adr_mask[18];
  assign index_l0_10 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1726" *) free_adr_mask[20];
  assign index_l0_11 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1727" *) free_adr_mask[22];
  assign index_l0_12 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1728" *) free_adr_mask[24];
  assign index_l0_13 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1729" *) free_adr_mask[26];
  assign index_l0_14 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1730" *) free_adr_mask[28];
  assign index_l0_15 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1731" *) free_adr_mask[30];
  assign index_l0_16 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1732" *) free_adr_mask[32];
  assign index_l0_17 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1733" *) free_adr_mask[34];
  assign index_l0_18 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1734" *) free_adr_mask[36];
  assign index_l0_19 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1735" *) free_adr_mask[38];
  assign index_l0_20 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1736" *) free_adr_mask[40];
  assign index_l0_21 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1737" *) free_adr_mask[42];
  assign index_l0_22 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1738" *) free_adr_mask[44];
  assign index_l0_23 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1739" *) free_adr_mask[46];
  assign index_l0_24 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1740" *) free_adr_mask[48];
  assign index_l0_25 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1741" *) free_adr_mask[50];
  assign index_l0_26 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1742" *) free_adr_mask[52];
  assign index_l0_27 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1743" *) free_adr_mask[54];
  assign index_l0_28 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1744" *) free_adr_mask[56];
  assign index_l0_29 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1745" *) free_adr_mask[58];
  assign index_l0_30 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1746" *) free_adr_mask[60];
  assign index_l0_31 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1747" *) free_adr_mask[62];
  assign index_l0_32 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1748" *) free_adr_mask[64];
  assign index_l0_33 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1749" *) free_adr_mask[66];
  assign index_l0_34 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1750" *) free_adr_mask[68];
  assign index_l0_35 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1751" *) free_adr_mask[70];
  assign index_l0_36 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1752" *) free_adr_mask[72];
  assign index_l0_37 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1753" *) free_adr_mask[74];
  assign index_l0_38 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1754" *) free_adr_mask[76];
  assign index_l0_39 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1755" *) free_adr_mask[78];
  assign index_l0_40 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1756" *) free_adr_mask[80];
  assign index_l0_41 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1757" *) free_adr_mask[82];
  assign index_l0_42 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1758" *) free_adr_mask[84];
  assign index_l0_43 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1759" *) free_adr_mask[86];
  assign index_l0_44 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1760" *) free_adr_mask[88];
  assign index_l0_45 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1761" *) free_adr_mask[90];
  assign index_l0_46 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1762" *) free_adr_mask[92];
  assign index_l0_47 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1763" *) free_adr_mask[94];
  assign index_l0_48 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1764" *) free_adr_mask[96];
  assign index_l0_49 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1765" *) free_adr_mask[98];
  assign index_l0_50 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1766" *) free_adr_mask[100];
  assign index_l0_51 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1767" *) free_adr_mask[102];
  assign index_l0_52 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1768" *) free_adr_mask[104];
  assign index_l0_53 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1769" *) free_adr_mask[106];
  assign index_l0_54 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1770" *) free_adr_mask[108];
  assign index_l0_55 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1771" *) free_adr_mask[110];
  assign index_l0_56 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1772" *) free_adr_mask[112];
  assign index_l0_57 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1773" *) free_adr_mask[114];
  assign index_l0_58 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1774" *) free_adr_mask[116];
  assign index_l0_59 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1775" *) free_adr_mask[118];
  assign index_l0_60 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1776" *) free_adr_mask[120];
  assign index_l0_61 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1777" *) free_adr_mask[122];
  assign index_l0_62 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1778" *) free_adr_mask[124];
  assign index_l0_63 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1779" *) free_adr_mask[126];
  assign index_l0_64 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1780" *) free_adr_mask[128];
  assign index_l0_65 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1781" *) free_adr_mask[130];
  assign index_l0_66 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1782" *) free_adr_mask[132];
  assign index_l0_67 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1783" *) free_adr_mask[134];
  assign index_l0_68 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1784" *) free_adr_mask[136];
  assign index_l0_69 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1785" *) free_adr_mask[138];
  assign index_l0_70 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1786" *) free_adr_mask[140];
  assign index_l0_71 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1787" *) free_adr_mask[142];
  assign index_l0_72 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1788" *) free_adr_mask[144];
  assign index_l0_73 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1789" *) free_adr_mask[146];
  assign index_l0_74 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1790" *) free_adr_mask[148];
  assign index_l0_75 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1791" *) free_adr_mask[150];
  assign index_l0_76 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1792" *) free_adr_mask[152];
  assign index_l0_77 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1793" *) free_adr_mask[154];
  assign index_l0_78 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1794" *) free_adr_mask[156];
  assign index_l0_79 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1795" *) free_adr_mask[158];
  assign index_l0_80 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1796" *) free_adr_mask[160];
  assign index_l0_81 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1797" *) free_adr_mask[162];
  assign index_l0_82 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1798" *) free_adr_mask[164];
  assign index_l0_83 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1799" *) free_adr_mask[166];
  assign index_l0_84 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1800" *) free_adr_mask[168];
  assign index_l0_85 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1801" *) free_adr_mask[170];
  assign index_l0_86 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1802" *) free_adr_mask[172];
  assign index_l0_87 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1803" *) free_adr_mask[174];
  assign index_l0_88 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1804" *) free_adr_mask[176];
  assign index_l0_89 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1805" *) free_adr_mask[178];
  assign index_l0_90 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1806" *) free_adr_mask[180];
  assign index_l0_91 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1807" *) free_adr_mask[182];
  assign index_l0_92 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1808" *) free_adr_mask[184];
  assign index_l0_93 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1809" *) free_adr_mask[186];
  assign index_l0_94 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1810" *) free_adr_mask[188];
  assign index_l0_95 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1811" *) free_adr_mask[190];
  assign index_l0_96 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1812" *) free_adr_mask[192];
  assign index_l0_97 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1813" *) free_adr_mask[194];
  assign index_l0_98 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1814" *) free_adr_mask[196];
  assign index_l0_99 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1815" *) free_adr_mask[198];
  assign index_l0_100 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1816" *) free_adr_mask[200];
  assign index_l0_101 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1817" *) free_adr_mask[202];
  assign index_l0_102 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1818" *) free_adr_mask[204];
  assign index_l0_103 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1819" *) free_adr_mask[206];
  assign index_l0_104 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1820" *) free_adr_mask[208];
  assign index_l0_105 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1821" *) free_adr_mask[210];
  assign index_l0_106 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1822" *) free_adr_mask[212];
  assign index_l0_107 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1823" *) free_adr_mask[214];
  assign index_l0_108 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1824" *) free_adr_mask[216];
  assign index_l0_109 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1825" *) free_adr_mask[218];
  assign index_l0_110 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1826" *) free_adr_mask[220];
  assign index_l0_111 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1827" *) free_adr_mask[222];
  assign index_l0_112 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1828" *) free_adr_mask[224];
  assign index_l0_113 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1829" *) free_adr_mask[226];
  assign index_l0_114 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1830" *) free_adr_mask[228];
  assign index_l0_115 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1831" *) free_adr_mask[230];
  assign index_l0_116 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1832" *) free_adr_mask[232];
  assign index_l0_117 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1833" *) free_adr_mask[234];
  assign index_l0_118 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1834" *) free_adr_mask[236];
  assign index_l0_119 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1835" *) free_adr_mask[238];
  assign index_l0_120 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1836" *) free_adr_mask[240];
  assign index_l0_121 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1837" *) free_adr_mask[242];
  assign index_l0_122 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1838" *) free_adr_mask[244];
  assign index_l0_123 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1839" *) free_adr_mask[246];
  assign index_l0_124 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1840" *) free_adr_mask[248];
  assign index_l0_125 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1841" *) free_adr_mask[250];
  assign index_l0_126 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1842" *) free_adr_mask[252];
  assign index_l0_127 = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1843" *) free_adr_mask[254];
  assign index_l1_0[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1844" *) flag_l0_0;
  assign index_l1_1[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1845" *) flag_l0_2;
  assign index_l1_2[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1846" *) flag_l0_4;
  assign index_l1_3[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1847" *) flag_l0_6;
  assign index_l1_4[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1848" *) flag_l0_8;
  assign index_l1_5[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1849" *) flag_l0_10;
  assign index_l1_6[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1850" *) flag_l0_12;
  assign index_l1_7[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1851" *) flag_l0_14;
  assign index_l1_8[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1852" *) flag_l0_16;
  assign index_l1_9[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1853" *) flag_l0_18;
  assign index_l1_10[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1854" *) flag_l0_20;
  assign index_l1_11[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1855" *) flag_l0_22;
  assign index_l1_12[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1856" *) flag_l0_24;
  assign index_l1_13[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1857" *) flag_l0_26;
  assign index_l1_14[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1858" *) flag_l0_28;
  assign index_l1_15[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1859" *) flag_l0_30;
  assign index_l1_16[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1860" *) flag_l0_32;
  assign index_l1_17[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1861" *) flag_l0_34;
  assign index_l1_18[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1862" *) flag_l0_36;
  assign index_l1_19[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1863" *) flag_l0_38;
  assign index_l1_20[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1864" *) flag_l0_40;
  assign index_l1_21[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1865" *) flag_l0_42;
  assign index_l1_22[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1866" *) flag_l0_44;
  assign index_l1_23[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1867" *) flag_l0_46;
  assign index_l1_24[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1868" *) flag_l0_48;
  assign index_l1_25[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1869" *) flag_l0_50;
  assign index_l1_26[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1870" *) flag_l0_52;
  assign index_l1_27[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1871" *) flag_l0_54;
  assign index_l1_28[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1872" *) flag_l0_56;
  assign index_l1_29[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1873" *) flag_l0_58;
  assign index_l1_30[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1874" *) flag_l0_60;
  assign index_l1_31[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1875" *) flag_l0_62;
  assign index_l1_32[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1876" *) flag_l0_64;
  assign index_l1_33[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1877" *) flag_l0_66;
  assign index_l1_34[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1878" *) flag_l0_68;
  assign index_l1_35[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1879" *) flag_l0_70;
  assign index_l1_36[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1880" *) flag_l0_72;
  assign index_l1_37[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1881" *) flag_l0_74;
  assign index_l1_38[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1882" *) flag_l0_76;
  assign index_l1_39[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1883" *) flag_l0_78;
  assign index_l1_40[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1884" *) flag_l0_80;
  assign index_l1_41[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1885" *) flag_l0_82;
  assign index_l1_42[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1886" *) flag_l0_84;
  assign index_l1_43[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1887" *) flag_l0_86;
  assign index_l1_44[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1888" *) flag_l0_88;
  assign index_l1_45[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1889" *) flag_l0_90;
  assign index_l1_46[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1890" *) flag_l0_92;
  assign index_l1_47[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1891" *) flag_l0_94;
  assign index_l1_48[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1892" *) flag_l0_96;
  assign index_l1_49[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1893" *) flag_l0_98;
  assign index_l1_50[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1894" *) flag_l0_100;
  assign index_l1_51[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1895" *) flag_l0_102;
  assign index_l1_52[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1896" *) flag_l0_104;
  assign index_l1_53[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1897" *) flag_l0_106;
  assign index_l1_54[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1898" *) flag_l0_108;
  assign index_l1_55[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1899" *) flag_l0_110;
  assign index_l1_56[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1900" *) flag_l0_112;
  assign index_l1_57[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1901" *) flag_l0_114;
  assign index_l1_58[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1902" *) flag_l0_116;
  assign index_l1_59[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1903" *) flag_l0_118;
  assign index_l1_60[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1904" *) flag_l0_120;
  assign index_l1_61[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1905" *) flag_l0_122;
  assign index_l1_62[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1906" *) flag_l0_124;
  assign index_l1_63[1] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1907" *) flag_l0_126;
  assign index_l2_0[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1908" *) flag_l1_0;
  assign index_l2_1[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1909" *) flag_l1_2;
  assign index_l2_2[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1910" *) flag_l1_4;
  assign index_l2_3[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1911" *) flag_l1_6;
  assign index_l2_4[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1912" *) flag_l1_8;
  assign index_l2_5[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1913" *) flag_l1_10;
  assign index_l2_6[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1914" *) flag_l1_12;
  assign index_l2_7[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1915" *) flag_l1_14;
  assign index_l2_8[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1916" *) flag_l1_16;
  assign index_l2_9[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1917" *) flag_l1_18;
  assign index_l2_10[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1918" *) flag_l1_20;
  assign index_l2_11[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1919" *) flag_l1_22;
  assign index_l2_12[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1920" *) flag_l1_24;
  assign index_l2_13[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1921" *) flag_l1_26;
  assign index_l2_14[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1922" *) flag_l1_28;
  assign index_l2_15[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1923" *) flag_l1_30;
  assign index_l2_16[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1924" *) flag_l1_32;
  assign index_l2_17[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1925" *) flag_l1_34;
  assign index_l2_18[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1926" *) flag_l1_36;
  assign index_l2_19[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1927" *) flag_l1_38;
  assign index_l2_20[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1928" *) flag_l1_40;
  assign index_l2_21[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1929" *) flag_l1_42;
  assign index_l2_22[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1930" *) flag_l1_44;
  assign index_l2_23[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1931" *) flag_l1_46;
  assign index_l2_24[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1932" *) flag_l1_48;
  assign index_l2_25[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1933" *) flag_l1_50;
  assign index_l2_26[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1934" *) flag_l1_52;
  assign index_l2_27[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1935" *) flag_l1_54;
  assign index_l2_28[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1936" *) flag_l1_56;
  assign index_l2_29[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1937" *) flag_l1_58;
  assign index_l2_30[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1938" *) flag_l1_60;
  assign index_l2_31[2] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1939" *) flag_l1_62;
  assign index_l3_0[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1940" *) flag_l2_0;
  assign index_l3_1[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1941" *) flag_l2_2;
  assign index_l3_2[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1942" *) flag_l2_4;
  assign index_l3_3[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1943" *) flag_l2_6;
  assign index_l3_4[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1944" *) flag_l2_8;
  assign index_l3_5[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1945" *) flag_l2_10;
  assign index_l3_6[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1946" *) flag_l2_12;
  assign index_l3_7[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1947" *) flag_l2_14;
  assign index_l3_8[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1948" *) flag_l2_16;
  assign index_l3_9[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1949" *) flag_l2_18;
  assign index_l3_10[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1950" *) flag_l2_20;
  assign index_l3_11[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1951" *) flag_l2_22;
  assign index_l3_12[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1952" *) flag_l2_24;
  assign index_l3_13[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1953" *) flag_l2_26;
  assign index_l3_14[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1954" *) flag_l2_28;
  assign index_l3_15[3] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1955" *) flag_l2_30;
  assign index_l4_0[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1956" *) flag_l3_0;
  assign index_l4_1[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1957" *) flag_l3_2;
  assign index_l4_2[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1958" *) flag_l3_4;
  assign index_l4_3[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1959" *) flag_l3_6;
  assign index_l4_4[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1960" *) flag_l3_8;
  assign index_l4_5[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1961" *) flag_l3_10;
  assign index_l4_6[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1962" *) flag_l3_12;
  assign index_l4_7[4] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1963" *) flag_l3_14;
  assign index_l5_0[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1964" *) flag_l4_0;
  assign index_l5_1[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1965" *) flag_l4_2;
  assign index_l5_2[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1966" *) flag_l4_4;
  assign index_l5_3[5] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1967" *) flag_l4_6;
  assign index_l6_0[6] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1968" *) flag_l5_0;
  assign index_l6_1[6] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1969" *) flag_l5_2;
  assign adr_ram_wr_data[7] = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1970" *) flag_l6_0;
  assign _1550_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) rd_skid0_0_vld;
  assign _1551_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) rd_skid0_1_vld;
  assign _1552_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *) rd_skid0_2_vld;
  assign _1553_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *) _1103_;
  assign _1554_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) rd_take_n_dly[0];
  assign cq_wr_prdy = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) cq_wr_busy_int;
  assign _1555_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) cq_rd_credit[0];
  assign _1556_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) cq_rd0_prdy_d;
  assign _1557_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) _1123_;
  assign _1558_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) rd_skid1_0_vld;
  assign _1559_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) rd_skid1_1_vld;
  assign _1560_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *) rd_skid1_2_vld;
  assign _1561_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *) _1127_;
  assign _1562_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) rd_take_n_dly[1];
  assign _1563_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) cq_rd_credit[1];
  assign _1564_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) cq_rd1_prdy_d;
  assign _1565_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) _1147_;
  assign _1566_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) rd_skid2_0_vld;
  assign _1567_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) rd_skid2_1_vld;
  assign _1568_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *) rd_skid2_2_vld;
  assign _1569_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *) _1150_;
  assign _1570_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) rd_take_n_dly[2];
  assign _1571_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) cq_rd_credit[2];
  assign _1572_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) cq_rd2_prdy_d;
  assign _1573_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) _1171_;
  assign _1574_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) rd_skid3_0_vld;
  assign _1575_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) rd_skid3_1_vld;
  assign _1576_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *) rd_skid3_2_vld;
  assign _1577_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *) _1174_;
  assign _1578_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) rd_take_n_dly[3];
  assign _1579_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) cq_rd_credit[3];
  assign _1580_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) cq_rd3_prdy_d;
  assign _1581_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) _1195_;
  assign _1582_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) rd_skid4_0_vld;
  assign _1583_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) rd_skid4_1_vld;
  assign _1584_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *) rd_skid4_2_vld;
  assign _1585_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *) _1198_;
  assign _1586_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) rd_take_n_dly[4];
  assign _1587_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) cq_rd_credit[4];
  assign _1588_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) cq_rd4_prdy_d;
  assign _1589_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) _1218_;
  assign _1590_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2802" *) cq_rd_take_elig[0];
  assign _1591_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2803" *) cq_rd_take_elig[4];
  assign _1592_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2804" *) cq_rd_take_elig[3];
  assign _1593_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2805" *) cq_rd_take_elig[2];
  assign _1594_ = ! (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2808" *) cq_rd_take_elig[1];
  assign _1595_ = rd_take_dly || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:180" *) rd_pushing;
  assign _1596_ = rd_pushing || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing_q;
  assign update_rd_take_n_dly = cq_rd_take || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2016" *) rd_take_dly;
  assign _1597_ = rd_pushing || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2131" *) cq_rd_take;
  assign _1598_ = _1066_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *) _1068_;
  assign _1599_ = _1069_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *) _1071_;
  assign _1600_ = _1073_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *) _1075_;
  assign _1601_ = _1076_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *) _1078_;
  assign _1602_ = _1080_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *) _1082_;
  assign cq_rd0_pvld = rd_skid0_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2334" *) rd_pre_bypassing0;
  assign _1603_ = rd_bypassing0 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) rd_take_n_dly[0];
  assign _1604_ = _1550_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) _1104_;
  assign _1605_ = _1551_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *) _1107_;
  assign _1606_ = rd_skid0_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *) _1553_;
  assign _1607_ = rd_skid0_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *) _1114_;
  assign _1608_ = _1607_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *) rd_take_n_dly[0];
  assign _1609_ = rd_skid0_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *) rd_bypassing0;
  assign _1610_ = _1609_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *) rd_take_n_dly[0];
  assign _1611_ = rd_skid0_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *) _1115_;
  assign _1612_ = rd_skid0_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *) _1111_;
  assign _1613_ = cq_rd0_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) _1550_;
  assign _1614_ = _1613_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) _1551_;
  assign _1615_ = _1614_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) _1118_;
  assign _1616_ = cq_rd_credit[0] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2392" *) cq_rd0_credits_ne0;
  assign _1617_ = _1554_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2394" *) rd_skid0_0_vld;
  assign _1618_ = _1552_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) _1551_;
  assign _1619_ = _1618_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2395" *) _1557_;
  assign cq_rd1_pvld = rd_skid1_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2430" *) rd_pre_bypassing1;
  assign _1620_ = rd_bypassing1 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) rd_take_n_dly[1];
  assign _1621_ = _1558_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) _1128_;
  assign _1622_ = _1559_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *) _1131_;
  assign _1623_ = rd_skid1_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *) _1561_;
  assign _1624_ = rd_skid1_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *) _1138_;
  assign _1625_ = _1624_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *) rd_take_n_dly[1];
  assign _1626_ = rd_skid1_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *) rd_bypassing1;
  assign _1627_ = _1626_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *) rd_take_n_dly[1];
  assign _1628_ = rd_skid1_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *) _1139_;
  assign _1629_ = rd_skid1_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *) _1135_;
  assign _1630_ = cq_rd1_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) _1558_;
  assign _1631_ = _1630_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) _1559_;
  assign _1632_ = _1631_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) _1142_;
  assign _1633_ = cq_rd_credit[1] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2488" *) cq_rd1_credits_ne0;
  assign _1634_ = _1562_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2490" *) rd_skid1_0_vld;
  assign _1635_ = _1560_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) _1559_;
  assign _1636_ = _1635_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2491" *) _1565_;
  assign cq_rd2_pvld = rd_skid2_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2526" *) rd_pre_bypassing2;
  assign _1637_ = rd_bypassing2 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) rd_take_n_dly[2];
  assign _1638_ = _1566_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) _1151_;
  assign _1639_ = _1567_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *) _1155_;
  assign _1640_ = rd_skid2_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *) _1569_;
  assign _1641_ = rd_skid2_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *) _1162_;
  assign _1642_ = _1641_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *) rd_take_n_dly[2];
  assign _1643_ = rd_skid2_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *) rd_bypassing2;
  assign _1644_ = _1643_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *) rd_take_n_dly[2];
  assign _1645_ = rd_skid2_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *) _1163_;
  assign _1646_ = rd_skid2_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *) _1159_;
  assign _1647_ = cq_rd2_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) _1566_;
  assign _1648_ = _1647_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) _1567_;
  assign _1649_ = _1648_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) _1166_;
  assign _1650_ = cq_rd_credit[2] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2584" *) cq_rd2_credits_ne0;
  assign _1651_ = _1570_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2586" *) rd_skid2_0_vld;
  assign _1652_ = _1568_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) _1567_;
  assign _1653_ = _1652_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2587" *) _1573_;
  assign cq_rd3_pvld = rd_skid3_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2622" *) rd_pre_bypassing3;
  assign _1654_ = rd_bypassing3 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) rd_take_n_dly[3];
  assign _1655_ = _1574_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) _1175_;
  assign _1656_ = _1575_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *) _1179_;
  assign _1657_ = rd_skid3_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *) _1577_;
  assign _1658_ = rd_skid3_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *) _1186_;
  assign _1659_ = _1658_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *) rd_take_n_dly[3];
  assign _1660_ = rd_skid3_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *) rd_bypassing3;
  assign _1661_ = _1660_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *) rd_take_n_dly[3];
  assign _1662_ = rd_skid3_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *) _1187_;
  assign _1663_ = rd_skid3_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *) _1182_;
  assign _1664_ = cq_rd3_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) _1574_;
  assign _1665_ = _1664_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) _1575_;
  assign _1666_ = _1665_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) _1190_;
  assign _1667_ = cq_rd_credit[3] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2680" *) cq_rd3_credits_ne0;
  assign _1668_ = _1578_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2682" *) rd_skid3_0_vld;
  assign _1669_ = _1576_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) _1575_;
  assign _1670_ = _1669_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2683" *) _1581_;
  assign cq_rd4_pvld = rd_skid4_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2718" *) rd_pre_bypassing4;
  assign _1671_ = rd_bypassing4 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) rd_take_n_dly[4];
  assign _1672_ = _1582_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) _1199_;
  assign _1673_ = _1583_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *) _1203_;
  assign _1674_ = rd_skid4_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *) _1585_;
  assign _1675_ = rd_skid4_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *) _1210_;
  assign _1676_ = _1675_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *) rd_take_n_dly[4];
  assign _1677_ = rd_skid4_0_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *) rd_bypassing4;
  assign _1678_ = _1677_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *) rd_take_n_dly[4];
  assign _1679_ = rd_skid4_2_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *) _1211_;
  assign _1680_ = rd_skid4_1_vld || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *) _1206_;
  assign _1681_ = cq_rd4_prdy_d || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) _1582_;
  assign _1682_ = _1681_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) _1583_;
  assign _1683_ = _1682_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) _1213_;
  assign _1684_ = cq_rd_credit[4] || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2776" *) cq_rd4_credits_ne0;
  assign _1685_ = _1586_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2778" *) rd_skid4_0_vld;
  assign _1686_ = _1584_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) _1583_;
  assign _1687_ = _1686_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2779" *) _1589_;
  assign _1688_ = rd_bypassing0 || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *) rd_bypassing1;
  assign _1689_ = _1688_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *) rd_bypassing2;
  assign _1690_ = _1689_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *) rd_bypassing3;
  assign wr_bypassing = _1690_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2843" *) rd_bypassing4;
  assign _1691_ = wr_reserving || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) rd_pushing;
  assign _1692_ = _1691_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) rd_take_dly;
  assign _1693_ = _1692_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) wr_reserving;
  assign _1694_ = _1693_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) _1722_;
  assign _1695_ = _1694_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) rd_take_dly;
  assign _1696_ = _1597_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) _1723_;
  assign _1697_ = _1696_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) rd_take_dly;
  assign nvdla_core_clk_mgated_enable = _1695_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) _1697_;
  assign _1698_ = nvdla_core_clk_mgated_enable || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) _1103_;
  assign _1699_ = _1698_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) rd_bypassing0;
  assign _1700_ = _1699_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) _1127_;
  assign _1701_ = _1700_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) rd_bypassing1;
  assign _1702_ = _1701_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) _1150_;
  assign _1703_ = _1702_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) rd_bypassing2;
  assign _1704_ = _1703_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) _1174_;
  assign _1705_ = _1704_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) rd_bypassing3;
  assign _1706_ = _1705_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2878" *) _1198_;
  assign nvdla_core_clk_mgated_skid_enable = _1706_ || (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2889" *) rd_bypassing4;
  assign _1707_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2244" *) cq_rd_count0;
  assign _1708_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2245" *) cq_rd_count1;
  assign _1709_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2246" *) cq_rd_count2;
  assign _1710_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2247" *) cq_rd_count3;
  assign _1711_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2248" *) cq_rd_count4;
  assign _1712_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2403" *) cq_rd0_credits_w_take_next;
  assign _1713_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2403" *) cq_rd0_credits_wo_take_next;
  assign _1714_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2499" *) cq_rd1_credits_w_take_next;
  assign _1715_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2499" *) cq_rd1_credits_wo_take_next;
  assign _1716_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2595" *) cq_rd2_credits_w_take_next;
  assign _1717_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2595" *) cq_rd2_credits_wo_take_next;
  assign _1718_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2691" *) cq_rd3_credits_w_take_next;
  assign _1719_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2691" *) cq_rd3_credits_wo_take_next;
  assign _1720_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2787" *) cq_rd4_credits_w_take_next;
  assign _1721_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2787" *) cq_rd4_credits_wo_take_next;
  assign _1722_ = cq_wr_busy_int != (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) cq_wr_busy_next;
  assign _1723_ = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2866" *) cq_rd_credit;
  assign flag_l0_0 = free_adr_mask[1] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1469" *) free_adr_mask[0];
  assign flag_l0_1 = free_adr_mask[3] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1470" *) free_adr_mask[2];
  assign flag_l0_2 = free_adr_mask[5] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1471" *) free_adr_mask[4];
  assign flag_l0_3 = free_adr_mask[7] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1472" *) free_adr_mask[6];
  assign flag_l0_4 = free_adr_mask[9] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1473" *) free_adr_mask[8];
  assign flag_l0_5 = free_adr_mask[11] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1474" *) free_adr_mask[10];
  assign flag_l0_6 = free_adr_mask[13] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1475" *) free_adr_mask[12];
  assign flag_l0_7 = free_adr_mask[15] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1476" *) free_adr_mask[14];
  assign flag_l0_8 = free_adr_mask[17] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1477" *) free_adr_mask[16];
  assign flag_l0_9 = free_adr_mask[19] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1478" *) free_adr_mask[18];
  assign flag_l0_10 = free_adr_mask[21] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1479" *) free_adr_mask[20];
  assign flag_l0_11 = free_adr_mask[23] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1480" *) free_adr_mask[22];
  assign flag_l0_12 = free_adr_mask[25] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1481" *) free_adr_mask[24];
  assign flag_l0_13 = free_adr_mask[27] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1482" *) free_adr_mask[26];
  assign flag_l0_14 = free_adr_mask[29] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1483" *) free_adr_mask[28];
  assign flag_l0_15 = free_adr_mask[31] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1484" *) free_adr_mask[30];
  assign flag_l0_16 = free_adr_mask[33] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1485" *) free_adr_mask[32];
  assign flag_l0_17 = free_adr_mask[35] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1486" *) free_adr_mask[34];
  assign flag_l0_18 = free_adr_mask[37] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1487" *) free_adr_mask[36];
  assign flag_l0_19 = free_adr_mask[39] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1488" *) free_adr_mask[38];
  assign flag_l0_20 = free_adr_mask[41] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1489" *) free_adr_mask[40];
  assign flag_l0_21 = free_adr_mask[43] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1490" *) free_adr_mask[42];
  assign flag_l0_22 = free_adr_mask[45] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1491" *) free_adr_mask[44];
  assign flag_l0_23 = free_adr_mask[47] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1492" *) free_adr_mask[46];
  assign flag_l0_24 = free_adr_mask[49] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1493" *) free_adr_mask[48];
  assign flag_l0_25 = free_adr_mask[51] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1494" *) free_adr_mask[50];
  assign flag_l0_26 = free_adr_mask[53] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1495" *) free_adr_mask[52];
  assign flag_l0_27 = free_adr_mask[55] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1496" *) free_adr_mask[54];
  assign flag_l0_28 = free_adr_mask[57] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1497" *) free_adr_mask[56];
  assign flag_l0_29 = free_adr_mask[59] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1498" *) free_adr_mask[58];
  assign flag_l0_30 = free_adr_mask[61] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1499" *) free_adr_mask[60];
  assign flag_l0_31 = free_adr_mask[63] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1500" *) free_adr_mask[62];
  assign flag_l0_32 = free_adr_mask[65] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1501" *) free_adr_mask[64];
  assign flag_l0_33 = free_adr_mask[67] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1502" *) free_adr_mask[66];
  assign flag_l0_34 = free_adr_mask[69] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1503" *) free_adr_mask[68];
  assign flag_l0_35 = free_adr_mask[71] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1504" *) free_adr_mask[70];
  assign flag_l0_36 = free_adr_mask[73] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1505" *) free_adr_mask[72];
  assign flag_l0_37 = free_adr_mask[75] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1506" *) free_adr_mask[74];
  assign flag_l0_38 = free_adr_mask[77] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1507" *) free_adr_mask[76];
  assign flag_l0_39 = free_adr_mask[79] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1508" *) free_adr_mask[78];
  assign flag_l0_40 = free_adr_mask[81] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1509" *) free_adr_mask[80];
  assign flag_l0_41 = free_adr_mask[83] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1510" *) free_adr_mask[82];
  assign flag_l0_42 = free_adr_mask[85] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1511" *) free_adr_mask[84];
  assign flag_l0_43 = free_adr_mask[87] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1512" *) free_adr_mask[86];
  assign flag_l0_44 = free_adr_mask[89] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1513" *) free_adr_mask[88];
  assign flag_l0_45 = free_adr_mask[91] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1514" *) free_adr_mask[90];
  assign flag_l0_46 = free_adr_mask[93] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1515" *) free_adr_mask[92];
  assign flag_l0_47 = free_adr_mask[95] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1516" *) free_adr_mask[94];
  assign flag_l0_48 = free_adr_mask[97] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1517" *) free_adr_mask[96];
  assign flag_l0_49 = free_adr_mask[99] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1518" *) free_adr_mask[98];
  assign flag_l0_50 = free_adr_mask[101] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1519" *) free_adr_mask[100];
  assign flag_l0_51 = free_adr_mask[103] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1520" *) free_adr_mask[102];
  assign flag_l0_52 = free_adr_mask[105] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1521" *) free_adr_mask[104];
  assign flag_l0_53 = free_adr_mask[107] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1522" *) free_adr_mask[106];
  assign flag_l0_54 = free_adr_mask[109] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1523" *) free_adr_mask[108];
  assign flag_l0_55 = free_adr_mask[111] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1524" *) free_adr_mask[110];
  assign flag_l0_56 = free_adr_mask[113] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1525" *) free_adr_mask[112];
  assign flag_l0_57 = free_adr_mask[115] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1526" *) free_adr_mask[114];
  assign flag_l0_58 = free_adr_mask[117] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1527" *) free_adr_mask[116];
  assign flag_l0_59 = free_adr_mask[119] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1528" *) free_adr_mask[118];
  assign flag_l0_60 = free_adr_mask[121] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1529" *) free_adr_mask[120];
  assign flag_l0_61 = free_adr_mask[123] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1530" *) free_adr_mask[122];
  assign flag_l0_62 = free_adr_mask[125] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1531" *) free_adr_mask[124];
  assign flag_l0_63 = free_adr_mask[127] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1532" *) free_adr_mask[126];
  assign flag_l0_64 = free_adr_mask[129] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1533" *) free_adr_mask[128];
  assign flag_l0_65 = free_adr_mask[131] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1534" *) free_adr_mask[130];
  assign flag_l0_66 = free_adr_mask[133] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1535" *) free_adr_mask[132];
  assign flag_l0_67 = free_adr_mask[135] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1536" *) free_adr_mask[134];
  assign flag_l0_68 = free_adr_mask[137] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1537" *) free_adr_mask[136];
  assign flag_l0_69 = free_adr_mask[139] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1538" *) free_adr_mask[138];
  assign flag_l0_70 = free_adr_mask[141] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1539" *) free_adr_mask[140];
  assign flag_l0_71 = free_adr_mask[143] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1540" *) free_adr_mask[142];
  assign flag_l0_72 = free_adr_mask[145] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1541" *) free_adr_mask[144];
  assign flag_l0_73 = free_adr_mask[147] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1542" *) free_adr_mask[146];
  assign flag_l0_74 = free_adr_mask[149] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1543" *) free_adr_mask[148];
  assign flag_l0_75 = free_adr_mask[151] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1544" *) free_adr_mask[150];
  assign flag_l0_76 = free_adr_mask[153] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1545" *) free_adr_mask[152];
  assign flag_l0_77 = free_adr_mask[155] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1546" *) free_adr_mask[154];
  assign flag_l0_78 = free_adr_mask[157] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1547" *) free_adr_mask[156];
  assign flag_l0_79 = free_adr_mask[159] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1548" *) free_adr_mask[158];
  assign flag_l0_80 = free_adr_mask[161] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1549" *) free_adr_mask[160];
  assign flag_l0_81 = free_adr_mask[163] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1550" *) free_adr_mask[162];
  assign flag_l0_82 = free_adr_mask[165] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1551" *) free_adr_mask[164];
  assign flag_l0_83 = free_adr_mask[167] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1552" *) free_adr_mask[166];
  assign flag_l0_84 = free_adr_mask[169] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1553" *) free_adr_mask[168];
  assign flag_l0_85 = free_adr_mask[171] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1554" *) free_adr_mask[170];
  assign flag_l0_86 = free_adr_mask[173] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1555" *) free_adr_mask[172];
  assign flag_l0_87 = free_adr_mask[175] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1556" *) free_adr_mask[174];
  assign flag_l0_88 = free_adr_mask[177] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1557" *) free_adr_mask[176];
  assign flag_l0_89 = free_adr_mask[179] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1558" *) free_adr_mask[178];
  assign flag_l0_90 = free_adr_mask[181] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1559" *) free_adr_mask[180];
  assign flag_l0_91 = free_adr_mask[183] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1560" *) free_adr_mask[182];
  assign flag_l0_92 = free_adr_mask[185] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1561" *) free_adr_mask[184];
  assign flag_l0_93 = free_adr_mask[187] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1562" *) free_adr_mask[186];
  assign flag_l0_94 = free_adr_mask[189] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1563" *) free_adr_mask[188];
  assign flag_l0_95 = free_adr_mask[191] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1564" *) free_adr_mask[190];
  assign flag_l0_96 = free_adr_mask[193] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1565" *) free_adr_mask[192];
  assign flag_l0_97 = free_adr_mask[195] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1566" *) free_adr_mask[194];
  assign flag_l0_98 = free_adr_mask[197] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1567" *) free_adr_mask[196];
  assign flag_l0_99 = free_adr_mask[199] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1568" *) free_adr_mask[198];
  assign flag_l0_100 = free_adr_mask[201] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1569" *) free_adr_mask[200];
  assign flag_l0_101 = free_adr_mask[203] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1570" *) free_adr_mask[202];
  assign flag_l0_102 = free_adr_mask[205] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1571" *) free_adr_mask[204];
  assign flag_l0_103 = free_adr_mask[207] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1572" *) free_adr_mask[206];
  assign flag_l0_104 = free_adr_mask[209] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1573" *) free_adr_mask[208];
  assign flag_l0_105 = free_adr_mask[211] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1574" *) free_adr_mask[210];
  assign flag_l0_106 = free_adr_mask[213] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1575" *) free_adr_mask[212];
  assign flag_l0_107 = free_adr_mask[215] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1576" *) free_adr_mask[214];
  assign flag_l0_108 = free_adr_mask[217] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1577" *) free_adr_mask[216];
  assign flag_l0_109 = free_adr_mask[219] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1578" *) free_adr_mask[218];
  assign flag_l0_110 = free_adr_mask[221] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1579" *) free_adr_mask[220];
  assign flag_l0_111 = free_adr_mask[223] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1580" *) free_adr_mask[222];
  assign flag_l0_112 = free_adr_mask[225] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1581" *) free_adr_mask[224];
  assign flag_l0_113 = free_adr_mask[227] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1582" *) free_adr_mask[226];
  assign flag_l0_114 = free_adr_mask[229] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1583" *) free_adr_mask[228];
  assign flag_l0_115 = free_adr_mask[231] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1584" *) free_adr_mask[230];
  assign flag_l0_116 = free_adr_mask[233] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1585" *) free_adr_mask[232];
  assign flag_l0_117 = free_adr_mask[235] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1586" *) free_adr_mask[234];
  assign flag_l0_118 = free_adr_mask[237] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1587" *) free_adr_mask[236];
  assign flag_l0_119 = free_adr_mask[239] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1588" *) free_adr_mask[238];
  assign flag_l0_120 = free_adr_mask[241] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1589" *) free_adr_mask[240];
  assign flag_l0_121 = free_adr_mask[243] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1590" *) free_adr_mask[242];
  assign flag_l0_122 = free_adr_mask[245] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1591" *) free_adr_mask[244];
  assign flag_l0_123 = free_adr_mask[247] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1592" *) free_adr_mask[246];
  assign flag_l0_124 = free_adr_mask[249] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1593" *) free_adr_mask[248];
  assign flag_l0_125 = free_adr_mask[251] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1594" *) free_adr_mask[250];
  assign flag_l0_126 = free_adr_mask[253] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1595" *) free_adr_mask[252];
  assign flag_l1_0 = flag_l0_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1596" *) flag_l0_0;
  assign flag_l1_1 = flag_l0_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1597" *) flag_l0_2;
  assign flag_l1_2 = flag_l0_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1598" *) flag_l0_4;
  assign flag_l1_3 = flag_l0_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1599" *) flag_l0_6;
  assign flag_l1_4 = flag_l0_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1600" *) flag_l0_8;
  assign flag_l1_5 = flag_l0_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1601" *) flag_l0_10;
  assign flag_l1_6 = flag_l0_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1602" *) flag_l0_12;
  assign flag_l1_7 = flag_l0_15 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1603" *) flag_l0_14;
  assign flag_l1_8 = flag_l0_17 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1604" *) flag_l0_16;
  assign flag_l1_9 = flag_l0_19 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1605" *) flag_l0_18;
  assign flag_l1_10 = flag_l0_21 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1606" *) flag_l0_20;
  assign flag_l1_11 = flag_l0_23 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1607" *) flag_l0_22;
  assign flag_l1_12 = flag_l0_25 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1608" *) flag_l0_24;
  assign flag_l1_13 = flag_l0_27 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1609" *) flag_l0_26;
  assign flag_l1_14 = flag_l0_29 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1610" *) flag_l0_28;
  assign flag_l1_15 = flag_l0_31 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1611" *) flag_l0_30;
  assign flag_l1_16 = flag_l0_33 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1612" *) flag_l0_32;
  assign flag_l1_17 = flag_l0_35 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1613" *) flag_l0_34;
  assign flag_l1_18 = flag_l0_37 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1614" *) flag_l0_36;
  assign flag_l1_19 = flag_l0_39 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1615" *) flag_l0_38;
  assign flag_l1_20 = flag_l0_41 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1616" *) flag_l0_40;
  assign flag_l1_21 = flag_l0_43 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1617" *) flag_l0_42;
  assign flag_l1_22 = flag_l0_45 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1618" *) flag_l0_44;
  assign flag_l1_23 = flag_l0_47 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1619" *) flag_l0_46;
  assign flag_l1_24 = flag_l0_49 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1620" *) flag_l0_48;
  assign flag_l1_25 = flag_l0_51 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1621" *) flag_l0_50;
  assign flag_l1_26 = flag_l0_53 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1622" *) flag_l0_52;
  assign flag_l1_27 = flag_l0_55 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1623" *) flag_l0_54;
  assign flag_l1_28 = flag_l0_57 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1624" *) flag_l0_56;
  assign flag_l1_29 = flag_l0_59 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1625" *) flag_l0_58;
  assign flag_l1_30 = flag_l0_61 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1626" *) flag_l0_60;
  assign flag_l1_31 = flag_l0_63 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1627" *) flag_l0_62;
  assign flag_l1_32 = flag_l0_65 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1628" *) flag_l0_64;
  assign flag_l1_33 = flag_l0_67 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1629" *) flag_l0_66;
  assign flag_l1_34 = flag_l0_69 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1630" *) flag_l0_68;
  assign flag_l1_35 = flag_l0_71 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1631" *) flag_l0_70;
  assign flag_l1_36 = flag_l0_73 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1632" *) flag_l0_72;
  assign flag_l1_37 = flag_l0_75 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1633" *) flag_l0_74;
  assign flag_l1_38 = flag_l0_77 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1634" *) flag_l0_76;
  assign flag_l1_39 = flag_l0_79 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1635" *) flag_l0_78;
  assign flag_l1_40 = flag_l0_81 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1636" *) flag_l0_80;
  assign flag_l1_41 = flag_l0_83 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1637" *) flag_l0_82;
  assign flag_l1_42 = flag_l0_85 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1638" *) flag_l0_84;
  assign flag_l1_43 = flag_l0_87 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1639" *) flag_l0_86;
  assign flag_l1_44 = flag_l0_89 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1640" *) flag_l0_88;
  assign flag_l1_45 = flag_l0_91 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1641" *) flag_l0_90;
  assign flag_l1_46 = flag_l0_93 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1642" *) flag_l0_92;
  assign flag_l1_47 = flag_l0_95 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1643" *) flag_l0_94;
  assign flag_l1_48 = flag_l0_97 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1644" *) flag_l0_96;
  assign flag_l1_49 = flag_l0_99 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1645" *) flag_l0_98;
  assign flag_l1_50 = flag_l0_101 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1646" *) flag_l0_100;
  assign flag_l1_51 = flag_l0_103 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1647" *) flag_l0_102;
  assign flag_l1_52 = flag_l0_105 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1648" *) flag_l0_104;
  assign flag_l1_53 = flag_l0_107 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1649" *) flag_l0_106;
  assign flag_l1_54 = flag_l0_109 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1650" *) flag_l0_108;
  assign flag_l1_55 = flag_l0_111 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1651" *) flag_l0_110;
  assign flag_l1_56 = flag_l0_113 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1652" *) flag_l0_112;
  assign flag_l1_57 = flag_l0_115 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1653" *) flag_l0_114;
  assign flag_l1_58 = flag_l0_117 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1654" *) flag_l0_116;
  assign flag_l1_59 = flag_l0_119 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1655" *) flag_l0_118;
  assign flag_l1_60 = flag_l0_121 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1656" *) flag_l0_120;
  assign flag_l1_61 = flag_l0_123 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1657" *) flag_l0_122;
  assign flag_l1_62 = flag_l0_125 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1658" *) flag_l0_124;
  assign flag_l2_0 = flag_l1_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1659" *) flag_l1_0;
  assign flag_l2_1 = flag_l1_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1660" *) flag_l1_2;
  assign flag_l2_2 = flag_l1_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1661" *) flag_l1_4;
  assign flag_l2_3 = flag_l1_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1662" *) flag_l1_6;
  assign flag_l2_4 = flag_l1_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1663" *) flag_l1_8;
  assign flag_l2_5 = flag_l1_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1664" *) flag_l1_10;
  assign flag_l2_6 = flag_l1_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1665" *) flag_l1_12;
  assign flag_l2_7 = flag_l1_15 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1666" *) flag_l1_14;
  assign flag_l2_8 = flag_l1_17 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1667" *) flag_l1_16;
  assign flag_l2_9 = flag_l1_19 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1668" *) flag_l1_18;
  assign flag_l2_10 = flag_l1_21 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1669" *) flag_l1_20;
  assign flag_l2_11 = flag_l1_23 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1670" *) flag_l1_22;
  assign flag_l2_12 = flag_l1_25 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1671" *) flag_l1_24;
  assign flag_l2_13 = flag_l1_27 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1672" *) flag_l1_26;
  assign flag_l2_14 = flag_l1_29 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1673" *) flag_l1_28;
  assign flag_l2_15 = flag_l1_31 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1674" *) flag_l1_30;
  assign flag_l2_16 = flag_l1_33 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1675" *) flag_l1_32;
  assign flag_l2_17 = flag_l1_35 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1676" *) flag_l1_34;
  assign flag_l2_18 = flag_l1_37 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1677" *) flag_l1_36;
  assign flag_l2_19 = flag_l1_39 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1678" *) flag_l1_38;
  assign flag_l2_20 = flag_l1_41 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1679" *) flag_l1_40;
  assign flag_l2_21 = flag_l1_43 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1680" *) flag_l1_42;
  assign flag_l2_22 = flag_l1_45 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1681" *) flag_l1_44;
  assign flag_l2_23 = flag_l1_47 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1682" *) flag_l1_46;
  assign flag_l2_24 = flag_l1_49 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1683" *) flag_l1_48;
  assign flag_l2_25 = flag_l1_51 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1684" *) flag_l1_50;
  assign flag_l2_26 = flag_l1_53 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1685" *) flag_l1_52;
  assign flag_l2_27 = flag_l1_55 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1686" *) flag_l1_54;
  assign flag_l2_28 = flag_l1_57 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1687" *) flag_l1_56;
  assign flag_l2_29 = flag_l1_59 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1688" *) flag_l1_58;
  assign flag_l2_30 = flag_l1_61 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1689" *) flag_l1_60;
  assign flag_l3_0 = flag_l2_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1690" *) flag_l2_0;
  assign flag_l3_1 = flag_l2_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1691" *) flag_l2_2;
  assign flag_l3_2 = flag_l2_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1692" *) flag_l2_4;
  assign flag_l3_3 = flag_l2_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1693" *) flag_l2_6;
  assign flag_l3_4 = flag_l2_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1694" *) flag_l2_8;
  assign flag_l3_5 = flag_l2_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1695" *) flag_l2_10;
  assign flag_l3_6 = flag_l2_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1696" *) flag_l2_12;
  assign flag_l3_7 = flag_l2_15 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1697" *) flag_l2_14;
  assign flag_l3_8 = flag_l2_17 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1698" *) flag_l2_16;
  assign flag_l3_9 = flag_l2_19 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1699" *) flag_l2_18;
  assign flag_l3_10 = flag_l2_21 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1700" *) flag_l2_20;
  assign flag_l3_11 = flag_l2_23 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1701" *) flag_l2_22;
  assign flag_l3_12 = flag_l2_25 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1702" *) flag_l2_24;
  assign flag_l3_13 = flag_l2_27 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1703" *) flag_l2_26;
  assign flag_l3_14 = flag_l2_29 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1704" *) flag_l2_28;
  assign flag_l4_0 = flag_l3_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1705" *) flag_l3_0;
  assign flag_l4_1 = flag_l3_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1706" *) flag_l3_2;
  assign flag_l4_2 = flag_l3_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1707" *) flag_l3_4;
  assign flag_l4_3 = flag_l3_7 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1708" *) flag_l3_6;
  assign flag_l4_4 = flag_l3_9 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1709" *) flag_l3_8;
  assign flag_l4_5 = flag_l3_11 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1710" *) flag_l3_10;
  assign flag_l4_6 = flag_l3_13 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1711" *) flag_l3_12;
  assign flag_l5_0 = flag_l4_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1712" *) flag_l4_0;
  assign flag_l5_1 = flag_l4_3 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1713" *) flag_l4_2;
  assign flag_l5_2 = flag_l4_5 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1714" *) flag_l4_4;
  assign flag_l6_0 = flag_l5_1 | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1715" *) flag_l5_0;
  assign _1724_ = cq_rd_credit[0] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2401" *) rd_take0;
  assign _1725_ = cq_rd_credit[1] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2497" *) rd_take1;
  assign _1726_ = cq_rd_credit[2] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2593" *) rd_take2;
  assign _1727_ = cq_rd_credit[3] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2689" *) rd_take3;
  assign _1728_ = cq_rd_credit[4] | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2785" *) rd_take4;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_take_thread_id_last <= 3'b000;
    else
      cq_rd_take_thread_id_last <= _0016_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd4_credits <= 9'b000000000;
    else
      cq_rd4_credits <= _0008_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd4_credits_ne0 <= 1'b0;
    else
      cq_rd4_credits_ne0 <= _0009_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid4_0_vld <= 1'b0;
    else
      rd_skid4_0_vld <= _0051_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid4_1_vld <= 1'b0;
    else
      rd_skid4_1_vld <= _0053_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid4_2_vld <= 1'b0;
    else
      rd_skid4_2_vld <= _0055_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid4_0 <= _0050_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid4_1 <= _0052_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid4_2 <= _0054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd4_prdy_d <= 1'b1;
    else
      cq_rd4_prdy_d <= cq_rd4_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd3_credits <= 9'b000000000;
    else
      cq_rd3_credits <= _0006_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd3_credits_ne0 <= 1'b0;
    else
      cq_rd3_credits_ne0 <= _0007_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid3_0_vld <= 1'b0;
    else
      rd_skid3_0_vld <= _0045_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid3_1_vld <= 1'b0;
    else
      rd_skid3_1_vld <= _0047_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid3_2_vld <= 1'b0;
    else
      rd_skid3_2_vld <= _0049_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid3_0 <= _0044_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid3_1 <= _0046_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid3_2 <= _0048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd3_prdy_d <= 1'b1;
    else
      cq_rd3_prdy_d <= cq_rd3_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd2_credits <= 9'b000000000;
    else
      cq_rd2_credits <= _0004_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd2_credits_ne0 <= 1'b0;
    else
      cq_rd2_credits_ne0 <= _0005_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid2_0_vld <= 1'b0;
    else
      rd_skid2_0_vld <= _0039_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid2_1_vld <= 1'b0;
    else
      rd_skid2_1_vld <= _0041_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid2_2_vld <= 1'b0;
    else
      rd_skid2_2_vld <= _0043_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid2_0 <= _0038_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid2_1 <= _0040_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid2_2 <= _0042_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd2_prdy_d <= 1'b1;
    else
      cq_rd2_prdy_d <= cq_rd2_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd1_credits <= 9'b000000000;
    else
      cq_rd1_credits <= _0002_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd1_credits_ne0 <= 1'b0;
    else
      cq_rd1_credits_ne0 <= _0003_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid1_0_vld <= 1'b0;
    else
      rd_skid1_0_vld <= _0033_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid1_1_vld <= 1'b0;
    else
      rd_skid1_1_vld <= _0035_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid1_2_vld <= 1'b0;
    else
      rd_skid1_2_vld <= _0037_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid1_0 <= _0032_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid1_1 <= _0034_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid1_2 <= _0036_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd1_prdy_d <= 1'b1;
    else
      cq_rd1_prdy_d <= cq_rd1_prdy;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd0_credits <= 9'b000000000;
    else
      cq_rd0_credits <= _0000_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd0_credits_ne0 <= 1'b0;
    else
      cq_rd0_credits_ne0 <= _0001_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid0_0_vld <= 1'b0;
    else
      rd_skid0_0_vld <= _0027_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid0_1_vld <= 1'b0;
    else
      rd_skid0_1_vld <= _0029_;
  always @(posedge nvdla_core_clk_mgated_skid or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_skid0_2_vld <= 1'b0;
    else
      rd_skid0_2_vld <= _0031_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid0_0 <= _0026_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid0_1 <= _0028_;
  always @(posedge nvdla_core_clk_mgated_skid)
      rd_skid0_2 <= _0030_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd0_prdy_d <= 1'b1;
    else
      cq_rd0_prdy_d <= cq_rd0_prdy;
  always @(posedge nvdla_core_clk_mgated)
      rd_adr_dly <= _0024_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_take_dly <= 1'b0;
    else
      rd_take_dly <= cq_rd_take;
  always @(posedge nvdla_core_clk_mgated)
      head0 <= _0019_;
  always @(posedge nvdla_core_clk_mgated)
      tail0 <= _0057_;
  always @(posedge nvdla_core_clk_mgated)
      head1 <= _0020_;
  always @(posedge nvdla_core_clk_mgated)
      tail1 <= _0058_;
  always @(posedge nvdla_core_clk_mgated)
      head2 <= _0021_;
  always @(posedge nvdla_core_clk_mgated)
      tail2 <= _0059_;
  always @(posedge nvdla_core_clk_mgated)
      head3 <= _0022_;
  always @(posedge nvdla_core_clk_mgated)
      tail3 <= _0060_;
  always @(posedge nvdla_core_clk_mgated)
      head4 <= _0023_;
  always @(posedge nvdla_core_clk_mgated)
      tail4 <= _0061_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      update_head <= 5'b00000;
    else
      update_head <= _0062_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count0 <= 9'b000000000;
    else
      cq_rd_count0 <= _0010_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count1 <= 9'b000000000;
    else
      cq_rd_count1 <= _0011_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count2 <= 9'b000000000;
    else
      cq_rd_count2 <= _0012_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count3 <= 9'b000000000;
    else
      cq_rd_count3 <= _0013_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_count4 <= 9'b000000000;
    else
      cq_rd_count4 <= _0014_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_take_n_dly <= 5'b00000;
    else
      rd_take_n_dly <= _0056_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_rd_credit <= 5'b00000;
    else
      cq_rd_credit <= _0015_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      rd_pushing_q <= 1'b0;
    else
      rd_pushing_q <= _0025_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      free_adr_mask <= 255'b111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111;
    else
      free_adr_mask <= _0018_;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_wr_busy_int <= 1'b0;
    else
      cq_wr_busy_int <= cq_wr_busy_next;
  always @(posedge nvdla_core_clk_mgated or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      cq_wr_count <= 9'b000000000;
    else
      cq_wr_count <= _0017_;
  assign _0016_ = cq_rd_take ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2832" *) cq_rd_take_thread_id : cq_rd_take_thread_id_last;
  assign _0009_ = _1728_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2785" *) _1785_ : cq_rd4_credits_ne0;
  assign _0008_ = _1728_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2785" *) cq_rd4_credits_next : cq_rd4_credits;
  assign _0054_ = _1208_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2745" *) _1784_ : rd_skid4_2;
  assign _1729_ = _1205_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2735" *) rd_skid4_2 : rd_skid4_1;
  assign _0052_ = _1204_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2733" *) _1784_ : _1729_;
  assign _1730_ = _1201_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2723" *) rd_skid4_1 : rd_skid4_0;
  assign _0050_ = _1200_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2721" *) _1783_ : _1730_;
  assign _0007_ = _1727_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2689" *) _1782_ : cq_rd3_credits_ne0;
  assign _0006_ = _1727_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2689" *) cq_rd3_credits_next : cq_rd3_credits;
  assign _0048_ = _1184_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2649" *) _1781_ : rd_skid3_2;
  assign _1731_ = _1181_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2639" *) rd_skid3_2 : rd_skid3_1;
  assign _0046_ = _1180_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2637" *) _1781_ : _1731_;
  assign _1732_ = _1177_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2627" *) rd_skid3_1 : rd_skid3_0;
  assign _0044_ = _1176_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2625" *) _1780_ : _1732_;
  assign _0005_ = _1726_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2593" *) _1779_ : cq_rd2_credits_ne0;
  assign _0004_ = _1726_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2593" *) cq_rd2_credits_next : cq_rd2_credits;
  assign _0042_ = _1161_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2553" *) _1778_ : rd_skid2_2;
  assign _1733_ = _1157_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2543" *) rd_skid2_2 : rd_skid2_1;
  assign _0040_ = _1156_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2541" *) _1778_ : _1733_;
  assign _1734_ = _1154_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2531" *) rd_skid2_1 : rd_skid2_0;
  assign _0038_ = _1152_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2529" *) _1777_ : _1734_;
  assign _0003_ = _1725_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2497" *) _1776_ : cq_rd1_credits_ne0;
  assign _0002_ = _1725_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2497" *) cq_rd1_credits_next : cq_rd1_credits;
  assign _0036_ = _1137_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2457" *) _1775_ : rd_skid1_2;
  assign _1735_ = _1133_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2447" *) rd_skid1_2 : rd_skid1_1;
  assign _0034_ = _1132_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2445" *) _1775_ : _1735_;
  assign _1736_ = _1130_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2435" *) rd_skid1_1 : rd_skid1_0;
  assign _0032_ = _1129_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2433" *) _1774_ : _1736_;
  assign _0001_ = _1724_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2401" *) _1773_ : cq_rd0_credits_ne0;
  assign _0000_ = _1724_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2401" *) cq_rd0_credits_next : cq_rd0_credits;
  assign _0030_ = _1113_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2361" *) _1772_ : rd_skid0_2;
  assign _1737_ = _1110_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2351" *) rd_skid0_2 : rd_skid0_1;
  assign _0028_ = _1108_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2349" *) _1772_ : _1737_;
  assign _1738_ = _1106_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2339" *) rd_skid0_1 : rd_skid0_0;
  assign _0026_ = _1105_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2337" *) _1771_ : _1738_;
  assign _0024_ = cq_rd_take ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2305" *) adr_ram_rd_adr : rd_adr_dly;
  function [7:0] _3874_;
    input [7:0] a;
    input [39:0] b;
    input [4:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2284|./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2279" *)
    (* parallel_case *)
    casez (s)
      5'b????1:
        _3874_ = b[7:0];
      5'b???1?:
        _3874_ = b[15:8];
      5'b??1??:
        _3874_ = b[23:16];
      5'b?1???:
        _3874_ = b[31:24];
      5'b1????:
        _3874_ = b[39:32];
      default:
        _3874_ = a;
    endcase
  endfunction
  assign adr_ram_rd_adr = _3874_(8'b00000000, { _1766_, _1767_, _1768_, _1769_, _1770_ }, { _0519_, _0521_, _0522_, _0523_, _0524_ });
  function [0:0] _3875_;
    input [0:0] a;
    input [4:0] b;
    input [4:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2260|./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2255" *)
    (* parallel_case *)
    casez (s)
      5'b????1:
        _3875_ = b[0:0];
      5'b???1?:
        _3875_ = b[1:1];
      5'b??1??:
        _3875_ = b[2:2];
      5'b?1???:
        _3875_ = b[3:3];
      5'b1????:
        _3875_ = b[4:4];
      default:
        _3875_ = a;
    endcase
  endfunction
  assign adr_ram_rd_enable = _3875_(1'b0, { _1090_, _1091_, _1092_, _1093_, _1094_ }, { _0519_, _0521_, _0522_, _0523_, _0524_ });
  function [0:0] _3876_;
    input [0:0] a;
    input [4:0] b;
    input [4:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2248|./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2243" *)
    (* parallel_case *)
    casez (s)
      5'b????1:
        _3876_ = b[0:0];
      5'b???1?:
        _3876_ = b[1:1];
      5'b??1??:
        _3876_ = b[2:2];
      5'b?1???:
        _3876_ = b[3:3];
      5'b1????:
        _3876_ = b[4:4];
      default:
        _3876_ = a;
    endcase
  endfunction
  assign adr_ram_wr_enable = _3876_(1'b0, { _1084_, _1085_, _1086_, _1087_, _1088_ }, { _0514_, _0515_, _0516_, _0517_, _0518_ });
  function [7:0] _3877_;
    input [7:0] a;
    input [39:0] b;
    input [4:0] s;
    (* full_case = 32'd1 *)
    (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2236|./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2231" *)
    (* parallel_case *)
    casez (s)
      5'b????1:
        _3877_ = b[7:0];
      5'b???1?:
        _3877_ = b[15:8];
      5'b??1??:
        _3877_ = b[23:16];
      5'b?1???:
        _3877_ = b[31:24];
      5'b1????:
        _3877_ = b[39:32];
      default:
        _3877_ = a;
    endcase
  endfunction
  assign adr_ram_wr_adr = _3877_(8'b00000000, { tail0, tail1, tail2, tail3, tail4 }, { _0514_, _0515_, _0516_, _0517_, _0518_ });
  assign _0061_ = rd_pushing4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2203" *) adr_ram_wr_data : tail4;
  assign _1739_ = update_head[4] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2215" *) adr_ram_rd_data : head4;
  assign _0023_ = _1602_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2213" *) adr_ram_wr_data : _1739_;
  assign _0060_ = rd_pushing3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2188" *) adr_ram_wr_data : tail3;
  assign _1740_ = update_head[3] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2200" *) adr_ram_rd_data : head3;
  assign _0022_ = _1601_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2198" *) adr_ram_wr_data : _1740_;
  assign _0059_ = rd_pushing2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2173" *) adr_ram_wr_data : tail2;
  assign _1741_ = update_head[2] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2185" *) adr_ram_rd_data : head2;
  assign _0021_ = _1600_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2183" *) adr_ram_wr_data : _1741_;
  assign _0058_ = rd_pushing1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2158" *) adr_ram_wr_data : tail1;
  assign _1742_ = update_head[1] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2170" *) adr_ram_rd_data : head1;
  assign _0020_ = _1599_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2168" *) adr_ram_wr_data : _1742_;
  assign _0057_ = rd_pushing0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2143" *) adr_ram_wr_data : tail0;
  assign _1743_ = update_head[0] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2155" *) adr_ram_rd_data : head0;
  assign _0019_ = _1598_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2153" *) adr_ram_wr_data : _1743_;
  assign _0062_ = _1597_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2131" *) update_head_next : update_head;
  assign _0014_ = _1744_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2109" *) rd_count4_next : cq_rd_count4;
  assign _0013_ = _1745_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2100" *) rd_count3_next : cq_rd_count3;
  assign _0012_ = _1746_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2091" *) rd_count2_next : cq_rd_count2;
  assign _0011_ = _1747_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2082" *) rd_count1_next : cq_rd_count1;
  assign _0010_ = _1748_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2073" *) rd_count0_next : cq_rd_count0;
  assign _0056_ = update_rd_take_n_dly ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2023" *) { rd_take4, rd_take3, rd_take2, rd_take1, rd_take0 } : rd_take_n_dly;
  assign _0015_[4] = _1596_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing4 : cq_rd_credit[4];
  assign _0015_[3] = _1596_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing3 : cq_rd_credit[3];
  assign _0015_[2] = _1596_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing2 : cq_rd_credit[2];
  assign _0015_[1] = _1596_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing1 : cq_rd_credit[1];
  assign _0015_[0] = _1596_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing0 : cq_rd_credit[0];
  assign _0025_ = _1596_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1984" *) rd_pushing : rd_pushing_q;
  assign _0291_ = _1055_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1465" *) 1'b0 : free_adr_mask[254];
  assign free_adr_mask_next[254] = _1054_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1463" *) 1'b1 : _0291_;
  assign _0289_ = _1053_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1460" *) 1'b0 : free_adr_mask[253];
  assign free_adr_mask_next[253] = _1052_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1458" *) 1'b1 : _0289_;
  assign _0288_ = _1051_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1455" *) 1'b0 : free_adr_mask[252];
  assign free_adr_mask_next[252] = _1050_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1453" *) 1'b1 : _0288_;
  assign _0287_ = _1049_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1450" *) 1'b0 : free_adr_mask[251];
  assign free_adr_mask_next[251] = _1048_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1448" *) 1'b1 : _0287_;
  assign _0286_ = _1047_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1445" *) 1'b0 : free_adr_mask[250];
  assign free_adr_mask_next[250] = _1046_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1443" *) 1'b1 : _0286_;
  assign _0285_ = _1045_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1440" *) 1'b0 : free_adr_mask[249];
  assign free_adr_mask_next[249] = _1044_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1438" *) 1'b1 : _0285_;
  assign _0283_ = _1043_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1435" *) 1'b0 : free_adr_mask[248];
  assign free_adr_mask_next[248] = _1042_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1433" *) 1'b1 : _0283_;
  assign _0282_ = _1041_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1430" *) 1'b0 : free_adr_mask[247];
  assign free_adr_mask_next[247] = _1040_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1428" *) 1'b1 : _0282_;
  assign _0281_ = _1039_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1425" *) 1'b0 : free_adr_mask[246];
  assign free_adr_mask_next[246] = _1038_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1423" *) 1'b1 : _0281_;
  assign _0280_ = _1037_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1420" *) 1'b0 : free_adr_mask[245];
  assign free_adr_mask_next[245] = _1036_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1418" *) 1'b1 : _0280_;
  assign _0279_ = _1035_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1415" *) 1'b0 : free_adr_mask[244];
  assign free_adr_mask_next[244] = _1034_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1413" *) 1'b1 : _0279_;
  assign _0277_ = _1033_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1410" *) 1'b0 : free_adr_mask[243];
  assign free_adr_mask_next[243] = _1032_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1408" *) 1'b1 : _0277_;
  assign _0276_ = _1031_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1405" *) 1'b0 : free_adr_mask[242];
  assign free_adr_mask_next[242] = _1030_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1403" *) 1'b1 : _0276_;
  assign _0275_ = _1029_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1400" *) 1'b0 : free_adr_mask[241];
  assign free_adr_mask_next[241] = _1028_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1398" *) 1'b1 : _0275_;
  assign _0274_ = _1027_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1395" *) 1'b0 : free_adr_mask[240];
  assign free_adr_mask_next[240] = _1026_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1393" *) 1'b1 : _0274_;
  assign _0273_ = _1025_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1390" *) 1'b0 : free_adr_mask[239];
  assign free_adr_mask_next[239] = _1024_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1388" *) 1'b1 : _0273_;
  assign _0272_ = _1023_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1385" *) 1'b0 : free_adr_mask[238];
  assign free_adr_mask_next[238] = _1022_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1383" *) 1'b1 : _0272_;
  assign _0271_ = _1021_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1380" *) 1'b0 : free_adr_mask[237];
  assign free_adr_mask_next[237] = _1020_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1378" *) 1'b1 : _0271_;
  assign _0270_ = _1019_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1375" *) 1'b0 : free_adr_mask[236];
  assign free_adr_mask_next[236] = _1018_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1373" *) 1'b1 : _0270_;
  assign _0269_ = _1017_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1370" *) 1'b0 : free_adr_mask[235];
  assign free_adr_mask_next[235] = _1016_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1368" *) 1'b1 : _0269_;
  assign _0268_ = _1015_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1365" *) 1'b0 : free_adr_mask[234];
  assign free_adr_mask_next[234] = _1014_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1363" *) 1'b1 : _0268_;
  assign _0266_ = _1013_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1360" *) 1'b0 : free_adr_mask[233];
  assign free_adr_mask_next[233] = _1012_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1358" *) 1'b1 : _0266_;
  assign _0265_ = _1011_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1355" *) 1'b0 : free_adr_mask[232];
  assign free_adr_mask_next[232] = _1010_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1353" *) 1'b1 : _0265_;
  assign _0264_ = _1009_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1350" *) 1'b0 : free_adr_mask[231];
  assign free_adr_mask_next[231] = _1008_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1348" *) 1'b1 : _0264_;
  assign _0263_ = _1007_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1345" *) 1'b0 : free_adr_mask[230];
  assign free_adr_mask_next[230] = _1006_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1343" *) 1'b1 : _0263_;
  assign _0262_ = _1005_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1340" *) 1'b0 : free_adr_mask[229];
  assign free_adr_mask_next[229] = _1004_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1338" *) 1'b1 : _0262_;
  assign _0261_ = _1003_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1335" *) 1'b0 : free_adr_mask[228];
  assign free_adr_mask_next[228] = _1002_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1333" *) 1'b1 : _0261_;
  assign _0260_ = _1001_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1330" *) 1'b0 : free_adr_mask[227];
  assign free_adr_mask_next[227] = _1000_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1328" *) 1'b1 : _0260_;
  assign _0259_ = _0999_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1325" *) 1'b0 : free_adr_mask[226];
  assign free_adr_mask_next[226] = _0998_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1323" *) 1'b1 : _0259_;
  assign _0258_ = _0997_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1320" *) 1'b0 : free_adr_mask[225];
  assign free_adr_mask_next[225] = _0996_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1318" *) 1'b1 : _0258_;
  assign _0257_ = _0995_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1315" *) 1'b0 : free_adr_mask[224];
  assign free_adr_mask_next[224] = _0994_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1313" *) 1'b1 : _0257_;
  assign _0255_ = _0993_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1310" *) 1'b0 : free_adr_mask[223];
  assign free_adr_mask_next[223] = _0992_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1308" *) 1'b1 : _0255_;
  assign _0254_ = _0991_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1305" *) 1'b0 : free_adr_mask[222];
  assign free_adr_mask_next[222] = _0990_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1303" *) 1'b1 : _0254_;
  assign _0253_ = _0989_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1300" *) 1'b0 : free_adr_mask[221];
  assign free_adr_mask_next[221] = _0988_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1298" *) 1'b1 : _0253_;
  assign _0252_ = _0987_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1295" *) 1'b0 : free_adr_mask[220];
  assign free_adr_mask_next[220] = _0986_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1293" *) 1'b1 : _0252_;
  assign _0251_ = _0985_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1290" *) 1'b0 : free_adr_mask[219];
  assign free_adr_mask_next[219] = _0984_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1288" *) 1'b1 : _0251_;
  assign _0250_ = _0983_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1285" *) 1'b0 : free_adr_mask[218];
  assign free_adr_mask_next[218] = _0982_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1283" *) 1'b1 : _0250_;
  assign _0249_ = _0981_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1280" *) 1'b0 : free_adr_mask[217];
  assign free_adr_mask_next[217] = _0980_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1278" *) 1'b1 : _0249_;
  assign _0248_ = _0979_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1275" *) 1'b0 : free_adr_mask[216];
  assign free_adr_mask_next[216] = _0978_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1273" *) 1'b1 : _0248_;
  assign _0247_ = _0977_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1270" *) 1'b0 : free_adr_mask[215];
  assign free_adr_mask_next[215] = _0976_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1268" *) 1'b1 : _0247_;
  assign _0246_ = _0975_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1265" *) 1'b0 : free_adr_mask[214];
  assign free_adr_mask_next[214] = _0974_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1263" *) 1'b1 : _0246_;
  assign _0244_ = _0973_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1260" *) 1'b0 : free_adr_mask[213];
  assign free_adr_mask_next[213] = _0972_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1258" *) 1'b1 : _0244_;
  assign _0243_ = _0971_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1255" *) 1'b0 : free_adr_mask[212];
  assign free_adr_mask_next[212] = _0970_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1253" *) 1'b1 : _0243_;
  assign _0242_ = _0969_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1250" *) 1'b0 : free_adr_mask[211];
  assign free_adr_mask_next[211] = _0968_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1248" *) 1'b1 : _0242_;
  assign _0241_ = _0967_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1245" *) 1'b0 : free_adr_mask[210];
  assign free_adr_mask_next[210] = _0966_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1243" *) 1'b1 : _0241_;
  assign _0240_ = _0965_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1240" *) 1'b0 : free_adr_mask[209];
  assign free_adr_mask_next[209] = _0964_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1238" *) 1'b1 : _0240_;
  assign _0239_ = _0963_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1235" *) 1'b0 : free_adr_mask[208];
  assign free_adr_mask_next[208] = _0962_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1233" *) 1'b1 : _0239_;
  assign _0238_ = _0961_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1230" *) 1'b0 : free_adr_mask[207];
  assign free_adr_mask_next[207] = _0960_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1228" *) 1'b1 : _0238_;
  assign _0237_ = _0959_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1225" *) 1'b0 : free_adr_mask[206];
  assign free_adr_mask_next[206] = _0958_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1223" *) 1'b1 : _0237_;
  assign _0236_ = _0957_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1220" *) 1'b0 : free_adr_mask[205];
  assign free_adr_mask_next[205] = _0956_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1218" *) 1'b1 : _0236_;
  assign _0235_ = _0955_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1215" *) 1'b0 : free_adr_mask[204];
  assign free_adr_mask_next[204] = _0954_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1213" *) 1'b1 : _0235_;
  assign _0233_ = _0953_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1210" *) 1'b0 : free_adr_mask[203];
  assign free_adr_mask_next[203] = _0952_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1208" *) 1'b1 : _0233_;
  assign _0232_ = _0951_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1205" *) 1'b0 : free_adr_mask[202];
  assign free_adr_mask_next[202] = _0950_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1203" *) 1'b1 : _0232_;
  assign _0231_ = _0949_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1200" *) 1'b0 : free_adr_mask[201];
  assign free_adr_mask_next[201] = _0948_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1198" *) 1'b1 : _0231_;
  assign _0230_ = _0947_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1195" *) 1'b0 : free_adr_mask[200];
  assign free_adr_mask_next[200] = _0946_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1193" *) 1'b1 : _0230_;
  assign _0229_ = _0945_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1190" *) 1'b0 : free_adr_mask[199];
  assign free_adr_mask_next[199] = _0944_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1188" *) 1'b1 : _0229_;
  assign _0228_ = _0943_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1185" *) 1'b0 : free_adr_mask[198];
  assign free_adr_mask_next[198] = _0942_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1183" *) 1'b1 : _0228_;
  assign _0227_ = _0941_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1180" *) 1'b0 : free_adr_mask[197];
  assign free_adr_mask_next[197] = _0940_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1178" *) 1'b1 : _0227_;
  assign _0226_ = _0939_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1175" *) 1'b0 : free_adr_mask[196];
  assign free_adr_mask_next[196] = _0938_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1173" *) 1'b1 : _0226_;
  assign _0225_ = _0937_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1170" *) 1'b0 : free_adr_mask[195];
  assign free_adr_mask_next[195] = _0936_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1168" *) 1'b1 : _0225_;
  assign _0224_ = _0935_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1165" *) 1'b0 : free_adr_mask[194];
  assign free_adr_mask_next[194] = _0934_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1163" *) 1'b1 : _0224_;
  assign _0222_ = _0933_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1160" *) 1'b0 : free_adr_mask[193];
  assign free_adr_mask_next[193] = _0932_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1158" *) 1'b1 : _0222_;
  assign _0221_ = _0931_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1155" *) 1'b0 : free_adr_mask[192];
  assign free_adr_mask_next[192] = _0930_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1153" *) 1'b1 : _0221_;
  assign _0220_ = _0929_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1150" *) 1'b0 : free_adr_mask[191];
  assign free_adr_mask_next[191] = _0928_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1148" *) 1'b1 : _0220_;
  assign _0219_ = _0927_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1145" *) 1'b0 : free_adr_mask[190];
  assign free_adr_mask_next[190] = _0926_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1143" *) 1'b1 : _0219_;
  assign _0218_ = _0925_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1140" *) 1'b0 : free_adr_mask[189];
  assign free_adr_mask_next[189] = _0924_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1138" *) 1'b1 : _0218_;
  assign _0217_ = _0923_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1135" *) 1'b0 : free_adr_mask[188];
  assign free_adr_mask_next[188] = _0922_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1133" *) 1'b1 : _0217_;
  assign _0216_ = _0921_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1130" *) 1'b0 : free_adr_mask[187];
  assign free_adr_mask_next[187] = _0920_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1128" *) 1'b1 : _0216_;
  assign _0215_ = _0919_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1125" *) 1'b0 : free_adr_mask[186];
  assign free_adr_mask_next[186] = _0918_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1123" *) 1'b1 : _0215_;
  assign _0214_ = _0917_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1120" *) 1'b0 : free_adr_mask[185];
  assign free_adr_mask_next[185] = _0916_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1118" *) 1'b1 : _0214_;
  assign _0213_ = _0915_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1115" *) 1'b0 : free_adr_mask[184];
  assign free_adr_mask_next[184] = _0914_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1113" *) 1'b1 : _0213_;
  assign _0211_ = _0913_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1110" *) 1'b0 : free_adr_mask[183];
  assign free_adr_mask_next[183] = _0912_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1108" *) 1'b1 : _0211_;
  assign _0210_ = _0911_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1105" *) 1'b0 : free_adr_mask[182];
  assign free_adr_mask_next[182] = _0910_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1103" *) 1'b1 : _0210_;
  assign _0209_ = _0909_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1100" *) 1'b0 : free_adr_mask[181];
  assign free_adr_mask_next[181] = _0908_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1098" *) 1'b1 : _0209_;
  assign _0208_ = _0907_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1095" *) 1'b0 : free_adr_mask[180];
  assign free_adr_mask_next[180] = _0906_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1093" *) 1'b1 : _0208_;
  assign _0207_ = _0905_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1090" *) 1'b0 : free_adr_mask[179];
  assign free_adr_mask_next[179] = _0904_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1088" *) 1'b1 : _0207_;
  assign _0206_ = _0903_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1085" *) 1'b0 : free_adr_mask[178];
  assign free_adr_mask_next[178] = _0902_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1083" *) 1'b1 : _0206_;
  assign _0205_ = _0901_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1080" *) 1'b0 : free_adr_mask[177];
  assign free_adr_mask_next[177] = _0900_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1078" *) 1'b1 : _0205_;
  assign _0204_ = _0899_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1075" *) 1'b0 : free_adr_mask[176];
  assign free_adr_mask_next[176] = _0898_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1073" *) 1'b1 : _0204_;
  assign _0203_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1070" *) 1'b0 : free_adr_mask[175];
  assign free_adr_mask_next[175] = _0896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1068" *) 1'b1 : _0203_;
  assign _0202_ = _0895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1065" *) 1'b0 : free_adr_mask[174];
  assign free_adr_mask_next[174] = _0894_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1063" *) 1'b1 : _0202_;
  assign _0200_ = _0893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1060" *) 1'b0 : free_adr_mask[173];
  assign free_adr_mask_next[173] = _0892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1058" *) 1'b1 : _0200_;
  assign _0199_ = _0891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1055" *) 1'b0 : free_adr_mask[172];
  assign free_adr_mask_next[172] = _0890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1053" *) 1'b1 : _0199_;
  assign _0198_ = _0889_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1050" *) 1'b0 : free_adr_mask[171];
  assign free_adr_mask_next[171] = _0888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1048" *) 1'b1 : _0198_;
  assign _0197_ = _0887_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1045" *) 1'b0 : free_adr_mask[170];
  assign free_adr_mask_next[170] = _0886_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1043" *) 1'b1 : _0197_;
  assign _0196_ = _0885_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1040" *) 1'b0 : free_adr_mask[169];
  assign free_adr_mask_next[169] = _0884_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1038" *) 1'b1 : _0196_;
  assign _0195_ = _0883_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1035" *) 1'b0 : free_adr_mask[168];
  assign free_adr_mask_next[168] = _0882_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1033" *) 1'b1 : _0195_;
  assign _0194_ = _0881_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1030" *) 1'b0 : free_adr_mask[167];
  assign free_adr_mask_next[167] = _0880_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1028" *) 1'b1 : _0194_;
  assign _0193_ = _0879_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1025" *) 1'b0 : free_adr_mask[166];
  assign free_adr_mask_next[166] = _0878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1023" *) 1'b1 : _0193_;
  assign _0192_ = _0877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1020" *) 1'b0 : free_adr_mask[165];
  assign free_adr_mask_next[165] = _0876_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1018" *) 1'b1 : _0192_;
  assign _0191_ = _0875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1015" *) 1'b0 : free_adr_mask[164];
  assign free_adr_mask_next[164] = _0874_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1013" *) 1'b1 : _0191_;
  assign _0189_ = _0873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1010" *) 1'b0 : free_adr_mask[163];
  assign free_adr_mask_next[163] = _0872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1008" *) 1'b1 : _0189_;
  assign _0188_ = _0871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1005" *) 1'b0 : free_adr_mask[162];
  assign free_adr_mask_next[162] = _0870_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1003" *) 1'b1 : _0188_;
  assign _0187_ = _0869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1000" *) 1'b0 : free_adr_mask[161];
  assign free_adr_mask_next[161] = _1548_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:998" *) 1'b1 : _0187_;
  assign _0186_ = _1547_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:995" *) 1'b0 : free_adr_mask[160];
  assign free_adr_mask_next[160] = _1546_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:993" *) 1'b1 : _0186_;
  assign _0185_ = _1545_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:990" *) 1'b0 : free_adr_mask[159];
  assign free_adr_mask_next[159] = _1544_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:988" *) 1'b1 : _0185_;
  assign _0184_ = _1543_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:985" *) 1'b0 : free_adr_mask[158];
  assign free_adr_mask_next[158] = _1542_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:983" *) 1'b1 : _0184_;
  assign _0183_ = _1541_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:980" *) 1'b0 : free_adr_mask[157];
  assign free_adr_mask_next[157] = _1540_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:978" *) 1'b1 : _0183_;
  assign _0182_ = _1539_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:975" *) 1'b0 : free_adr_mask[156];
  assign free_adr_mask_next[156] = _1538_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:973" *) 1'b1 : _0182_;
  assign _0181_ = _1537_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:970" *) 1'b0 : free_adr_mask[155];
  assign free_adr_mask_next[155] = _1536_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:968" *) 1'b1 : _0181_;
  assign _0180_ = _1535_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:965" *) 1'b0 : free_adr_mask[154];
  assign free_adr_mask_next[154] = _1534_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:963" *) 1'b1 : _0180_;
  assign _0178_ = _1533_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:960" *) 1'b0 : free_adr_mask[153];
  assign free_adr_mask_next[153] = _1532_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:958" *) 1'b1 : _0178_;
  assign _0177_ = _1531_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:955" *) 1'b0 : free_adr_mask[152];
  assign free_adr_mask_next[152] = _1530_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:953" *) 1'b1 : _0177_;
  assign _0176_ = _1529_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:950" *) 1'b0 : free_adr_mask[151];
  assign free_adr_mask_next[151] = _1528_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:948" *) 1'b1 : _0176_;
  assign _0175_ = _1527_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:945" *) 1'b0 : free_adr_mask[150];
  assign free_adr_mask_next[150] = _1526_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:943" *) 1'b1 : _0175_;
  assign _0174_ = _1525_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:940" *) 1'b0 : free_adr_mask[149];
  assign free_adr_mask_next[149] = _1524_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:938" *) 1'b1 : _0174_;
  assign _0172_ = _1523_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:935" *) 1'b0 : free_adr_mask[148];
  assign free_adr_mask_next[148] = _1522_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:933" *) 1'b1 : _0172_;
  assign _0171_ = _1521_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:930" *) 1'b0 : free_adr_mask[147];
  assign free_adr_mask_next[147] = _1520_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:928" *) 1'b1 : _0171_;
  assign _0170_ = _1519_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:925" *) 1'b0 : free_adr_mask[146];
  assign free_adr_mask_next[146] = _1518_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:923" *) 1'b1 : _0170_;
  assign _0169_ = _1517_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:920" *) 1'b0 : free_adr_mask[145];
  assign free_adr_mask_next[145] = _1516_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:918" *) 1'b1 : _0169_;
  assign _0168_ = _1515_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:915" *) 1'b0 : free_adr_mask[144];
  assign free_adr_mask_next[144] = _1514_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:913" *) 1'b1 : _0168_;
  assign _0166_ = _1513_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:910" *) 1'b0 : free_adr_mask[143];
  assign free_adr_mask_next[143] = _1512_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:908" *) 1'b1 : _0166_;
  assign _0165_ = _1511_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:905" *) 1'b0 : free_adr_mask[142];
  assign free_adr_mask_next[142] = _1510_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:903" *) 1'b1 : _0165_;
  assign _0164_ = _1509_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:900" *) 1'b0 : free_adr_mask[141];
  assign free_adr_mask_next[141] = _1508_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:898" *) 1'b1 : _0164_;
  assign _0163_ = _1507_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:895" *) 1'b0 : free_adr_mask[140];
  assign free_adr_mask_next[140] = _1506_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:893" *) 1'b1 : _0163_;
  assign _0162_ = _1505_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:890" *) 1'b0 : free_adr_mask[139];
  assign free_adr_mask_next[139] = _1504_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:888" *) 1'b1 : _0162_;
  assign _0161_ = _1503_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:885" *) 1'b0 : free_adr_mask[138];
  assign free_adr_mask_next[138] = _1502_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:883" *) 1'b1 : _0161_;
  assign _0160_ = _1501_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:880" *) 1'b0 : free_adr_mask[137];
  assign free_adr_mask_next[137] = _1500_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:878" *) 1'b1 : _0160_;
  assign _0159_ = _1499_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:875" *) 1'b0 : free_adr_mask[136];
  assign free_adr_mask_next[136] = _1498_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:873" *) 1'b1 : _0159_;
  assign _0158_ = _1497_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:870" *) 1'b0 : free_adr_mask[135];
  assign free_adr_mask_next[135] = _1496_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:868" *) 1'b1 : _0158_;
  assign _0157_ = _1495_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:865" *) 1'b0 : free_adr_mask[134];
  assign free_adr_mask_next[134] = _1494_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:863" *) 1'b1 : _0157_;
  assign _0155_ = _1493_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:860" *) 1'b0 : free_adr_mask[133];
  assign free_adr_mask_next[133] = _1492_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:858" *) 1'b1 : _0155_;
  assign _0154_ = _1491_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:855" *) 1'b0 : free_adr_mask[132];
  assign free_adr_mask_next[132] = _1490_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:853" *) 1'b1 : _0154_;
  assign _0153_ = _1489_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:850" *) 1'b0 : free_adr_mask[131];
  assign free_adr_mask_next[131] = _1488_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:848" *) 1'b1 : _0153_;
  assign _0152_ = _1487_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:845" *) 1'b0 : free_adr_mask[130];
  assign free_adr_mask_next[130] = _1486_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:843" *) 1'b1 : _0152_;
  assign _0151_ = _1485_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:840" *) 1'b0 : free_adr_mask[129];
  assign free_adr_mask_next[129] = _1484_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:838" *) 1'b1 : _0151_;
  assign _0150_ = _1483_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:835" *) 1'b0 : free_adr_mask[128];
  assign free_adr_mask_next[128] = _1482_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:833" *) 1'b1 : _0150_;
  assign _0149_ = _1481_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:830" *) 1'b0 : free_adr_mask[127];
  assign free_adr_mask_next[127] = _1480_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:828" *) 1'b1 : _0149_;
  assign _0148_ = _1479_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:825" *) 1'b0 : free_adr_mask[126];
  assign free_adr_mask_next[126] = _1478_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:823" *) 1'b1 : _0148_;
  assign _0147_ = _1477_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:820" *) 1'b0 : free_adr_mask[125];
  assign free_adr_mask_next[125] = _1476_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:818" *) 1'b1 : _0147_;
  assign _0146_ = _1475_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:815" *) 1'b0 : free_adr_mask[124];
  assign free_adr_mask_next[124] = _1474_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:813" *) 1'b1 : _0146_;
  assign _0144_ = _1473_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:810" *) 1'b0 : free_adr_mask[123];
  assign free_adr_mask_next[123] = _1472_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:808" *) 1'b1 : _0144_;
  assign _0143_ = _1471_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:805" *) 1'b0 : free_adr_mask[122];
  assign free_adr_mask_next[122] = _1470_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:803" *) 1'b1 : _0143_;
  assign _0142_ = _1469_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:800" *) 1'b0 : free_adr_mask[121];
  assign free_adr_mask_next[121] = _1468_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:798" *) 1'b1 : _0142_;
  assign _0141_ = _1467_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:795" *) 1'b0 : free_adr_mask[120];
  assign free_adr_mask_next[120] = _1466_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:793" *) 1'b1 : _0141_;
  assign _0140_ = _1465_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:790" *) 1'b0 : free_adr_mask[119];
  assign free_adr_mask_next[119] = _1464_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:788" *) 1'b1 : _0140_;
  assign _0139_ = _1463_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:785" *) 1'b0 : free_adr_mask[118];
  assign free_adr_mask_next[118] = _1462_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:783" *) 1'b1 : _0139_;
  assign _0138_ = _1461_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:780" *) 1'b0 : free_adr_mask[117];
  assign free_adr_mask_next[117] = _1460_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:778" *) 1'b1 : _0138_;
  assign _0137_ = _1459_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:775" *) 1'b0 : free_adr_mask[116];
  assign free_adr_mask_next[116] = _1458_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:773" *) 1'b1 : _0137_;
  assign _0136_ = _1457_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:770" *) 1'b0 : free_adr_mask[115];
  assign free_adr_mask_next[115] = _1456_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:768" *) 1'b1 : _0136_;
  assign _0135_ = _1455_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:765" *) 1'b0 : free_adr_mask[114];
  assign free_adr_mask_next[114] = _1454_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:763" *) 1'b1 : _0135_;
  assign _0133_ = _1453_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:760" *) 1'b0 : free_adr_mask[113];
  assign free_adr_mask_next[113] = _1452_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:758" *) 1'b1 : _0133_;
  assign _0132_ = _1451_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:755" *) 1'b0 : free_adr_mask[112];
  assign free_adr_mask_next[112] = _1450_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:753" *) 1'b1 : _0132_;
  assign _0131_ = _1449_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:750" *) 1'b0 : free_adr_mask[111];
  assign free_adr_mask_next[111] = _1448_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:748" *) 1'b1 : _0131_;
  assign _0130_ = _1447_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:745" *) 1'b0 : free_adr_mask[110];
  assign free_adr_mask_next[110] = _1446_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:743" *) 1'b1 : _0130_;
  assign _0129_ = _1445_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:740" *) 1'b0 : free_adr_mask[109];
  assign free_adr_mask_next[109] = _1444_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:738" *) 1'b1 : _0129_;
  assign _0128_ = _1443_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:735" *) 1'b0 : free_adr_mask[108];
  assign free_adr_mask_next[108] = _1442_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:733" *) 1'b1 : _0128_;
  assign _0127_ = _1441_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:730" *) 1'b0 : free_adr_mask[107];
  assign free_adr_mask_next[107] = _1440_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:728" *) 1'b1 : _0127_;
  assign _0126_ = _1439_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:725" *) 1'b0 : free_adr_mask[106];
  assign free_adr_mask_next[106] = _1438_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:723" *) 1'b1 : _0126_;
  assign _0125_ = _1437_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:720" *) 1'b0 : free_adr_mask[105];
  assign free_adr_mask_next[105] = _1436_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:718" *) 1'b1 : _0125_;
  assign _0124_ = _1435_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:715" *) 1'b0 : free_adr_mask[104];
  assign free_adr_mask_next[104] = _1434_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:713" *) 1'b1 : _0124_;
  assign _0122_ = _1433_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:710" *) 1'b0 : free_adr_mask[103];
  assign free_adr_mask_next[103] = _1432_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:708" *) 1'b1 : _0122_;
  assign _0121_ = _1431_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:705" *) 1'b0 : free_adr_mask[102];
  assign free_adr_mask_next[102] = _1430_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:703" *) 1'b1 : _0121_;
  assign _0120_ = _1429_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:700" *) 1'b0 : free_adr_mask[101];
  assign free_adr_mask_next[101] = _1428_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:698" *) 1'b1 : _0120_;
  assign _0119_ = _1427_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:695" *) 1'b0 : free_adr_mask[100];
  assign free_adr_mask_next[100] = _1426_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:693" *) 1'b1 : _0119_;
  assign _0118_ = _1425_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:690" *) 1'b0 : free_adr_mask[99];
  assign free_adr_mask_next[99] = _1424_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:688" *) 1'b1 : _0118_;
  assign _0117_ = _1423_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:685" *) 1'b0 : free_adr_mask[98];
  assign free_adr_mask_next[98] = _1422_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:683" *) 1'b1 : _0117_;
  assign _0116_ = _1421_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:680" *) 1'b0 : free_adr_mask[97];
  assign free_adr_mask_next[97] = _1420_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:678" *) 1'b1 : _0116_;
  assign _0115_ = _1419_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:675" *) 1'b0 : free_adr_mask[96];
  assign free_adr_mask_next[96] = _1418_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:673" *) 1'b1 : _0115_;
  assign _0114_ = _1417_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:670" *) 1'b0 : free_adr_mask[95];
  assign free_adr_mask_next[95] = _1416_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:668" *) 1'b1 : _0114_;
  assign _0113_ = _1415_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:665" *) 1'b0 : free_adr_mask[94];
  assign free_adr_mask_next[94] = _1414_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:663" *) 1'b1 : _0113_;
  assign _0111_ = _1413_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:660" *) 1'b0 : free_adr_mask[93];
  assign free_adr_mask_next[93] = _1412_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:658" *) 1'b1 : _0111_;
  assign _0110_ = _1411_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:655" *) 1'b0 : free_adr_mask[92];
  assign free_adr_mask_next[92] = _1410_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:653" *) 1'b1 : _0110_;
  assign _0109_ = _1409_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:650" *) 1'b0 : free_adr_mask[91];
  assign free_adr_mask_next[91] = _1408_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:648" *) 1'b1 : _0109_;
  assign _0108_ = _1407_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:645" *) 1'b0 : free_adr_mask[90];
  assign free_adr_mask_next[90] = _1406_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:643" *) 1'b1 : _0108_;
  assign _0107_ = _1405_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:640" *) 1'b0 : free_adr_mask[89];
  assign free_adr_mask_next[89] = _1404_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:638" *) 1'b1 : _0107_;
  assign _0106_ = _1403_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:635" *) 1'b0 : free_adr_mask[88];
  assign free_adr_mask_next[88] = _1402_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:633" *) 1'b1 : _0106_;
  assign _0105_ = _1401_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:630" *) 1'b0 : free_adr_mask[87];
  assign free_adr_mask_next[87] = _1400_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:628" *) 1'b1 : _0105_;
  assign _0104_ = _1399_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:625" *) 1'b0 : free_adr_mask[86];
  assign free_adr_mask_next[86] = _1398_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:623" *) 1'b1 : _0104_;
  assign _0103_ = _1397_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:620" *) 1'b0 : free_adr_mask[85];
  assign free_adr_mask_next[85] = _1396_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:618" *) 1'b1 : _0103_;
  assign _0102_ = _1395_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:615" *) 1'b0 : free_adr_mask[84];
  assign free_adr_mask_next[84] = _1394_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:613" *) 1'b1 : _0102_;
  assign _0100_ = _1393_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:610" *) 1'b0 : free_adr_mask[83];
  assign free_adr_mask_next[83] = _1392_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:608" *) 1'b1 : _0100_;
  assign _0099_ = _1391_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:605" *) 1'b0 : free_adr_mask[82];
  assign free_adr_mask_next[82] = _1390_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:603" *) 1'b1 : _0099_;
  assign _0098_ = _1389_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:600" *) 1'b0 : free_adr_mask[81];
  assign free_adr_mask_next[81] = _1388_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:598" *) 1'b1 : _0098_;
  assign _0097_ = _1387_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:595" *) 1'b0 : free_adr_mask[80];
  assign free_adr_mask_next[80] = _1386_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:593" *) 1'b1 : _0097_;
  assign _0096_ = _1385_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:590" *) 1'b0 : free_adr_mask[79];
  assign free_adr_mask_next[79] = _1384_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:588" *) 1'b1 : _0096_;
  assign _0095_ = _1383_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:585" *) 1'b0 : free_adr_mask[78];
  assign free_adr_mask_next[78] = _1382_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:583" *) 1'b1 : _0095_;
  assign _0094_ = _1381_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:580" *) 1'b0 : free_adr_mask[77];
  assign free_adr_mask_next[77] = _1380_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:578" *) 1'b1 : _0094_;
  assign _0093_ = _1379_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:575" *) 1'b0 : free_adr_mask[76];
  assign free_adr_mask_next[76] = _1378_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:573" *) 1'b1 : _0093_;
  assign _0092_ = _1377_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:570" *) 1'b0 : free_adr_mask[75];
  assign free_adr_mask_next[75] = _1376_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:568" *) 1'b1 : _0092_;
  assign _0091_ = _1375_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:565" *) 1'b0 : free_adr_mask[74];
  assign free_adr_mask_next[74] = _1374_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:563" *) 1'b1 : _0091_;
  assign _0089_ = _1373_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:560" *) 1'b0 : free_adr_mask[73];
  assign free_adr_mask_next[73] = _1372_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:558" *) 1'b1 : _0089_;
  assign _0088_ = _1371_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:555" *) 1'b0 : free_adr_mask[72];
  assign free_adr_mask_next[72] = _1370_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:553" *) 1'b1 : _0088_;
  assign _0087_ = _1369_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:550" *) 1'b0 : free_adr_mask[71];
  assign free_adr_mask_next[71] = _1368_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:548" *) 1'b1 : _0087_;
  assign _0086_ = _1367_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:545" *) 1'b0 : free_adr_mask[70];
  assign free_adr_mask_next[70] = _1366_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:543" *) 1'b1 : _0086_;
  assign _0085_ = _1365_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:540" *) 1'b0 : free_adr_mask[69];
  assign free_adr_mask_next[69] = _1364_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:538" *) 1'b1 : _0085_;
  assign _0084_ = _1363_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:535" *) 1'b0 : free_adr_mask[68];
  assign free_adr_mask_next[68] = _1362_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:533" *) 1'b1 : _0084_;
  assign _0083_ = _1361_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:530" *) 1'b0 : free_adr_mask[67];
  assign free_adr_mask_next[67] = _1360_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:528" *) 1'b1 : _0083_;
  assign _0082_ = _1359_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:525" *) 1'b0 : free_adr_mask[66];
  assign free_adr_mask_next[66] = _1358_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:523" *) 1'b1 : _0082_;
  assign _0081_ = _1357_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:520" *) 1'b0 : free_adr_mask[65];
  assign free_adr_mask_next[65] = _1356_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:518" *) 1'b1 : _0081_;
  assign _0080_ = _1355_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:515" *) 1'b0 : free_adr_mask[64];
  assign free_adr_mask_next[64] = _1354_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:513" *) 1'b1 : _0080_;
  assign _0078_ = _1353_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:510" *) 1'b0 : free_adr_mask[63];
  assign free_adr_mask_next[63] = _1352_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:508" *) 1'b1 : _0078_;
  assign _0077_ = _1351_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:505" *) 1'b0 : free_adr_mask[62];
  assign free_adr_mask_next[62] = _1350_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:503" *) 1'b1 : _0077_;
  assign _0076_ = _1349_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:500" *) 1'b0 : free_adr_mask[61];
  assign free_adr_mask_next[61] = _1348_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:498" *) 1'b1 : _0076_;
  assign _0075_ = _1347_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:495" *) 1'b0 : free_adr_mask[60];
  assign free_adr_mask_next[60] = _1346_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:493" *) 1'b1 : _0075_;
  assign _0074_ = _1345_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:490" *) 1'b0 : free_adr_mask[59];
  assign free_adr_mask_next[59] = _1344_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:488" *) 1'b1 : _0074_;
  assign _0073_ = _1343_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:485" *) 1'b0 : free_adr_mask[58];
  assign free_adr_mask_next[58] = _1342_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:483" *) 1'b1 : _0073_;
  assign _0072_ = _1341_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:480" *) 1'b0 : free_adr_mask[57];
  assign free_adr_mask_next[57] = _1340_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:478" *) 1'b1 : _0072_;
  assign _0071_ = _1339_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:475" *) 1'b0 : free_adr_mask[56];
  assign free_adr_mask_next[56] = _1338_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:473" *) 1'b1 : _0071_;
  assign _0070_ = _1337_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:470" *) 1'b0 : free_adr_mask[55];
  assign free_adr_mask_next[55] = _1336_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:468" *) 1'b1 : _0070_;
  assign _0069_ = _1335_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:465" *) 1'b0 : free_adr_mask[54];
  assign free_adr_mask_next[54] = _1334_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:463" *) 1'b1 : _0069_;
  assign _0067_ = _1333_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:460" *) 1'b0 : free_adr_mask[53];
  assign free_adr_mask_next[53] = _1332_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:458" *) 1'b1 : _0067_;
  assign _0066_ = _1331_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:455" *) 1'b0 : free_adr_mask[52];
  assign free_adr_mask_next[52] = _1330_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:453" *) 1'b1 : _0066_;
  assign _0065_ = _1329_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:450" *) 1'b0 : free_adr_mask[51];
  assign free_adr_mask_next[51] = _1328_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:448" *) 1'b1 : _0065_;
  assign _0064_ = _1327_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:445" *) 1'b0 : free_adr_mask[50];
  assign free_adr_mask_next[50] = _1326_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:443" *) 1'b1 : _0064_;
  assign _0063_ = _1325_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:440" *) 1'b0 : free_adr_mask[49];
  assign free_adr_mask_next[49] = _1324_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:438" *) 1'b1 : _0063_;
  assign _0317_ = _1323_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:435" *) 1'b0 : free_adr_mask[48];
  assign free_adr_mask_next[48] = _1322_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:433" *) 1'b1 : _0317_;
  assign _0316_ = _1321_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:430" *) 1'b0 : free_adr_mask[47];
  assign free_adr_mask_next[47] = _1320_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:428" *) 1'b1 : _0316_;
  assign _0315_ = _1319_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:425" *) 1'b0 : free_adr_mask[46];
  assign free_adr_mask_next[46] = _1318_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:423" *) 1'b1 : _0315_;
  assign _0314_ = _1317_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:420" *) 1'b0 : free_adr_mask[45];
  assign free_adr_mask_next[45] = _1316_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:418" *) 1'b1 : _0314_;
  assign _0313_ = _1315_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:415" *) 1'b0 : free_adr_mask[44];
  assign free_adr_mask_next[44] = _1314_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:413" *) 1'b1 : _0313_;
  assign _0311_ = _1313_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:410" *) 1'b0 : free_adr_mask[43];
  assign free_adr_mask_next[43] = _1312_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:408" *) 1'b1 : _0311_;
  assign _0310_ = _1311_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:405" *) 1'b0 : free_adr_mask[42];
  assign free_adr_mask_next[42] = _1310_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:403" *) 1'b1 : _0310_;
  assign _0309_ = _1309_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:400" *) 1'b0 : free_adr_mask[41];
  assign free_adr_mask_next[41] = _1308_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:398" *) 1'b1 : _0309_;
  assign _0308_ = _1307_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:395" *) 1'b0 : free_adr_mask[40];
  assign free_adr_mask_next[40] = _1306_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:393" *) 1'b1 : _0308_;
  assign _0307_ = _1305_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:390" *) 1'b0 : free_adr_mask[39];
  assign free_adr_mask_next[39] = _1304_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:388" *) 1'b1 : _0307_;
  assign _0306_ = _1303_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:385" *) 1'b0 : free_adr_mask[38];
  assign free_adr_mask_next[38] = _1302_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:383" *) 1'b1 : _0306_;
  assign _0305_ = _1301_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:380" *) 1'b0 : free_adr_mask[37];
  assign free_adr_mask_next[37] = _1300_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:378" *) 1'b1 : _0305_;
  assign _0304_ = _1299_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:375" *) 1'b0 : free_adr_mask[36];
  assign free_adr_mask_next[36] = _1298_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:373" *) 1'b1 : _0304_;
  assign _0303_ = _1297_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:370" *) 1'b0 : free_adr_mask[35];
  assign free_adr_mask_next[35] = _1296_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:368" *) 1'b1 : _0303_;
  assign _0302_ = _1295_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:365" *) 1'b0 : free_adr_mask[34];
  assign free_adr_mask_next[34] = _1294_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:363" *) 1'b1 : _0302_;
  assign _0300_ = _1293_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:360" *) 1'b0 : free_adr_mask[33];
  assign free_adr_mask_next[33] = _1292_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:358" *) 1'b1 : _0300_;
  assign _0299_ = _1291_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:355" *) 1'b0 : free_adr_mask[32];
  assign free_adr_mask_next[32] = _1290_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:353" *) 1'b1 : _0299_;
  assign _0298_ = _1289_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:350" *) 1'b0 : free_adr_mask[31];
  assign free_adr_mask_next[31] = _1288_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:348" *) 1'b1 : _0298_;
  assign _0297_ = _1287_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:345" *) 1'b0 : free_adr_mask[30];
  assign free_adr_mask_next[30] = _1286_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:343" *) 1'b1 : _0297_;
  assign _0296_ = _1285_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:340" *) 1'b0 : free_adr_mask[29];
  assign free_adr_mask_next[29] = _1284_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:338" *) 1'b1 : _0296_;
  assign _0295_ = _1283_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:335" *) 1'b0 : free_adr_mask[28];
  assign free_adr_mask_next[28] = _1282_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:333" *) 1'b1 : _0295_;
  assign _0294_ = _1281_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:330" *) 1'b0 : free_adr_mask[27];
  assign free_adr_mask_next[27] = _1280_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:328" *) 1'b1 : _0294_;
  assign _0293_ = _1279_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:325" *) 1'b0 : free_adr_mask[26];
  assign free_adr_mask_next[26] = _1278_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:323" *) 1'b1 : _0293_;
  assign _0292_ = _1277_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:320" *) 1'b0 : free_adr_mask[25];
  assign free_adr_mask_next[25] = _1276_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:318" *) 1'b1 : _0292_;
  assign _0290_ = _1275_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:315" *) 1'b0 : free_adr_mask[24];
  assign free_adr_mask_next[24] = _1274_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:313" *) 1'b1 : _0290_;
  assign _0278_ = _1273_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:310" *) 1'b0 : free_adr_mask[23];
  assign free_adr_mask_next[23] = _1272_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:308" *) 1'b1 : _0278_;
  assign _0267_ = _1271_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:305" *) 1'b0 : free_adr_mask[22];
  assign free_adr_mask_next[22] = _1270_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:303" *) 1'b1 : _0267_;
  assign _0256_ = _1269_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:300" *) 1'b0 : free_adr_mask[21];
  assign free_adr_mask_next[21] = _1268_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:298" *) 1'b1 : _0256_;
  assign _0245_ = _1267_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:295" *) 1'b0 : free_adr_mask[20];
  assign free_adr_mask_next[20] = _1266_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:293" *) 1'b1 : _0245_;
  assign _0234_ = _1265_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:290" *) 1'b0 : free_adr_mask[19];
  assign free_adr_mask_next[19] = _1264_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:288" *) 1'b1 : _0234_;
  assign _0223_ = _1263_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:285" *) 1'b0 : free_adr_mask[18];
  assign free_adr_mask_next[18] = _1262_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:283" *) 1'b1 : _0223_;
  assign _0212_ = _1221_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:280" *) 1'b0 : free_adr_mask[17];
  assign free_adr_mask_next[17] = _1220_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:278" *) 1'b1 : _0212_;
  assign _0201_ = _1209_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:275" *) 1'b0 : free_adr_mask[16];
  assign free_adr_mask_next[16] = _1202_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:273" *) 1'b1 : _0201_;
  assign _0190_ = _1197_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:270" *) 1'b0 : free_adr_mask[15];
  assign free_adr_mask_next[15] = _1189_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:268" *) 1'b1 : _0190_;
  assign _0179_ = _1185_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:265" *) 1'b0 : free_adr_mask[14];
  assign free_adr_mask_next[14] = _1178_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:263" *) 1'b1 : _0179_;
  assign _0167_ = _1173_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:260" *) 1'b0 : free_adr_mask[13];
  assign free_adr_mask_next[13] = _1165_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:258" *) 1'b1 : _0167_;
  assign _0156_ = _1158_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:255" *) 1'b0 : free_adr_mask[12];
  assign free_adr_mask_next[12] = _1153_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:253" *) 1'b1 : _0156_;
  assign _0145_ = _1149_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:250" *) 1'b0 : free_adr_mask[11];
  assign free_adr_mask_next[11] = _1141_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:248" *) 1'b1 : _0145_;
  assign _0134_ = _1134_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:245" *) 1'b0 : free_adr_mask[10];
  assign free_adr_mask_next[10] = _1126_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:243" *) 1'b1 : _0134_;
  assign _0123_ = _1125_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:240" *) 1'b0 : free_adr_mask[9];
  assign free_adr_mask_next[9] = _1116_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:238" *) 1'b1 : _0123_;
  assign _0112_ = _1109_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:235" *) 1'b0 : free_adr_mask[8];
  assign free_adr_mask_next[8] = _1102_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:233" *) 1'b1 : _0112_;
  assign _0101_ = _1101_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:230" *) 1'b0 : free_adr_mask[7];
  assign free_adr_mask_next[7] = _1100_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:228" *) 1'b1 : _0101_;
  assign _0090_ = _1089_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:225" *) 1'b0 : free_adr_mask[6];
  assign free_adr_mask_next[6] = _1083_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:223" *) 1'b1 : _0090_;
  assign _0079_ = _1079_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:220" *) 1'b0 : free_adr_mask[5];
  assign free_adr_mask_next[5] = _1072_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:218" *) 1'b1 : _0079_;
  assign _0068_ = _1065_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:215" *) 1'b0 : free_adr_mask[4];
  assign free_adr_mask_next[4] = _1064_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:213" *) 1'b1 : _0068_;
  assign _0312_ = _1063_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:210" *) 1'b0 : free_adr_mask[3];
  assign free_adr_mask_next[3] = _1062_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:208" *) 1'b1 : _0312_;
  assign _0301_ = _1061_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:205" *) 1'b0 : free_adr_mask[2];
  assign free_adr_mask_next[2] = _1060_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:203" *) 1'b1 : _0301_;
  assign _0284_ = _1059_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:200" *) 1'b0 : free_adr_mask[1];
  assign free_adr_mask_next[1] = _1058_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:198" *) 1'b1 : _0284_;
  assign _0173_ = _1057_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:195" *) 1'b0 : free_adr_mask[0];
  assign free_adr_mask_next[0] = _1056_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:193" *) 1'b1 : _0173_;
  assign _0018_ = _1595_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:180" *) free_adr_mask_next : free_adr_mask;
  assign _0017_ = _1749_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:129" *) wr_count_next : cq_wr_count;
  assign cq_rd_take = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2799" *) { cq_rd_take_elig[0], cq_rd_take_elig[1], cq_rd_take_elig[2], cq_rd_take_elig[3], cq_rd_take_elig[4] };
  assign cq_rd_take_thread_id[0] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2825" *) { cq_rd_take_thread_id_is_1[0], cq_rd_take_thread_id_is_1[1], cq_rd_take_thread_id_is_1[2], cq_rd_take_thread_id_is_1[3], cq_rd_take_thread_id_is_1[4], cq_rd_take_thread_id_is_3[0], cq_rd_take_thread_id_is_3[1], cq_rd_take_thread_id_is_3[2], cq_rd_take_thread_id_is_3[3], cq_rd_take_thread_id_is_3[4] };
  assign cq_rd_take_thread_id[1] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2826" *) { cq_rd_take_thread_id_is_2[0], cq_rd_take_thread_id_is_2[1], cq_rd_take_thread_id_is_2[2], cq_rd_take_thread_id_is_2[3], cq_rd_take_thread_id_is_2[4], cq_rd_take_thread_id_is_3[0], cq_rd_take_thread_id_is_3[1], cq_rd_take_thread_id_is_3[2], cq_rd_take_thread_id_is_3[3], cq_rd_take_thread_id_is_3[4] };
  assign cq_rd_take_thread_id[2] = | (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2827" *) { cq_rd_take_thread_id_is_4[0], cq_rd_take_thread_id_is_4[1], cq_rd_take_thread_id_is_4[2], cq_rd_take_thread_id_is_4[3], cq_rd_take_thread_id_is_4[4] };
  assign _1750_ = cq_rd_count0 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2052" *) 1'b1;
  assign _1751_ = cq_rd_count1 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2055" *) 1'b1;
  assign _1752_ = cq_rd_count2 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2058" *) 1'b1;
  assign _1753_ = cq_rd_count3 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2061" *) 1'b1;
  assign _1754_ = cq_rd_count4 - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2064" *) 1'b1;
  assign cq_rd0_credits_w_take_next = cq_rd0_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2387" *) 1'b1;
  assign cq_rd1_credits_w_take_next = cq_rd1_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2483" *) 1'b1;
  assign cq_rd2_credits_w_take_next = cq_rd2_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2579" *) 1'b1;
  assign cq_rd3_credits_w_take_next = cq_rd3_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2675" *) 1'b1;
  assign cq_rd4_credits_w_take_next = cq_rd4_credits_wo_take_next - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2771" *) 1'b1;
  assign _1755_ = cq_wr_count - (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:93" *) 1'b1;
  assign index_l1_0[0] = flag_l0_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1844" *) index_l0_0 : index_l0_1;
  assign index_l1_1[0] = flag_l0_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1845" *) index_l0_2 : index_l0_3;
  assign index_l1_2[0] = flag_l0_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1846" *) index_l0_4 : index_l0_5;
  assign index_l1_3[0] = flag_l0_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1847" *) index_l0_6 : index_l0_7;
  assign index_l1_4[0] = flag_l0_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1848" *) index_l0_8 : index_l0_9;
  assign index_l1_5[0] = flag_l0_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1849" *) index_l0_10 : index_l0_11;
  assign index_l1_6[0] = flag_l0_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1850" *) index_l0_12 : index_l0_13;
  assign index_l1_7[0] = flag_l0_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1851" *) index_l0_14 : index_l0_15;
  assign index_l1_8[0] = flag_l0_16 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1852" *) index_l0_16 : index_l0_17;
  assign index_l1_9[0] = flag_l0_18 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1853" *) index_l0_18 : index_l0_19;
  assign index_l1_10[0] = flag_l0_20 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1854" *) index_l0_20 : index_l0_21;
  assign index_l1_11[0] = flag_l0_22 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1855" *) index_l0_22 : index_l0_23;
  assign index_l1_12[0] = flag_l0_24 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1856" *) index_l0_24 : index_l0_25;
  assign index_l1_13[0] = flag_l0_26 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1857" *) index_l0_26 : index_l0_27;
  assign index_l1_14[0] = flag_l0_28 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1858" *) index_l0_28 : index_l0_29;
  assign index_l1_15[0] = flag_l0_30 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1859" *) index_l0_30 : index_l0_31;
  assign index_l1_16[0] = flag_l0_32 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1860" *) index_l0_32 : index_l0_33;
  assign index_l1_17[0] = flag_l0_34 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1861" *) index_l0_34 : index_l0_35;
  assign index_l1_18[0] = flag_l0_36 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1862" *) index_l0_36 : index_l0_37;
  assign index_l1_19[0] = flag_l0_38 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1863" *) index_l0_38 : index_l0_39;
  assign index_l1_20[0] = flag_l0_40 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1864" *) index_l0_40 : index_l0_41;
  assign index_l1_21[0] = flag_l0_42 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1865" *) index_l0_42 : index_l0_43;
  assign index_l1_22[0] = flag_l0_44 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1866" *) index_l0_44 : index_l0_45;
  assign index_l1_23[0] = flag_l0_46 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1867" *) index_l0_46 : index_l0_47;
  assign index_l1_24[0] = flag_l0_48 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1868" *) index_l0_48 : index_l0_49;
  assign index_l1_25[0] = flag_l0_50 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1869" *) index_l0_50 : index_l0_51;
  assign index_l1_26[0] = flag_l0_52 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1870" *) index_l0_52 : index_l0_53;
  assign index_l1_27[0] = flag_l0_54 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1871" *) index_l0_54 : index_l0_55;
  assign index_l1_28[0] = flag_l0_56 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1872" *) index_l0_56 : index_l0_57;
  assign index_l1_29[0] = flag_l0_58 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1873" *) index_l0_58 : index_l0_59;
  assign index_l1_30[0] = flag_l0_60 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1874" *) index_l0_60 : index_l0_61;
  assign index_l1_31[0] = flag_l0_62 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1875" *) index_l0_62 : index_l0_63;
  assign index_l1_32[0] = flag_l0_64 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1876" *) index_l0_64 : index_l0_65;
  assign index_l1_33[0] = flag_l0_66 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1877" *) index_l0_66 : index_l0_67;
  assign index_l1_34[0] = flag_l0_68 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1878" *) index_l0_68 : index_l0_69;
  assign index_l1_35[0] = flag_l0_70 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1879" *) index_l0_70 : index_l0_71;
  assign index_l1_36[0] = flag_l0_72 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1880" *) index_l0_72 : index_l0_73;
  assign index_l1_37[0] = flag_l0_74 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1881" *) index_l0_74 : index_l0_75;
  assign index_l1_38[0] = flag_l0_76 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1882" *) index_l0_76 : index_l0_77;
  assign index_l1_39[0] = flag_l0_78 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1883" *) index_l0_78 : index_l0_79;
  assign index_l1_40[0] = flag_l0_80 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1884" *) index_l0_80 : index_l0_81;
  assign index_l1_41[0] = flag_l0_82 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1885" *) index_l0_82 : index_l0_83;
  assign index_l1_42[0] = flag_l0_84 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1886" *) index_l0_84 : index_l0_85;
  assign index_l1_43[0] = flag_l0_86 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1887" *) index_l0_86 : index_l0_87;
  assign index_l1_44[0] = flag_l0_88 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1888" *) index_l0_88 : index_l0_89;
  assign index_l1_45[0] = flag_l0_90 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1889" *) index_l0_90 : index_l0_91;
  assign index_l1_46[0] = flag_l0_92 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1890" *) index_l0_92 : index_l0_93;
  assign index_l1_47[0] = flag_l0_94 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1891" *) index_l0_94 : index_l0_95;
  assign index_l1_48[0] = flag_l0_96 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1892" *) index_l0_96 : index_l0_97;
  assign index_l1_49[0] = flag_l0_98 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1893" *) index_l0_98 : index_l0_99;
  assign index_l1_50[0] = flag_l0_100 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1894" *) index_l0_100 : index_l0_101;
  assign index_l1_51[0] = flag_l0_102 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1895" *) index_l0_102 : index_l0_103;
  assign index_l1_52[0] = flag_l0_104 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1896" *) index_l0_104 : index_l0_105;
  assign index_l1_53[0] = flag_l0_106 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1897" *) index_l0_106 : index_l0_107;
  assign index_l1_54[0] = flag_l0_108 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1898" *) index_l0_108 : index_l0_109;
  assign index_l1_55[0] = flag_l0_110 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1899" *) index_l0_110 : index_l0_111;
  assign index_l1_56[0] = flag_l0_112 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1900" *) index_l0_112 : index_l0_113;
  assign index_l1_57[0] = flag_l0_114 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1901" *) index_l0_114 : index_l0_115;
  assign index_l1_58[0] = flag_l0_116 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1902" *) index_l0_116 : index_l0_117;
  assign index_l1_59[0] = flag_l0_118 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1903" *) index_l0_118 : index_l0_119;
  assign index_l1_60[0] = flag_l0_120 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1904" *) index_l0_120 : index_l0_121;
  assign index_l1_61[0] = flag_l0_122 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1905" *) index_l0_122 : index_l0_123;
  assign index_l1_62[0] = flag_l0_124 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1906" *) index_l0_124 : index_l0_125;
  assign index_l1_63[0] = flag_l0_126 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1907" *) index_l0_126 : index_l0_127;
  assign index_l2_0[1:0] = flag_l1_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1908" *) index_l1_0 : index_l1_1;
  assign index_l2_1[1:0] = flag_l1_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1909" *) index_l1_2 : index_l1_3;
  assign index_l2_2[1:0] = flag_l1_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1910" *) index_l1_4 : index_l1_5;
  assign index_l2_3[1:0] = flag_l1_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1911" *) index_l1_6 : index_l1_7;
  assign index_l2_4[1:0] = flag_l1_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1912" *) index_l1_8 : index_l1_9;
  assign index_l2_5[1:0] = flag_l1_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1913" *) index_l1_10 : index_l1_11;
  assign index_l2_6[1:0] = flag_l1_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1914" *) index_l1_12 : index_l1_13;
  assign index_l2_7[1:0] = flag_l1_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1915" *) index_l1_14 : index_l1_15;
  assign index_l2_8[1:0] = flag_l1_16 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1916" *) index_l1_16 : index_l1_17;
  assign index_l2_9[1:0] = flag_l1_18 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1917" *) index_l1_18 : index_l1_19;
  assign index_l2_10[1:0] = flag_l1_20 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1918" *) index_l1_20 : index_l1_21;
  assign index_l2_11[1:0] = flag_l1_22 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1919" *) index_l1_22 : index_l1_23;
  assign index_l2_12[1:0] = flag_l1_24 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1920" *) index_l1_24 : index_l1_25;
  assign index_l2_13[1:0] = flag_l1_26 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1921" *) index_l1_26 : index_l1_27;
  assign index_l2_14[1:0] = flag_l1_28 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1922" *) index_l1_28 : index_l1_29;
  assign index_l2_15[1:0] = flag_l1_30 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1923" *) index_l1_30 : index_l1_31;
  assign index_l2_16[1:0] = flag_l1_32 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1924" *) index_l1_32 : index_l1_33;
  assign index_l2_17[1:0] = flag_l1_34 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1925" *) index_l1_34 : index_l1_35;
  assign index_l2_18[1:0] = flag_l1_36 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1926" *) index_l1_36 : index_l1_37;
  assign index_l2_19[1:0] = flag_l1_38 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1927" *) index_l1_38 : index_l1_39;
  assign index_l2_20[1:0] = flag_l1_40 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1928" *) index_l1_40 : index_l1_41;
  assign index_l2_21[1:0] = flag_l1_42 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1929" *) index_l1_42 : index_l1_43;
  assign index_l2_22[1:0] = flag_l1_44 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1930" *) index_l1_44 : index_l1_45;
  assign index_l2_23[1:0] = flag_l1_46 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1931" *) index_l1_46 : index_l1_47;
  assign index_l2_24[1:0] = flag_l1_48 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1932" *) index_l1_48 : index_l1_49;
  assign index_l2_25[1:0] = flag_l1_50 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1933" *) index_l1_50 : index_l1_51;
  assign index_l2_26[1:0] = flag_l1_52 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1934" *) index_l1_52 : index_l1_53;
  assign index_l2_27[1:0] = flag_l1_54 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1935" *) index_l1_54 : index_l1_55;
  assign index_l2_28[1:0] = flag_l1_56 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1936" *) index_l1_56 : index_l1_57;
  assign index_l2_29[1:0] = flag_l1_58 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1937" *) index_l1_58 : index_l1_59;
  assign index_l2_30[1:0] = flag_l1_60 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1938" *) index_l1_60 : index_l1_61;
  assign index_l2_31[1:0] = flag_l1_62 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1939" *) index_l1_62 : index_l1_63;
  assign index_l3_0[2:0] = flag_l2_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1940" *) index_l2_0 : index_l2_1;
  assign index_l3_1[2:0] = flag_l2_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1941" *) index_l2_2 : index_l2_3;
  assign index_l3_2[2:0] = flag_l2_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1942" *) index_l2_4 : index_l2_5;
  assign index_l3_3[2:0] = flag_l2_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1943" *) index_l2_6 : index_l2_7;
  assign index_l3_4[2:0] = flag_l2_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1944" *) index_l2_8 : index_l2_9;
  assign index_l3_5[2:0] = flag_l2_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1945" *) index_l2_10 : index_l2_11;
  assign index_l3_6[2:0] = flag_l2_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1946" *) index_l2_12 : index_l2_13;
  assign index_l3_7[2:0] = flag_l2_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1947" *) index_l2_14 : index_l2_15;
  assign index_l3_8[2:0] = flag_l2_16 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1948" *) index_l2_16 : index_l2_17;
  assign index_l3_9[2:0] = flag_l2_18 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1949" *) index_l2_18 : index_l2_19;
  assign index_l3_10[2:0] = flag_l2_20 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1950" *) index_l2_20 : index_l2_21;
  assign index_l3_11[2:0] = flag_l2_22 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1951" *) index_l2_22 : index_l2_23;
  assign index_l3_12[2:0] = flag_l2_24 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1952" *) index_l2_24 : index_l2_25;
  assign index_l3_13[2:0] = flag_l2_26 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1953" *) index_l2_26 : index_l2_27;
  assign index_l3_14[2:0] = flag_l2_28 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1954" *) index_l2_28 : index_l2_29;
  assign index_l3_15[2:0] = flag_l2_30 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1955" *) index_l2_30 : index_l2_31;
  assign index_l4_0[3:0] = flag_l3_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1956" *) index_l3_0 : index_l3_1;
  assign index_l4_1[3:0] = flag_l3_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1957" *) index_l3_2 : index_l3_3;
  assign index_l4_2[3:0] = flag_l3_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1958" *) index_l3_4 : index_l3_5;
  assign index_l4_3[3:0] = flag_l3_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1959" *) index_l3_6 : index_l3_7;
  assign index_l4_4[3:0] = flag_l3_8 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1960" *) index_l3_8 : index_l3_9;
  assign index_l4_5[3:0] = flag_l3_10 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1961" *) index_l3_10 : index_l3_11;
  assign index_l4_6[3:0] = flag_l3_12 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1962" *) index_l3_12 : index_l3_13;
  assign index_l4_7[3:0] = flag_l3_14 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1963" *) index_l3_14 : index_l3_15;
  assign index_l5_0[4:0] = flag_l4_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1964" *) index_l4_0 : index_l4_1;
  assign index_l5_1[4:0] = flag_l4_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1965" *) index_l4_2 : index_l4_3;
  assign index_l5_2[4:0] = flag_l4_4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1966" *) index_l4_4 : index_l4_5;
  assign index_l5_3[4:0] = flag_l4_6 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1967" *) index_l4_6 : index_l4_7;
  assign index_l6_0[5:0] = flag_l5_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1968" *) index_l5_0 : index_l5_1;
  assign index_l6_1[5:0] = flag_l5_2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1969" *) index_l5_2 : index_l5_3;
  assign adr_ram_wr_data[6:0] = flag_l6_0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:1970" *) index_l6_0 : index_l6_1;
  assign _1756_ = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2051" *) cq_rd_count0 : _0318_;
  assign _1757_ = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2052" *) _1750_ : cq_rd_count0;
  assign rd_count0_next = rd_pushing0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2052" *) _1756_ : _1757_;
  assign _1758_ = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2054" *) cq_rd_count1 : _0319_;
  assign _1759_ = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2055" *) _1751_ : cq_rd_count1;
  assign rd_count1_next = rd_pushing1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2055" *) _1758_ : _1759_;
  assign _1760_ = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2057" *) cq_rd_count2 : _0320_;
  assign _1761_ = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2058" *) _1752_ : cq_rd_count2;
  assign rd_count2_next = rd_pushing2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2058" *) _1760_ : _1761_;
  assign _1762_ = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2060" *) cq_rd_count3 : _0321_;
  assign _1763_ = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2061" *) _1753_ : cq_rd_count3;
  assign rd_count3_next = rd_pushing3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2061" *) _1762_ : _1763_;
  assign _1764_ = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2063" *) cq_rd_count4 : _0322_;
  assign _1765_ = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2064" *) _1754_ : cq_rd_count4;
  assign rd_count4_next = rd_pushing4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2064" *) _1764_ : _1765_;
  assign _1766_ = _1095_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2268" *) adr_ram_rd_data : head0;
  assign _1767_ = _1096_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2269" *) adr_ram_rd_data : head1;
  assign _1768_ = _1097_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2270" *) adr_ram_rd_data : head2;
  assign _1769_ = _1098_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2271" *) adr_ram_rd_data : head3;
  assign _1770_ = _1099_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2272" *) adr_ram_rd_data : head4;
  assign cq_rd0_pd = rd_skid0_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2335" *) rd_skid0_0 : cq_wr_pd;
  assign _1771_ = rd_take_n_dly[0] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2338" *) cq_rd_pd_p : cq_wr_pd;
  assign _1772_ = rd_bypassing0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2350" *) cq_wr_pd : cq_rd_pd_p;
  assign _0027_ = _1103_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2377" *) _1608_ : _1610_;
  assign _0029_ = _1103_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2378" *) _1611_ : _1612_;
  assign _0031_ = _1103_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2380" *) _1117_ : _1611_;
  assign cq_rd0_credits_next = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2389" *) cq_rd0_credits_w_take_next : cq_rd0_credits_wo_take_next;
  assign _1773_ = rd_take0 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2403" *) _1712_ : _1713_;
  assign cq_rd1_pd = rd_skid1_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2431" *) rd_skid1_0 : cq_wr_pd;
  assign _1774_ = rd_take_n_dly[1] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2434" *) cq_rd_pd_p : cq_wr_pd;
  assign _1775_ = rd_bypassing1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2446" *) cq_wr_pd : cq_rd_pd_p;
  assign _0033_ = _1127_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2473" *) _1625_ : _1627_;
  assign _0035_ = _1127_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2474" *) _1628_ : _1629_;
  assign _0037_ = _1127_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2476" *) _1140_ : _1628_;
  assign cq_rd1_credits_next = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2485" *) cq_rd1_credits_w_take_next : cq_rd1_credits_wo_take_next;
  assign _1776_ = rd_take1 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2499" *) _1714_ : _1715_;
  assign cq_rd2_pd = rd_skid2_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2527" *) rd_skid2_0 : cq_wr_pd;
  assign _1777_ = rd_take_n_dly[2] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2530" *) cq_rd_pd_p : cq_wr_pd;
  assign _1778_ = rd_bypassing2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2542" *) cq_wr_pd : cq_rd_pd_p;
  assign _0039_ = _1150_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2569" *) _1642_ : _1644_;
  assign _0041_ = _1150_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2570" *) _1645_ : _1646_;
  assign _0043_ = _1150_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2572" *) _1164_ : _1645_;
  assign cq_rd2_credits_next = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2581" *) cq_rd2_credits_w_take_next : cq_rd2_credits_wo_take_next;
  assign _1779_ = rd_take2 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2595" *) _1716_ : _1717_;
  assign cq_rd3_pd = rd_skid3_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2623" *) rd_skid3_0 : cq_wr_pd;
  assign _1780_ = rd_take_n_dly[3] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2626" *) cq_rd_pd_p : cq_wr_pd;
  assign _1781_ = rd_bypassing3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2638" *) cq_wr_pd : cq_rd_pd_p;
  assign _0045_ = _1174_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2665" *) _1659_ : _1661_;
  assign _0047_ = _1174_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2666" *) _1662_ : _1663_;
  assign _0049_ = _1174_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2668" *) _1188_ : _1662_;
  assign cq_rd3_credits_next = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2677" *) cq_rd3_credits_w_take_next : cq_rd3_credits_wo_take_next;
  assign _1782_ = rd_take3 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2691" *) _1718_ : _1719_;
  assign cq_rd4_pd = rd_skid4_0_vld ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2719" *) rd_skid4_0 : cq_wr_pd;
  assign _1783_ = rd_take_n_dly[4] ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2722" *) cq_rd_pd_p : cq_wr_pd;
  assign _1784_ = rd_bypassing4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2734" *) cq_wr_pd : cq_rd_pd_p;
  assign _0051_ = _1198_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2761" *) _1676_ : _1678_;
  assign _0053_ = _1198_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2762" *) _1679_ : _1680_;
  assign _0055_ = _1198_ ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2764" *) _1212_ : _1679_;
  assign cq_rd4_credits_next = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2773" *) cq_rd4_credits_w_take_next : cq_rd4_credits_wo_take_next;
  assign _1785_ = rd_take4 ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2787" *) _1720_ : _1721_;
  assign wr_count_next_wr_popping = rd_pushing ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:93" *) cq_wr_count : _1755_;
  assign wr_count_next_no_wr_popping = rd_pushing ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:94" *) _0323_ : cq_wr_count;
  assign wr_count_next = rd_take_dly ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:96" *) wr_count_next_wr_popping : wr_count_next_no_wr_popping;
  assign cq_wr_busy_next = rd_take_dly ? (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:99" *) 1'b0 : wr_count_next_no_wr_popping_is_256;
  assign _1749_ = rd_pushing ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:129" *) rd_take_dly;
  assign _1748_ = rd_pushing0 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2073" *) rd_take0;
  assign _1747_ = rd_pushing1 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2082" *) rd_take1;
  assign _1746_ = rd_pushing2 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2091" *) rd_take2;
  assign _1745_ = rd_pushing3 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2100" *) rd_take3;
  assign _1744_ = rd_pushing4 ^ (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2109" *) rd_take4;
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:2219" *)
  nv_ram_rwst_256x8 adr_ram (
    .clk(nvdla_core_clk),
    .di(adr_ram_wr_data),
    .dout(adr_ram_rd_data),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(adr_ram_rd_adr),
    .re(adr_ram_rd_enable),
    .wa(adr_ram_wr_adr),
    .we(adr_ram_wr_enable)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:76" *)
  NV_CLK_gate_power nvdla_core_clk_mgate (
    .clk(nvdla_core_clk),
    .clk_en(nvdla_core_clk_mgated_enable),
    .clk_gated(nvdla_core_clk_mgated),
    .reset_(nvdla_core_rstn)
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:73" *)
  NV_CLK_gate_power nvdla_core_clk_rd_mgate_skid (
    .clk(nvdla_core_clk),
    .clk_en(nvdla_core_clk_mgated_skid_enable),
    .clk_gated(nvdla_core_clk_mgated_skid),
    .reset_(nvdla_core_rstn)
  );
  (* src = "./vmod/nvdla/nocif/NV_NVDLA_CVIF_WRITE_cq.v:151" *)
  \$paramod\nv_ram_rws_256x3\FORCE_CONTENTION_ASSERTION_RESET_ACTIVE=1'1  ram (
    .clk(nvdla_core_clk),
    .di(cq_wr_pd),
    .dout(cq_rd_pd_p),
    .pwrbus_ram_pd(pwrbus_ram_pd),
    .ra(adr_ram_rd_adr),
    .re(cq_rd_take),
    .wa(adr_ram_wr_data),
    .we(rd_pushing)
  );
  assign cq_rd_adr = adr_ram_rd_adr;
  assign cq_rd_adr_p = adr_ram_rd_adr;
  assign cq_wr_adr = adr_ram_wr_data;
  assign free_adr_index = adr_ram_wr_data;
  assign index_l7_0 = adr_ram_wr_data;
  assign rd_enable = cq_rd_take;
  assign rd_popping = rd_take_dly;
  assign rd_popping_adr = rd_adr_dly;
  assign rd_pushing_adr = adr_ram_wr_data;
  assign rd_pushing_thread_id = cq_wr_thread_id;
  assign rd_take_dly_cg = rd_take_dly;
  assign wr_adr_popping = rd_pushing;
  assign wr_count_next_is_256 = cq_wr_busy_next;
  assign wr_limit_muxed = 9'b000000000;
  assign wr_limit_reg = 9'b000000000;
  assign wr_popping = rd_take_dly;
  assign wr_pushing = rd_pushing;
  assign wr_pushing_thread_id = cq_wr_thread_id;
  assign wr_reserving_and_not_bypassing = rd_pushing;
endmodule
