module CSC_chn_data_in_rsci_unreg(in_0, outsig);
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:507" *)
  input in_0;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:508" *)
  output outsig;
  assign outsig = in_0;
endmodule
