module FP16_TO_FP32_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp16_to_fp32.v:206" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp16_to_fp32.v:207" *)
  output outsig;
  assign outsig = in_0;
endmodule
