module CSC_leading_sign_23_0(mantissa, rtn);
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:455" *)
  wire _000_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *)
  wire _001_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:466" *)
  wire _002_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *)
  wire _003_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *)
  wire _004_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:468" *)
  wire _005_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *)
  wire _006_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *)
  wire _007_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _008_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _009_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _010_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _011_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _012_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _013_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _014_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _015_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _016_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _017_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *)
  wire _018_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *)
  wire _019_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *)
  wire _020_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:447" *)
  wire _021_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:454" *)
  wire _022_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _023_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:443" *)
  wire _024_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:444" *)
  wire _025_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:445" *)
  wire _026_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:449" *)
  wire _027_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:450" *)
  wire _028_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:451" *)
  wire _029_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:456" *)
  wire _030_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:457" *)
  wire _031_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:458" *)
  wire _032_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *)
  wire _033_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _034_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _035_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _036_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _037_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:461" *)
  wire _038_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *)
  wire _039_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *)
  wire _040_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *)
  wire _041_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *)
  wire _042_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *)
  wire _043_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *)
  wire _044_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *)
  wire _045_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *)
  wire _046_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _047_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _048_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _049_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _050_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _051_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _052_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _053_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _054_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _055_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _056_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _057_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _058_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _059_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _060_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *)
  wire _061_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *)
  wire _062_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *)
  wire _063_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:465" *)
  wire _064_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *)
  wire _065_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *)
  wire _066_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *)
  wire _067_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _068_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *)
  wire _069_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *)
  wire _070_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *)
  wire _071_;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:441" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:439" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:438" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:440" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:428" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:423" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:429" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:424" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:430" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:425" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:431" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:426" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:432" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:427" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:422" *)
  wire IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:437" *)
  wire c_h_1_10;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:433" *)
  wire c_h_1_2;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:434" *)
  wire c_h_1_5;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:435" *)
  wire c_h_1_6;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:436" *)
  wire c_h_1_9;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:419" *)
  input [22:0] mantissa;
  (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:420" *)
  output [4:0] rtn;
  assign c_h_1_2 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:446" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3 = _021_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:448" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1;
  assign c_h_1_5 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:452" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2;
  assign c_h_1_6 = c_h_1_2 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:453" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign _000_ = _022_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:455" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4 = _000_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:455" *) c_h_1_5;
  assign c_h_1_9 = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:459" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2;
  assign c_h_1_10 = c_h_1_6 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:460" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl = c_h_1_6 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:461" *) _038_;
  assign _001_ = c_h_1_2 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *) _062_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl = _001_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *) _063_;
  assign _002_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:466" *) _064_;
  assign _003_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *) _065_;
  assign _004_ = _041_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *) c_h_1_6;
  assign _005_ = _002_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:468" *) _042_;
  assign _006_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *) _066_;
  assign _007_ = _043_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *) c_h_1_10;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl = _005_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *) _044_;
  assign _008_ = _068_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) c_h_1_2;
  assign _009_ = _046_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _048_;
  assign _010_ = _070_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) c_h_1_5;
  assign _011_ = _050_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) _052_;
  assign _012_ = _053_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) c_h_1_6;
  assign _013_ = _009_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) _054_;
  assign _014_ = _057_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) c_h_1_9;
  assign _015_ = _056_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) _058_;
  assign _016_ = _059_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) c_h_1_10;
  assign _017_ = _013_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) _060_;
  assign _018_ = _061_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1;
  assign _019_ = _018_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *) c_h_1_9;
  assign _020_ = _019_ & (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *) c_h_1_10;
  assign _021_ = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:447" *) mantissa[16:15];
  assign _022_ = ! (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:454" *) mantissa[8:7];
  assign _023_ = mantissa[2:1] == (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) 1'b1;
  assign _024_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:443" *) mantissa[20:19];
  assign _025_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:444" *) mantissa[22:21];
  assign _026_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:445" *) mantissa[18:17];
  assign _027_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:449" *) mantissa[12:11];
  assign _028_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:450" *) mantissa[14:13];
  assign _029_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:451" *) mantissa[10:9];
  assign _030_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:456" *) mantissa[4:3];
  assign _031_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:457" *) mantissa[6:5];
  assign _032_ = | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:458" *) mantissa[2:1];
  assign _033_ = mantissa[21:20] != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *) 1'b1;
  assign _034_ = mantissa[17:16] != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) 1'b1;
  assign _035_ = mantissa[13:12] != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) 1'b1;
  assign _036_ = mantissa[9:8] != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) 1'b1;
  assign _037_ = mantissa[5:4] != (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) 1'b1;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_2 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:443" *) _024_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_6_2_sdt_1 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:444" *) _025_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:445" *) _026_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_2 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:449" *) _027_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_26_2_sdt_1 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:450" *) _028_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:451" *) _029_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_2 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:456" *) _030_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_50_2_sdt_1 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:457" *) _031_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:458" *) _032_;
  assign _038_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:461" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_42_4_sdt_4;
  assign _039_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *) IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_18_3_sdt_3;
  assign _040_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *) c_h_1_10;
  assign _041_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *) _003_;
  assign _042_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *) _004_;
  assign _043_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *) _006_;
  assign _044_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *) _007_;
  assign _045_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *) _033_;
  assign _046_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *) _067_;
  assign _047_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _034_;
  assign _048_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _008_;
  assign _049_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _035_;
  assign _050_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _069_;
  assign _051_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) _036_;
  assign _052_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) _010_;
  assign _053_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) _011_;
  assign _054_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) _012_;
  assign _055_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) _037_;
  assign _056_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) _071_;
  assign _057_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) _023_;
  assign _058_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) _014_;
  assign _059_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) _015_;
  assign _060_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) _016_;
  assign _061_ = ~ (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:475" *) mantissa[0];
  assign _062_ = c_h_1_5 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *) _039_;
  assign _063_ = c_h_1_9 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:463" *) _040_;
  assign _064_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_14_2_sdt_1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:465" *) _024_;
  assign _065_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_34_2_sdt_1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:467" *) _027_;
  assign _066_ = IntLeadZero_23U_leading_sign_23_0_rtn_wrs_c_56_2_sdt_1 | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:469" *) _030_;
  assign _067_ = mantissa[22] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:471" *) _045_;
  assign _068_ = mantissa[18] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _047_;
  assign _069_ = mantissa[14] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:472" *) _049_;
  assign _070_ = mantissa[10] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:473" *) _051_;
  assign _071_ = mantissa[6] | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:474" *) _055_;
  assign IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl = _017_ | (* src = "./vmod/nvdla/csc/NV_NVDLA_CSC_pra_cell.v:476" *) _020_;
  assign rtn = { c_h_1_10, IntLeadZero_23U_leading_sign_23_0_rtn_and_85_nl, IntLeadZero_23U_leading_sign_23_0_rtn_and_83_nl, IntLeadZero_23U_leading_sign_23_0_rtn_and_90_nl, IntLeadZero_23U_leading_sign_23_0_rtn_IntLeadZero_23U_leading_sign_23_0_rtn_or_2_nl };
endmodule
