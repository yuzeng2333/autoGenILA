module exp(input clk);
  reg [7:0] \buff[0] = 8'b00000000;
endmodule
