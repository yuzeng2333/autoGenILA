module bar__DOT__i1(
clk,
rst,
__ILA_bar_decode_of_i1__,
__ILA_bar_valid__,
i_wb_data,
kp,
ki,
kd,
sp,
pv,
RS,
un,
__COUNTER_start__n0
);
input            clk;
input            rst;
output            __ILA_bar_decode_of_i1__;
output            __ILA_bar_valid__;
output reg     [31:0] i_wb_data;
output reg      [1:0] kp;
output reg      [1:0] ki;
output reg      [1:0] kd;
output reg      [1:0] sp;
output reg      [1:0] pv;
output reg            RS;
output reg     [31:0] un;
output reg      [7:0] __COUNTER_start__n0;
wire            __ILA_bar_decode_of_i1__;
wire            __ILA_bar_valid__;
wire            bv_1_0_n74;
wire            bv_1_1_n2;
wire            clk;
wire            n1;
wire            n10;
wire            n100;
wire            n1000;
wire            n1001;
wire            n1002;
wire            n1003;
wire            n1004;
wire            n1005;
wire            n1006;
wire            n1007;
wire            n1008;
wire            n1009;
wire            n101;
wire            n1010;
wire            n1011;
wire            n1012;
wire            n1013;
wire            n1014;
wire            n1015;
wire            n1016;
wire            n1017;
wire            n1018;
wire            n1019;
wire            n102;
wire            n1020;
wire            n1021;
wire            n1022;
wire            n1023;
wire            n1024;
wire            n1025;
wire            n1026;
wire            n1027;
wire            n1028;
wire            n1029;
wire            n103;
wire            n1030;
wire            n1031;
wire            n1032;
wire            n1033;
wire            n1034;
wire            n1035;
wire            n1036;
wire            n1037;
wire            n1038;
wire            n1039;
wire            n104;
wire            n1040;
wire            n1041;
wire            n1042;
wire            n1043;
wire            n1044;
wire            n1045;
wire            n1046;
wire            n1047;
wire            n1048;
wire            n1049;
wire            n105;
wire            n1050;
wire            n1051;
wire            n1052;
wire            n1053;
wire            n1054;
wire            n1055;
wire            n1056;
wire            n1057;
wire            n1058;
wire            n1059;
wire            n106;
wire            n1060;
wire            n1061;
wire            n1062;
wire            n1063;
wire            n1064;
wire            n1065;
wire            n1066;
wire            n1067;
wire            n1068;
wire            n1069;
wire            n107;
wire            n1070;
wire            n1071;
wire            n1072;
wire            n1073;
wire            n1074;
wire            n1075;
wire            n1076;
wire            n1077;
wire            n1078;
wire            n1079;
wire            n108;
wire            n1080;
wire            n1081;
wire            n1082;
wire            n1083;
wire            n1084;
wire            n1085;
wire            n1086;
wire            n1087;
wire            n1088;
wire            n1089;
wire            n109;
wire            n1090;
wire            n1091;
wire            n1092;
wire            n1093;
wire            n1094;
wire            n1095;
wire            n1096;
wire            n1097;
wire            n1098;
wire            n1099;
wire            n11;
wire            n110;
wire            n1100;
wire            n1101;
wire            n1102;
wire            n1103;
wire            n1104;
wire            n1105;
wire            n1106;
wire            n1107;
wire            n1108;
wire            n1109;
wire            n111;
wire            n1110;
wire            n1111;
wire            n1112;
wire            n1113;
wire            n1114;
wire            n1115;
wire            n1116;
wire            n1117;
wire            n1118;
wire            n1119;
wire            n112;
wire            n1120;
wire            n1121;
wire            n1122;
wire            n1123;
wire            n1124;
wire            n1125;
wire            n1126;
wire            n1127;
wire            n1128;
wire            n1129;
wire            n113;
wire            n1130;
wire            n1131;
wire            n1132;
wire            n1133;
wire            n1134;
wire            n1135;
wire            n1136;
wire            n1137;
wire            n1138;
wire            n1139;
wire            n114;
wire            n1140;
wire            n1141;
wire            n1142;
wire            n1143;
wire            n1144;
wire            n1145;
wire            n1146;
wire            n1147;
wire            n1148;
wire            n1149;
wire            n115;
wire            n1150;
wire            n1151;
wire            n1152;
wire            n1153;
wire            n1154;
wire            n1155;
wire            n1156;
wire            n1157;
wire            n1158;
wire            n1159;
wire            n116;
wire            n1160;
wire            n1161;
wire            n1162;
wire            n1163;
wire            n1164;
wire            n1165;
wire            n1166;
wire            n1167;
wire            n1168;
wire            n1169;
wire            n117;
wire            n1170;
wire            n1171;
wire            n1172;
wire            n1173;
wire            n1174;
wire            n1175;
wire            n1176;
wire            n1177;
wire            n1178;
wire            n1179;
wire            n118;
wire            n1180;
wire            n1181;
wire            n1182;
wire            n1183;
wire            n1184;
wire            n1185;
wire            n1186;
wire            n1187;
wire            n1188;
wire            n1189;
wire            n119;
wire            n1190;
wire            n1191;
wire            n1192;
wire            n1193;
wire            n1194;
wire            n1195;
wire            n1196;
wire            n1197;
wire            n1198;
wire            n1199;
wire            n12;
wire            n120;
wire            n1200;
wire            n1201;
wire            n1202;
wire            n1203;
wire            n1204;
wire            n1205;
wire            n1206;
wire            n1207;
wire            n1208;
wire            n1209;
wire            n121;
wire            n1210;
wire            n1211;
wire            n1212;
wire            n1213;
wire            n1214;
wire            n1215;
wire            n1216;
wire            n1217;
wire            n1218;
wire            n1219;
wire            n122;
wire            n1220;
wire            n1221;
wire            n1222;
wire            n1223;
wire            n1224;
wire            n1225;
wire            n1226;
wire            n1227;
wire            n1228;
wire            n1229;
wire            n123;
wire            n1230;
wire            n1231;
wire            n1232;
wire            n1233;
wire            n1234;
wire            n1235;
wire            n1236;
wire            n1237;
wire            n1238;
wire            n1239;
wire            n124;
wire            n1240;
wire            n1241;
wire            n1242;
wire            n1243;
wire            n1244;
wire            n1245;
wire            n1246;
wire            n1247;
wire            n1248;
wire            n1249;
wire            n125;
wire            n1250;
wire            n1251;
wire            n1252;
wire            n1253;
wire            n1254;
wire            n1255;
wire            n1256;
wire            n1257;
wire            n1258;
wire            n1259;
wire            n126;
wire            n1260;
wire            n1261;
wire            n1262;
wire            n1263;
wire            n1264;
wire            n1265;
wire            n1266;
wire            n1267;
wire            n1268;
wire            n1269;
wire            n127;
wire            n1270;
wire            n1271;
wire            n1272;
wire            n1273;
wire            n1274;
wire            n1275;
wire            n1276;
wire            n1277;
wire            n1278;
wire            n1279;
wire            n128;
wire            n1280;
wire            n1281;
wire            n1282;
wire            n1283;
wire            n1284;
wire            n1285;
wire            n1286;
wire            n1287;
wire            n1288;
wire            n1289;
wire            n129;
wire            n1290;
wire            n1291;
wire            n1292;
wire            n1293;
wire            n1294;
wire            n1295;
wire            n1296;
wire            n1297;
wire            n1298;
wire            n1299;
wire            n13;
wire            n130;
wire            n1300;
wire            n1301;
wire            n1302;
wire            n1303;
wire            n1304;
wire            n1305;
wire            n1306;
wire            n1307;
wire            n1308;
wire            n1309;
wire            n131;
wire            n1310;
wire            n1311;
wire            n1312;
wire            n1313;
wire            n1314;
wire            n1315;
wire            n1316;
wire            n1317;
wire            n1318;
wire            n1319;
wire            n132;
wire            n1320;
wire            n1321;
wire            n1322;
wire            n1323;
wire            n1324;
wire            n1325;
wire            n1326;
wire            n1327;
wire            n1328;
wire            n1329;
wire            n133;
wire            n1330;
wire            n1331;
wire            n1332;
wire            n1333;
wire            n1334;
wire            n1335;
wire            n1336;
wire            n1337;
wire            n1338;
wire            n1339;
wire            n134;
wire            n1340;
wire            n1341;
wire            n1342;
wire            n1343;
wire            n1344;
wire            n1345;
wire            n1346;
wire            n1347;
wire            n1348;
wire            n1349;
wire            n135;
wire            n1350;
wire            n1351;
wire            n1352;
wire            n1353;
wire            n1354;
wire            n1355;
wire            n1356;
wire            n1357;
wire            n1358;
wire            n1359;
wire            n136;
wire            n1360;
wire            n1361;
wire            n1362;
wire            n1363;
wire            n1364;
wire            n1365;
wire            n1366;
wire            n1367;
wire            n1368;
wire            n1369;
wire            n137;
wire            n1370;
wire            n1371;
wire            n1372;
wire            n1373;
wire            n1374;
wire            n1375;
wire            n1376;
wire            n1377;
wire            n1378;
wire            n1379;
wire            n138;
wire            n1380;
wire            n1381;
wire            n1382;
wire            n1383;
wire            n1384;
wire            n1385;
wire            n1386;
wire            n1387;
wire            n1388;
wire            n1389;
wire            n139;
wire            n1390;
wire            n1391;
wire            n1392;
wire            n1393;
wire            n1394;
wire            n1395;
wire            n1396;
wire            n1397;
wire            n1398;
wire            n1399;
wire            n14;
wire            n140;
wire            n1400;
wire            n1401;
wire            n1402;
wire            n1403;
wire            n1404;
wire            n1405;
wire            n1406;
wire            n1407;
wire            n1408;
wire            n1409;
wire            n141;
wire            n1410;
wire            n1411;
wire            n1412;
wire            n1413;
wire            n1414;
wire            n1415;
wire            n1416;
wire            n1417;
wire            n1418;
wire            n1419;
wire            n142;
wire            n1420;
wire            n1421;
wire            n1422;
wire            n1423;
wire            n1424;
wire            n1425;
wire            n1426;
wire            n1427;
wire            n1428;
wire            n1429;
wire            n143;
wire            n1430;
wire            n1431;
wire            n1432;
wire            n1433;
wire            n1434;
wire            n1435;
wire            n1436;
wire            n1437;
wire            n1438;
wire            n1439;
wire            n144;
wire            n1440;
wire            n1441;
wire            n1442;
wire            n1443;
wire            n1444;
wire            n1445;
wire            n1446;
wire            n1447;
wire            n1448;
wire            n1449;
wire            n145;
wire            n1450;
wire            n1451;
wire            n1452;
wire            n1453;
wire            n1454;
wire            n1455;
wire            n1456;
wire            n1457;
wire            n1458;
wire            n1459;
wire            n146;
wire            n1460;
wire            n1461;
wire            n1462;
wire            n1463;
wire            n1464;
wire            n1465;
wire            n1466;
wire            n1467;
wire            n1468;
wire            n1469;
wire            n147;
wire            n1470;
wire            n1471;
wire            n1472;
wire            n1473;
wire            n1474;
wire            n1475;
wire            n1476;
wire            n1477;
wire            n1478;
wire            n1479;
wire            n148;
wire            n1480;
wire            n1481;
wire            n1482;
wire            n1483;
wire            n1484;
wire            n1485;
wire            n1486;
wire            n1487;
wire            n1488;
wire            n1489;
wire            n149;
wire            n1490;
wire            n1491;
wire            n1492;
wire            n1493;
wire            n1494;
wire            n1495;
wire            n1496;
wire            n1497;
wire            n1498;
wire            n1499;
wire            n15;
wire            n150;
wire            n1500;
wire            n1501;
wire            n1502;
wire            n1503;
wire            n1504;
wire            n1505;
wire            n1506;
wire            n1507;
wire            n1508;
wire            n1509;
wire            n151;
wire            n1510;
wire            n1511;
wire            n1512;
wire            n1513;
wire            n1514;
wire            n1515;
wire            n1516;
wire            n1517;
wire            n1518;
wire            n1519;
wire            n152;
wire            n1520;
wire            n1521;
wire            n1522;
wire            n1523;
wire            n1524;
wire            n1525;
wire            n1526;
wire            n1527;
wire            n1528;
wire            n1529;
wire            n153;
wire            n1530;
wire            n1531;
wire            n1532;
wire            n1533;
wire            n1534;
wire            n1535;
wire            n1536;
wire            n1537;
wire            n1538;
wire            n1539;
wire            n154;
wire            n1540;
wire            n1541;
wire            n1542;
wire            n1543;
wire            n1544;
wire            n1545;
wire            n1546;
wire            n1547;
wire            n1548;
wire            n1549;
wire            n155;
wire            n1550;
wire            n1551;
wire            n1552;
wire            n1553;
wire            n1554;
wire            n1555;
wire            n1556;
wire            n1557;
wire            n1558;
wire            n1559;
wire            n156;
wire            n1560;
wire            n1561;
wire            n1562;
wire            n1563;
wire            n1564;
wire            n1565;
wire            n1566;
wire            n1567;
wire            n1568;
wire            n1569;
wire            n157;
wire            n1570;
wire            n1571;
wire            n1572;
wire            n1573;
wire            n1574;
wire            n1575;
wire            n1576;
wire            n1577;
wire            n1578;
wire            n1579;
wire            n158;
wire            n1580;
wire            n1581;
wire            n1582;
wire            n1583;
wire            n1584;
wire            n1585;
wire            n1586;
wire            n1587;
wire            n1588;
wire            n1589;
wire            n159;
wire            n1590;
wire            n1591;
wire            n1592;
wire            n1593;
wire            n1594;
wire            n1595;
wire            n1596;
wire            n1597;
wire            n1598;
wire            n1599;
wire            n16;
wire            n160;
wire            n1600;
wire            n1601;
wire            n1602;
wire            n1603;
wire            n1604;
wire            n1605;
wire            n1606;
wire            n1607;
wire            n1608;
wire            n1609;
wire            n161;
wire            n1610;
wire            n1611;
wire            n1612;
wire            n1613;
wire            n1614;
wire            n1615;
wire            n1616;
wire            n1617;
wire            n1618;
wire            n1619;
wire            n162;
wire            n1620;
wire            n1621;
wire            n1622;
wire            n1623;
wire            n1624;
wire            n1625;
wire            n1626;
wire            n1627;
wire            n1628;
wire            n1629;
wire            n163;
wire            n1630;
wire            n1631;
wire            n1632;
wire            n1633;
wire            n1634;
wire            n1635;
wire            n1636;
wire            n1637;
wire            n1638;
wire            n1639;
wire            n164;
wire            n1640;
wire            n1641;
wire            n1642;
wire            n1643;
wire            n1644;
wire            n1645;
wire            n1646;
wire            n1647;
wire            n1648;
wire            n1649;
wire            n165;
wire            n1650;
wire            n1651;
wire            n1652;
wire            n1653;
wire            n1654;
wire            n1655;
wire            n1656;
wire            n1657;
wire            n1658;
wire            n1659;
wire            n166;
wire            n1660;
wire            n1661;
wire            n1662;
wire            n1663;
wire            n1664;
wire            n1665;
wire            n1666;
wire            n1667;
wire            n1668;
wire            n1669;
wire            n167;
wire            n1670;
wire            n1671;
wire            n1672;
wire            n1673;
wire            n1674;
wire            n1675;
wire            n1676;
wire            n1677;
wire            n1678;
wire            n1679;
wire            n168;
wire            n1680;
wire            n1681;
wire            n1682;
wire            n1683;
wire            n1684;
wire            n1685;
wire            n1686;
wire            n1687;
wire            n1688;
wire            n1689;
wire            n169;
wire            n1690;
wire            n1691;
wire            n1692;
wire            n1693;
wire            n1694;
wire            n1695;
wire            n1696;
wire            n1697;
wire            n1698;
wire            n1699;
wire            n17;
wire            n170;
wire            n1700;
wire            n1701;
wire            n1702;
wire            n1703;
wire            n1704;
wire            n1705;
wire            n1706;
wire            n1707;
wire            n1708;
wire            n1709;
wire            n171;
wire            n1710;
wire            n1711;
wire            n1712;
wire            n1713;
wire            n1714;
wire            n1715;
wire            n1716;
wire            n1717;
wire            n1718;
wire            n1719;
wire            n172;
wire            n1720;
wire            n1721;
wire            n1722;
wire            n1723;
wire            n1724;
wire            n1725;
wire            n1726;
wire            n1727;
wire            n1728;
wire            n1729;
wire            n173;
wire            n1730;
wire            n1731;
wire            n1732;
wire            n1733;
wire            n1734;
wire            n1735;
wire            n1736;
wire            n1737;
wire            n1738;
wire            n1739;
wire            n174;
wire            n1740;
wire            n1741;
wire            n1742;
wire            n1743;
wire            n1744;
wire            n1745;
wire            n1746;
wire            n1747;
wire            n1748;
wire            n1749;
wire            n175;
wire            n1750;
wire            n1751;
wire            n1752;
wire            n1753;
wire            n1754;
wire            n1755;
wire            n1756;
wire            n1757;
wire            n1758;
wire            n1759;
wire            n176;
wire            n1760;
wire            n1761;
wire            n1762;
wire            n1763;
wire            n1764;
wire            n1765;
wire            n1766;
wire            n1767;
wire            n1768;
wire            n1769;
wire            n177;
wire            n1770;
wire            n1771;
wire            n1772;
wire            n1773;
wire            n1774;
wire            n1775;
wire            n1776;
wire            n1777;
wire            n1778;
wire            n1779;
wire            n178;
wire            n1780;
wire            n1781;
wire            n1782;
wire            n1783;
wire            n1784;
wire            n1785;
wire            n1786;
wire            n1787;
wire            n1788;
wire            n1789;
wire            n179;
wire            n1790;
wire            n1791;
wire            n1792;
wire            n1793;
wire            n1794;
wire            n1795;
wire            n1796;
wire            n1797;
wire            n1798;
wire            n1799;
wire            n18;
wire            n180;
wire            n1800;
wire            n1801;
wire            n1802;
wire            n1803;
wire            n1804;
wire            n1805;
wire            n1806;
wire            n1807;
wire            n1808;
wire            n1809;
wire            n181;
wire            n1810;
wire            n1811;
wire            n1812;
wire            n1813;
wire            n1814;
wire            n1815;
wire            n1816;
wire            n1817;
wire            n1818;
wire            n1819;
wire            n182;
wire            n1820;
wire            n1821;
wire            n1822;
wire            n1823;
wire            n1824;
wire            n1825;
wire            n1826;
wire            n1827;
wire            n1828;
wire            n1829;
wire            n183;
wire            n1830;
wire            n1831;
wire            n1832;
wire            n1833;
wire            n1834;
wire            n1835;
wire            n1836;
wire            n1837;
wire            n1838;
wire            n1839;
wire            n184;
wire            n1840;
wire            n1841;
wire            n1842;
wire            n1843;
wire            n1844;
wire            n1845;
wire            n1846;
wire            n1847;
wire            n1848;
wire            n1849;
wire            n185;
wire            n1850;
wire            n1851;
wire            n1852;
wire            n1853;
wire            n1854;
wire            n1855;
wire            n1856;
wire            n1857;
wire            n1858;
wire            n1859;
wire            n186;
wire            n1860;
wire            n1861;
wire            n1862;
wire            n1863;
wire            n1864;
wire            n1865;
wire            n1866;
wire            n1867;
wire            n1868;
wire            n1869;
wire            n187;
wire            n1870;
wire            n1871;
wire            n1872;
wire            n1873;
wire            n1874;
wire            n1875;
wire            n1876;
wire            n1877;
wire            n1878;
wire            n1879;
wire            n188;
wire            n1880;
wire            n1881;
wire            n1882;
wire            n1883;
wire            n1884;
wire            n1885;
wire            n1886;
wire            n1887;
wire            n1888;
wire            n1889;
wire            n189;
wire            n1890;
wire            n1891;
wire            n1892;
wire            n1893;
wire            n1894;
wire            n1895;
wire            n1896;
wire            n1897;
wire            n1898;
wire            n1899;
wire            n19;
wire            n190;
wire            n1900;
wire            n1901;
wire            n1902;
wire            n1903;
wire            n1904;
wire            n1905;
wire            n1906;
wire            n1907;
wire            n1908;
wire            n1909;
wire            n191;
wire            n1910;
wire            n1911;
wire            n1912;
wire            n1913;
wire            n1914;
wire            n1915;
wire            n1916;
wire            n1917;
wire            n1918;
wire            n1919;
wire            n192;
wire            n1920;
wire            n1921;
wire            n1922;
wire            n1923;
wire            n1924;
wire            n1925;
wire            n1926;
wire            n1927;
wire            n1928;
wire            n1929;
wire            n193;
wire            n1930;
wire            n1931;
wire            n1932;
wire            n1933;
wire            n1934;
wire            n1935;
wire            n1936;
wire            n1937;
wire            n1938;
wire            n1939;
wire            n194;
wire            n1940;
wire            n1941;
wire            n1942;
wire            n1943;
wire            n1944;
wire            n1945;
wire            n1946;
wire            n1947;
wire            n1948;
wire            n1949;
wire            n195;
wire            n1950;
wire            n1951;
wire            n1952;
wire            n1953;
wire            n1954;
wire            n1955;
wire            n1956;
wire            n1957;
wire            n1958;
wire            n1959;
wire            n196;
wire            n1960;
wire            n1961;
wire            n1962;
wire            n1963;
wire            n1964;
wire            n1965;
wire            n1966;
wire            n1967;
wire            n1968;
wire            n1969;
wire            n197;
wire            n1970;
wire            n1971;
wire            n1972;
wire            n1973;
wire            n1974;
wire            n1975;
wire            n1976;
wire            n1977;
wire            n1978;
wire            n1979;
wire            n198;
wire            n1980;
wire            n1981;
wire            n1982;
wire            n1983;
wire            n1984;
wire            n1985;
wire            n1986;
wire            n1987;
wire            n1988;
wire            n1989;
wire            n199;
wire            n1990;
wire            n1991;
wire            n1992;
wire            n1993;
wire            n1994;
wire            n1995;
wire            n1996;
wire            n1997;
wire            n1998;
wire            n1999;
wire            n20;
wire            n200;
wire            n2000;
wire            n2001;
wire            n2002;
wire            n2003;
wire            n2004;
wire            n2005;
wire            n2006;
wire            n2007;
wire            n2008;
wire            n2009;
wire            n201;
wire            n2010;
wire            n2011;
wire            n2012;
wire            n2013;
wire            n2014;
wire            n2015;
wire            n2016;
wire            n2017;
wire            n2018;
wire            n2019;
wire            n202;
wire            n2020;
wire            n2021;
wire            n2022;
wire            n2023;
wire            n2024;
wire            n2025;
wire            n2026;
wire            n2027;
wire            n2028;
wire            n2029;
wire            n203;
wire            n2030;
wire            n2031;
wire            n2032;
wire            n2033;
wire            n2034;
wire            n2035;
wire            n2036;
wire            n2037;
wire            n2038;
wire            n2039;
wire            n204;
wire            n2040;
wire            n2041;
wire            n2042;
wire            n2043;
wire            n2044;
wire            n2045;
wire            n2046;
wire            n2047;
wire            n2048;
wire            n2049;
wire            n205;
wire            n2050;
wire            n2051;
wire            n2052;
wire            n2053;
wire            n2054;
wire            n2055;
wire            n2056;
wire            n2057;
wire            n2058;
wire            n2059;
wire            n206;
wire            n2060;
wire            n2061;
wire            n2062;
wire            n2063;
wire            n2064;
wire            n2065;
wire            n2066;
wire            n2067;
wire            n2068;
wire            n2069;
wire            n207;
wire            n2070;
wire            n2071;
wire            n2072;
wire            n2073;
wire            n2074;
wire            n2075;
wire            n2076;
wire            n2077;
wire            n2078;
wire            n2079;
wire            n208;
wire            n2080;
wire            n2081;
wire            n2082;
wire            n2083;
wire            n2084;
wire            n2085;
wire            n2086;
wire            n2087;
wire            n2088;
wire            n2089;
wire            n209;
wire            n2090;
wire            n2091;
wire            n2092;
wire            n2093;
wire            n2094;
wire            n2095;
wire            n2096;
wire            n2097;
wire            n2098;
wire            n2099;
wire            n21;
wire            n210;
wire            n2100;
wire            n2101;
wire            n2102;
wire            n2103;
wire            n2104;
wire            n2105;
wire            n2106;
wire            n2107;
wire            n2108;
wire            n2109;
wire            n211;
wire            n2110;
wire            n2111;
wire            n2112;
wire            n2113;
wire            n2114;
wire            n2115;
wire            n2116;
wire            n2117;
wire            n2118;
wire            n2119;
wire            n212;
wire            n2120;
wire            n2121;
wire            n2122;
wire            n2123;
wire            n2124;
wire            n2125;
wire            n2126;
wire            n2127;
wire            n2128;
wire            n2129;
wire            n213;
wire            n2130;
wire            n2131;
wire            n2132;
wire            n2133;
wire            n2134;
wire            n2135;
wire            n2136;
wire            n2137;
wire            n2138;
wire            n2139;
wire            n214;
wire            n2140;
wire            n2141;
wire            n2142;
wire            n2143;
wire            n2144;
wire            n2145;
wire            n2146;
wire            n2147;
wire            n2148;
wire            n2149;
wire            n215;
wire            n2150;
wire            n2151;
wire            n2152;
wire            n2153;
wire            n2154;
wire            n2155;
wire            n2156;
wire            n2157;
wire            n2158;
wire            n2159;
wire            n216;
wire            n2160;
wire            n2161;
wire            n2162;
wire            n2163;
wire            n2164;
wire            n2165;
wire            n2166;
wire            n2167;
wire            n2168;
wire            n2169;
wire            n217;
wire            n2170;
wire            n2171;
wire            n2172;
wire            n2173;
wire            n2174;
wire            n2175;
wire            n2176;
wire            n2177;
wire            n2178;
wire            n2179;
wire            n218;
wire            n2180;
wire            n2181;
wire            n2182;
wire            n2183;
wire            n2184;
wire            n2185;
wire            n2186;
wire            n2187;
wire            n2188;
wire            n2189;
wire            n219;
wire            n2190;
wire            n2191;
wire            n2192;
wire            n2193;
wire            n2194;
wire            n2195;
wire            n2196;
wire            n2197;
wire            n2198;
wire            n2199;
wire            n22;
wire            n220;
wire            n2200;
wire            n2201;
wire            n2202;
wire            n2203;
wire            n2204;
wire            n2205;
wire            n2206;
wire            n2207;
wire            n2208;
wire            n2209;
wire            n221;
wire            n2210;
wire            n2211;
wire            n2212;
wire            n2213;
wire            n2214;
wire            n2215;
wire            n2216;
wire            n2217;
wire            n2218;
wire            n2219;
wire            n222;
wire            n2220;
wire            n2221;
wire            n2222;
wire            n2223;
wire            n2224;
wire            n2225;
wire            n2226;
wire            n2227;
wire            n2228;
wire            n2229;
wire            n223;
wire            n2230;
wire            n2231;
wire            n2232;
wire            n2233;
wire            n2234;
wire            n2235;
wire            n2236;
wire            n2237;
wire            n2238;
wire            n2239;
wire            n224;
wire            n2240;
wire            n2241;
wire            n2242;
wire            n2243;
wire            n2244;
wire            n2245;
wire            n2246;
wire            n2247;
wire            n2248;
wire            n2249;
wire            n225;
wire            n2250;
wire            n2251;
wire            n2252;
wire            n2253;
wire            n2254;
wire            n2255;
wire            n2256;
wire            n2257;
wire            n2258;
wire            n2259;
wire            n226;
wire            n2260;
wire            n2261;
wire            n2262;
wire            n2263;
wire            n2264;
wire            n2265;
wire            n2266;
wire            n2267;
wire            n2268;
wire            n2269;
wire            n227;
wire            n2270;
wire            n2271;
wire            n2272;
wire            n2273;
wire            n2274;
wire            n2275;
wire            n2276;
wire            n2277;
wire            n2278;
wire            n2279;
wire            n228;
wire            n2280;
wire            n2281;
wire            n2282;
wire            n2283;
wire            n2284;
wire            n2285;
wire            n2286;
wire            n2287;
wire            n2288;
wire            n2289;
wire            n229;
wire            n2290;
wire            n2291;
wire            n2292;
wire            n2293;
wire            n2294;
wire            n2295;
wire            n2296;
wire            n2297;
wire            n2298;
wire            n2299;
wire            n23;
wire            n230;
wire            n2300;
wire            n2301;
wire            n2302;
wire            n2303;
wire            n2304;
wire            n2305;
wire            n2306;
wire            n2307;
wire            n2308;
wire            n2309;
wire            n231;
wire            n2310;
wire            n2311;
wire            n2312;
wire            n2313;
wire            n2314;
wire            n2315;
wire            n2316;
wire            n2317;
wire            n2318;
wire            n2319;
wire            n232;
wire            n2320;
wire            n2321;
wire            n2322;
wire            n2323;
wire            n2324;
wire            n2325;
wire            n2326;
wire            n2327;
wire            n2328;
wire            n2329;
wire            n233;
wire            n2330;
wire            n2331;
wire            n2332;
wire            n2333;
wire            n2334;
wire            n2335;
wire            n2336;
wire            n2337;
wire            n2338;
wire            n2339;
wire            n234;
wire            n2340;
wire            n2341;
wire            n2342;
wire            n2343;
wire            n2344;
wire            n2345;
wire            n2346;
wire            n2347;
wire            n2348;
wire            n2349;
wire            n235;
wire            n2350;
wire            n2351;
wire            n2352;
wire            n2353;
wire            n2354;
wire            n2355;
wire            n2356;
wire            n2357;
wire            n2358;
wire            n2359;
wire            n236;
wire            n2360;
wire            n2361;
wire            n2362;
wire            n2363;
wire            n2364;
wire            n2365;
wire            n2366;
wire            n2367;
wire            n2368;
wire            n2369;
wire            n237;
wire            n2370;
wire            n2371;
wire            n2372;
wire            n2373;
wire            n2374;
wire            n2375;
wire            n2376;
wire            n2377;
wire            n2378;
wire            n2379;
wire            n238;
wire            n2380;
wire            n2381;
wire            n2382;
wire            n2383;
wire            n2384;
wire            n2385;
wire            n2386;
wire            n2387;
wire            n2388;
wire            n2389;
wire            n239;
wire            n2390;
wire            n2391;
wire            n2392;
wire            n2393;
wire            n2394;
wire            n2395;
wire            n2396;
wire            n2397;
wire            n2398;
wire            n2399;
wire            n24;
wire            n240;
wire            n2400;
wire            n2401;
wire            n2402;
wire            n2403;
wire            n2404;
wire            n2405;
wire            n2406;
wire            n2407;
wire            n2408;
wire            n2409;
wire            n241;
wire            n2410;
wire            n2411;
wire            n2412;
wire            n2413;
wire            n2414;
wire            n2415;
wire            n2416;
wire            n2417;
wire            n2418;
wire            n2419;
wire            n242;
wire            n2420;
wire            n2421;
wire            n2422;
wire            n2423;
wire            n2424;
wire            n2425;
wire            n2426;
wire            n2427;
wire            n2428;
wire            n2429;
wire            n243;
wire            n2430;
wire            n2431;
wire            n2432;
wire            n2433;
wire            n2434;
wire            n2435;
wire            n2436;
wire            n2437;
wire            n2438;
wire            n2439;
wire            n244;
wire            n2440;
wire            n2441;
wire            n2442;
wire            n2443;
wire            n2444;
wire            n2445;
wire            n2446;
wire            n2447;
wire            n2448;
wire            n2449;
wire            n245;
wire            n2450;
wire            n2451;
wire            n2452;
wire            n2453;
wire            n2454;
wire            n2455;
wire            n2456;
wire            n2457;
wire            n2458;
wire            n2459;
wire            n246;
wire            n2460;
wire            n2461;
wire            n2462;
wire            n2463;
wire            n2464;
wire            n2465;
wire            n2466;
wire            n2467;
wire            n2468;
wire            n2469;
wire            n247;
wire            n2470;
wire            n2471;
wire            n2472;
wire            n2473;
wire            n2474;
wire            n2475;
wire            n2476;
wire            n2477;
wire            n2478;
wire            n2479;
wire            n248;
wire            n2480;
wire            n2481;
wire            n2482;
wire            n2483;
wire            n2484;
wire            n2485;
wire            n2486;
wire            n2487;
wire            n2488;
wire            n2489;
wire            n249;
wire            n2490;
wire            n2491;
wire            n2492;
wire            n2493;
wire            n2494;
wire            n2495;
wire            n2496;
wire            n2497;
wire            n2498;
wire            n2499;
wire            n25;
wire            n250;
wire            n2500;
wire            n2501;
wire            n2502;
wire            n2503;
wire            n2504;
wire            n2505;
wire            n2506;
wire            n2507;
wire            n2508;
wire            n2509;
wire            n251;
wire            n2510;
wire            n2511;
wire            n2512;
wire            n2513;
wire            n2514;
wire            n2515;
wire            n2516;
wire            n2517;
wire            n2518;
wire            n2519;
wire            n252;
wire            n2520;
wire            n2521;
wire            n2522;
wire            n2523;
wire            n2524;
wire            n2525;
wire            n2526;
wire            n2527;
wire            n2528;
wire            n2529;
wire            n253;
wire            n2530;
wire            n2531;
wire            n2532;
wire            n2533;
wire            n2534;
wire            n2535;
wire            n2536;
wire            n2537;
wire            n2538;
wire            n2539;
wire            n254;
wire            n2540;
wire            n2541;
wire            n2542;
wire            n2543;
wire            n2544;
wire            n2545;
wire            n2546;
wire            n2547;
wire            n2548;
wire            n2549;
wire            n255;
wire            n2550;
wire            n2551;
wire            n2552;
wire            n2553;
wire            n2554;
wire            n2555;
wire            n2556;
wire            n2557;
wire            n2558;
wire            n2559;
wire            n256;
wire            n2560;
wire            n2561;
wire            n2562;
wire            n2563;
wire            n2564;
wire            n2565;
wire            n2566;
wire            n2567;
wire            n2568;
wire            n2569;
wire            n257;
wire            n2570;
wire            n2571;
wire            n2572;
wire            n2573;
wire            n2574;
wire            n2575;
wire            n2576;
wire            n2577;
wire            n2578;
wire            n2579;
wire            n258;
wire            n2580;
wire            n2581;
wire            n2582;
wire            n2583;
wire            n2584;
wire            n2585;
wire            n2586;
wire            n2587;
wire            n2588;
wire            n2589;
wire            n259;
wire            n2590;
wire            n2591;
wire            n2592;
wire            n2593;
wire            n2594;
wire            n2595;
wire            n2596;
wire            n2597;
wire            n2598;
wire            n2599;
wire            n26;
wire            n260;
wire            n2600;
wire            n2601;
wire            n2602;
wire            n2603;
wire            n2604;
wire            n2605;
wire            n2606;
wire            n2607;
wire            n2608;
wire            n2609;
wire            n261;
wire            n2610;
wire            n2611;
wire            n2612;
wire            n2613;
wire            n2614;
wire            n2615;
wire            n2616;
wire            n2617;
wire            n2618;
wire            n2619;
wire            n262;
wire            n2620;
wire            n2621;
wire            n2622;
wire            n2623;
wire            n2624;
wire            n2625;
wire            n2626;
wire            n2627;
wire            n2628;
wire            n2629;
wire            n263;
wire            n2630;
wire            n2631;
wire            n2632;
wire            n2633;
wire            n2634;
wire            n2635;
wire            n2636;
wire            n2637;
wire            n2638;
wire            n2639;
wire            n264;
wire            n2640;
wire            n2641;
wire            n2642;
wire            n2643;
wire            n2644;
wire            n2645;
wire            n2646;
wire            n2647;
wire            n2648;
wire            n2649;
wire            n265;
wire            n2650;
wire            n2651;
wire            n2652;
wire            n2653;
wire            n2654;
wire            n2655;
wire            n2656;
wire            n2657;
wire            n2658;
wire            n2659;
wire            n266;
wire            n2660;
wire            n2661;
wire            n2662;
wire            n2663;
wire            n2664;
wire            n2665;
wire            n2666;
wire            n2667;
wire            n2668;
wire            n2669;
wire            n267;
wire            n2670;
wire            n2671;
wire            n2672;
wire            n2673;
wire            n2674;
wire            n2675;
wire            n2676;
wire            n2677;
wire            n2678;
wire            n2679;
wire            n268;
wire            n2680;
wire            n2681;
wire            n2682;
wire            n2683;
wire            n2684;
wire            n2685;
wire            n2686;
wire            n2687;
wire            n2688;
wire            n2689;
wire            n269;
wire            n2690;
wire            n2691;
wire            n2692;
wire            n2693;
wire            n2694;
wire            n2695;
wire            n2696;
wire            n2697;
wire            n2698;
wire            n2699;
wire            n27;
wire            n270;
wire            n2700;
wire            n2701;
wire            n2702;
wire            n2703;
wire            n2704;
wire            n2705;
wire            n2706;
wire            n2707;
wire            n2708;
wire            n2709;
wire            n271;
wire            n2710;
wire            n2711;
wire            n2712;
wire            n2713;
wire            n2714;
wire            n2715;
wire            n2716;
wire            n2717;
wire            n2718;
wire            n2719;
wire            n272;
wire            n2720;
wire            n2721;
wire            n2722;
wire            n2723;
wire            n2724;
wire            n2725;
wire            n2726;
wire            n2727;
wire            n2728;
wire            n2729;
wire            n273;
wire            n2730;
wire            n2731;
wire            n2732;
wire            n2733;
wire            n2734;
wire            n2735;
wire            n2736;
wire            n2737;
wire            n2738;
wire            n2739;
wire            n274;
wire            n2740;
wire            n2741;
wire            n2742;
wire            n2743;
wire            n2744;
wire            n2745;
wire            n2746;
wire            n2747;
wire            n2748;
wire            n2749;
wire            n275;
wire            n2750;
wire            n2751;
wire            n2752;
wire            n2753;
wire            n2754;
wire            n2755;
wire            n2756;
wire            n2757;
wire            n2758;
wire            n2759;
wire            n276;
wire            n2760;
wire            n2761;
wire            n2762;
wire            n2763;
wire            n2764;
wire            n2765;
wire            n2766;
wire            n2767;
wire            n2768;
wire            n2769;
wire            n277;
wire            n2770;
wire            n2771;
wire            n2772;
wire            n2773;
wire            n2774;
wire            n2775;
wire            n2776;
wire            n2777;
wire            n2778;
wire            n2779;
wire            n278;
wire            n2780;
wire            n2781;
wire            n2782;
wire            n2783;
wire            n2784;
wire            n2785;
wire            n2786;
wire            n2787;
wire            n2788;
wire            n2789;
wire            n279;
wire            n2790;
wire            n2791;
wire            n2792;
wire            n2793;
wire            n2794;
wire            n2795;
wire            n2796;
wire            n2797;
wire            n2798;
wire            n2799;
wire            n28;
wire            n280;
wire            n2800;
wire            n2801;
wire            n2802;
wire            n2803;
wire            n2804;
wire            n2805;
wire            n2806;
wire            n2807;
wire            n2808;
wire            n2809;
wire            n281;
wire            n2810;
wire            n2811;
wire            n2812;
wire            n2813;
wire            n2814;
wire            n2815;
wire            n2816;
wire            n2817;
wire            n2818;
wire            n2819;
wire            n282;
wire            n2820;
wire            n2821;
wire            n2822;
wire            n2823;
wire            n2824;
wire            n2825;
wire            n2826;
wire            n2827;
wire            n2828;
wire            n2829;
wire            n283;
wire            n2830;
wire            n2831;
wire            n2832;
wire            n2833;
wire            n2834;
wire            n2835;
wire            n2836;
wire            n2837;
wire            n2838;
wire            n2839;
wire            n284;
wire            n2840;
wire            n2841;
wire            n2842;
wire            n2843;
wire            n2844;
wire            n2845;
wire            n2846;
wire            n2847;
wire            n2848;
wire            n2849;
wire            n285;
wire            n2850;
wire            n2851;
wire            n2852;
wire            n2853;
wire            n2854;
wire            n2855;
wire            n2856;
wire            n2857;
wire            n2858;
wire            n2859;
wire            n286;
wire            n2860;
wire            n2861;
wire            n2862;
wire            n2863;
wire            n2864;
wire            n2865;
wire            n2866;
wire            n2867;
wire            n2868;
wire            n2869;
wire            n287;
wire            n2870;
wire            n2871;
wire            n2872;
wire            n2873;
wire            n2874;
wire            n2875;
wire            n2876;
wire            n2877;
wire            n2878;
wire            n2879;
wire            n288;
wire            n2880;
wire            n2881;
wire            n2882;
wire            n2883;
wire            n2884;
wire            n2885;
wire            n2886;
wire            n2887;
wire            n2888;
wire            n2889;
wire            n289;
wire            n2890;
wire            n2891;
wire            n2892;
wire            n2893;
wire            n2894;
wire            n2895;
wire            n2896;
wire            n2897;
wire            n2898;
wire            n2899;
wire            n29;
wire            n290;
wire            n2900;
wire            n2901;
wire            n2902;
wire            n2903;
wire            n2904;
wire            n2905;
wire            n2906;
wire            n2907;
wire            n2908;
wire            n2909;
wire            n291;
wire            n2910;
wire            n2911;
wire            n2912;
wire            n2913;
wire            n2914;
wire            n2915;
wire            n2916;
wire            n2917;
wire            n2918;
wire            n2919;
wire            n292;
wire            n2920;
wire            n2921;
wire            n2922;
wire            n2923;
wire            n2924;
wire            n2925;
wire            n2926;
wire            n2927;
wire            n2928;
wire            n2929;
wire            n293;
wire            n2930;
wire            n2931;
wire            n2932;
wire            n2933;
wire            n2934;
wire            n2935;
wire            n2936;
wire            n2937;
wire            n2938;
wire            n2939;
wire            n294;
wire            n2940;
wire            n2941;
wire            n2942;
wire            n2943;
wire            n2944;
wire            n2945;
wire            n2946;
wire            n2947;
wire            n2948;
wire            n2949;
wire            n295;
wire            n2950;
wire            n2951;
wire            n2952;
wire            n2953;
wire            n2954;
wire            n2955;
wire            n2956;
wire            n2957;
wire            n2958;
wire            n2959;
wire            n296;
wire            n2960;
wire            n2961;
wire            n2962;
wire            n2963;
wire            n2964;
wire            n2965;
wire            n2966;
wire            n2967;
wire            n2968;
wire            n2969;
wire            n297;
wire            n2970;
wire            n2971;
wire            n2972;
wire            n2973;
wire            n2974;
wire            n2975;
wire            n2976;
wire            n2977;
wire            n2978;
wire            n2979;
wire            n298;
wire            n2980;
wire            n2981;
wire            n2982;
wire            n2983;
wire            n2984;
wire            n2985;
wire            n2986;
wire            n2987;
wire            n2988;
wire            n2989;
wire            n299;
wire            n2990;
wire            n2991;
wire            n2992;
wire            n2993;
wire            n2994;
wire            n2995;
wire            n2996;
wire            n2997;
wire            n2998;
wire            n2999;
wire            n3;
wire            n30;
wire            n300;
wire            n3000;
wire            n3001;
wire            n3002;
wire            n3003;
wire            n3004;
wire            n3005;
wire            n3006;
wire            n3007;
wire            n3008;
wire            n3009;
wire            n301;
wire            n3010;
wire            n3011;
wire            n3012;
wire            n3013;
wire            n3014;
wire            n3015;
wire            n3016;
wire            n3017;
wire            n3018;
wire            n3019;
wire            n302;
wire            n3020;
wire            n3021;
wire            n3022;
wire            n3023;
wire            n3024;
wire            n3025;
wire            n3026;
wire            n3027;
wire            n3028;
wire            n3029;
wire            n303;
wire            n3030;
wire            n3031;
wire            n3032;
wire            n3033;
wire            n3034;
wire            n3035;
wire            n3036;
wire            n3037;
wire            n3038;
wire            n3039;
wire            n304;
wire            n3040;
wire            n3041;
wire            n3042;
wire            n3043;
wire            n3044;
wire            n3045;
wire            n3046;
wire            n3047;
wire            n3048;
wire            n3049;
wire            n305;
wire            n3050;
wire            n3051;
wire            n3052;
wire            n3053;
wire            n3054;
wire            n3055;
wire            n3056;
wire            n3057;
wire            n3058;
wire            n3059;
wire            n306;
wire            n3060;
wire            n3061;
wire            n3062;
wire            n3063;
wire            n3064;
wire            n3065;
wire            n3066;
wire            n3067;
wire            n3068;
wire            n3069;
wire            n307;
wire            n3070;
wire            n3071;
wire            n3072;
wire            n3073;
wire            n3074;
wire            n3075;
wire            n3076;
wire            n3077;
wire            n3078;
wire            n3079;
wire            n308;
wire            n3080;
wire            n3081;
wire            n3082;
wire            n3083;
wire            n3084;
wire            n3085;
wire            n3086;
wire            n3087;
wire            n3088;
wire            n3089;
wire            n309;
wire            n3090;
wire            n3091;
wire            n3092;
wire            n3093;
wire            n3094;
wire            n3095;
wire            n3096;
wire            n3097;
wire            n3098;
wire            n3099;
wire            n31;
wire            n310;
wire            n3100;
wire            n3101;
wire            n3102;
wire            n3103;
wire            n3104;
wire            n3105;
wire            n3106;
wire            n3107;
wire            n3108;
wire            n3109;
wire            n311;
wire            n3110;
wire            n3111;
wire            n3112;
wire            n3113;
wire            n3114;
wire            n3115;
wire            n3116;
wire            n3117;
wire            n3118;
wire            n3119;
wire            n312;
wire            n3120;
wire            n3121;
wire            n3122;
wire            n3123;
wire            n3124;
wire            n3125;
wire            n3126;
wire            n3127;
wire            n3128;
wire            n3129;
wire            n313;
wire            n3130;
wire            n3131;
wire            n3132;
wire            n3133;
wire            n3134;
wire            n3135;
wire            n3136;
wire            n3137;
wire            n3138;
wire            n3139;
wire            n314;
wire            n3140;
wire            n3141;
wire            n3142;
wire            n3143;
wire            n3144;
wire            n3145;
wire            n3146;
wire            n3147;
wire            n3148;
wire            n3149;
wire            n315;
wire            n3150;
wire            n3151;
wire            n3152;
wire            n3153;
wire            n3154;
wire            n3155;
wire            n3156;
wire            n3157;
wire            n3158;
wire            n3159;
wire            n316;
wire            n3160;
wire            n3161;
wire            n3162;
wire            n3163;
wire            n3164;
wire            n3165;
wire            n3166;
wire            n3167;
wire            n3168;
wire            n3169;
wire            n317;
wire            n3170;
wire            n3171;
wire            n3172;
wire            n3173;
wire            n3174;
wire            n3175;
wire            n3176;
wire            n3177;
wire            n3178;
wire            n3179;
wire            n318;
wire            n3180;
wire            n3181;
wire            n3182;
wire            n3183;
wire            n3184;
wire            n3185;
wire            n3186;
wire            n3187;
wire            n3188;
wire            n3189;
wire            n319;
wire            n3190;
wire            n3191;
wire            n3192;
wire            n3193;
wire            n3194;
wire            n3195;
wire            n3196;
wire            n3197;
wire            n3198;
wire            n3199;
wire            n32;
wire            n320;
wire            n3200;
wire            n3201;
wire            n3202;
wire            n3203;
wire            n3204;
wire            n3205;
wire            n3206;
wire            n3207;
wire            n3208;
wire            n3209;
wire            n321;
wire            n3210;
wire            n3211;
wire            n3212;
wire            n3213;
wire            n3214;
wire            n3215;
wire            n3216;
wire            n3217;
wire            n3218;
wire            n3219;
wire            n322;
wire            n3220;
wire            n3221;
wire            n3222;
wire            n3223;
wire            n3224;
wire            n3225;
wire            n3226;
wire            n3227;
wire            n3228;
wire            n3229;
wire            n323;
wire            n3230;
wire            n3231;
wire            n3232;
wire            n3233;
wire            n3234;
wire            n3235;
wire            n3236;
wire            n3237;
wire            n3238;
wire            n3239;
wire            n324;
wire            n3240;
wire            n3241;
wire            n3242;
wire            n3243;
wire            n3244;
wire            n3245;
wire            n3246;
wire            n3247;
wire            n3248;
wire            n3249;
wire            n325;
wire            n3250;
wire            n3251;
wire            n3252;
wire            n3253;
wire            n3254;
wire            n3255;
wire            n3256;
wire            n3257;
wire            n3258;
wire            n3259;
wire            n326;
wire            n3260;
wire            n3261;
wire            n3262;
wire            n3263;
wire            n3264;
wire            n3265;
wire            n3266;
wire            n3267;
wire            n3268;
wire            n3269;
wire            n327;
wire            n3270;
wire            n3271;
wire            n3272;
wire            n3273;
wire            n3274;
wire            n3275;
wire            n3276;
wire            n3277;
wire            n3278;
wire            n3279;
wire            n328;
wire            n3280;
wire            n3281;
wire            n3282;
wire            n3283;
wire            n3284;
wire            n3285;
wire            n3286;
wire            n3287;
wire            n3288;
wire            n3289;
wire            n329;
wire            n3290;
wire            n3291;
wire            n3292;
wire            n3293;
wire            n3294;
wire            n3295;
wire            n3296;
wire            n3297;
wire            n3298;
wire            n3299;
wire            n33;
wire            n330;
wire            n3300;
wire            n3301;
wire            n3302;
wire            n3303;
wire            n3304;
wire            n3305;
wire            n3306;
wire            n3307;
wire            n3308;
wire            n3309;
wire            n331;
wire            n3310;
wire            n3311;
wire            n3312;
wire            n3313;
wire            n3314;
wire            n3315;
wire            n3316;
wire            n3317;
wire            n3318;
wire            n3319;
wire            n332;
wire            n3320;
wire            n3321;
wire            n3322;
wire            n3323;
wire            n3324;
wire            n3325;
wire            n3326;
wire            n3327;
wire            n3328;
wire            n3329;
wire            n333;
wire            n3330;
wire            n3331;
wire            n3332;
wire            n3333;
wire            n3334;
wire            n3335;
wire            n3336;
wire            n3337;
wire            n3338;
wire            n3339;
wire            n334;
wire            n3340;
wire            n3341;
wire            n3342;
wire            n3343;
wire            n3344;
wire            n3345;
wire            n3346;
wire            n3347;
wire            n3348;
wire            n3349;
wire            n335;
wire            n3350;
wire            n3351;
wire            n3352;
wire            n3353;
wire            n3354;
wire            n3355;
wire            n3356;
wire            n3357;
wire            n3358;
wire            n3359;
wire            n336;
wire            n3360;
wire            n3361;
wire            n3362;
wire            n3363;
wire            n3364;
wire            n3365;
wire            n3366;
wire            n3367;
wire            n3368;
wire            n3369;
wire            n337;
wire            n3370;
wire            n3371;
wire            n3372;
wire            n3373;
wire            n3374;
wire            n3375;
wire            n3376;
wire            n3377;
wire            n3378;
wire            n3379;
wire            n338;
wire            n3380;
wire            n3381;
wire            n3382;
wire            n3383;
wire            n3384;
wire            n3385;
wire            n3386;
wire            n3387;
wire            n3388;
wire            n3389;
wire            n339;
wire            n3390;
wire            n3391;
wire            n3392;
wire            n3393;
wire            n3394;
wire            n3395;
wire            n3396;
wire            n3397;
wire            n3398;
wire            n3399;
wire            n34;
wire            n340;
wire            n3400;
wire            n3401;
wire            n3402;
wire            n3403;
wire            n3404;
wire            n3405;
wire            n3406;
wire            n3407;
wire            n3408;
wire            n3409;
wire            n341;
wire            n3410;
wire            n3411;
wire            n3412;
wire            n3413;
wire            n3414;
wire            n3415;
wire            n3416;
wire            n3417;
wire            n3418;
wire            n3419;
wire            n342;
wire            n3420;
wire            n3421;
wire            n3422;
wire            n3423;
wire            n3424;
wire            n3425;
wire            n3426;
wire            n3427;
wire            n3428;
wire            n3429;
wire            n343;
wire            n3430;
wire            n3431;
wire            n3432;
wire            n3433;
wire            n3434;
wire            n3435;
wire            n3436;
wire            n3437;
wire            n3438;
wire            n3439;
wire            n344;
wire            n3440;
wire            n3441;
wire            n3442;
wire            n3443;
wire            n3444;
wire            n3445;
wire            n3446;
wire            n3447;
wire            n3448;
wire            n3449;
wire            n345;
wire            n3450;
wire            n3451;
wire            n3452;
wire            n3453;
wire            n3454;
wire            n3455;
wire            n3456;
wire            n3457;
wire            n3458;
wire            n3459;
wire            n346;
wire            n3460;
wire            n3461;
wire            n3462;
wire            n3463;
wire            n3464;
wire            n3465;
wire            n3466;
wire            n3467;
wire            n3468;
wire            n3469;
wire            n347;
wire            n3470;
wire            n3471;
wire            n3472;
wire            n3473;
wire      [1:0] n3474;
wire            n3475;
wire            n3476;
wire            n3477;
wire            n3478;
wire            n3479;
wire            n348;
wire            n3480;
wire      [2:0] n3481;
wire            n3482;
wire            n3483;
wire            n3484;
wire            n3485;
wire            n3486;
wire            n3487;
wire            n3488;
wire            n3489;
wire            n349;
wire            n3490;
wire            n3491;
wire            n3492;
wire            n3493;
wire            n3494;
wire            n3495;
wire            n3496;
wire            n3497;
wire            n3498;
wire            n3499;
wire            n35;
wire            n350;
wire            n3500;
wire            n3501;
wire            n3502;
wire            n3503;
wire            n3504;
wire            n3505;
wire            n3506;
wire            n3507;
wire            n3508;
wire            n3509;
wire            n351;
wire            n3510;
wire            n3511;
wire            n3512;
wire            n3513;
wire            n3514;
wire            n3515;
wire            n3516;
wire            n3517;
wire            n3518;
wire            n3519;
wire            n352;
wire            n3520;
wire            n3521;
wire            n3522;
wire            n3523;
wire            n3524;
wire            n3525;
wire            n3526;
wire            n3527;
wire            n3528;
wire            n3529;
wire            n353;
wire            n3530;
wire            n3531;
wire            n3532;
wire            n3533;
wire            n3534;
wire            n3535;
wire            n3536;
wire            n3537;
wire            n3538;
wire            n3539;
wire            n354;
wire            n3540;
wire            n3541;
wire            n3542;
wire            n3543;
wire            n3544;
wire            n3545;
wire            n3546;
wire            n3547;
wire            n3548;
wire            n3549;
wire            n355;
wire            n3550;
wire            n3551;
wire            n3552;
wire            n3553;
wire            n3554;
wire            n3555;
wire            n3556;
wire            n3557;
wire            n3558;
wire            n3559;
wire            n356;
wire            n3560;
wire            n3561;
wire            n3562;
wire            n3563;
wire            n3564;
wire            n3565;
wire            n3566;
wire            n3567;
wire            n3568;
wire            n3569;
wire            n357;
wire            n3570;
wire            n3571;
wire            n3572;
wire            n3573;
wire            n3574;
wire            n3575;
wire            n3576;
wire            n3577;
wire            n3578;
wire            n3579;
wire            n358;
wire            n3580;
wire            n3581;
wire            n3582;
wire            n3583;
wire            n3584;
wire            n3585;
wire            n3586;
wire            n3587;
wire            n3588;
wire            n3589;
wire            n359;
wire            n3590;
wire            n3591;
wire            n3592;
wire            n3593;
wire            n3594;
wire            n3595;
wire            n3596;
wire            n3597;
wire            n3598;
wire            n3599;
wire            n36;
wire            n360;
wire            n3600;
wire            n3601;
wire            n3602;
wire            n3603;
wire            n3604;
wire            n3605;
wire            n3606;
wire            n3607;
wire            n3608;
wire      [3:0] n3609;
wire            n361;
wire            n3610;
wire            n3611;
wire            n3612;
wire            n3613;
wire            n3614;
wire            n3615;
wire      [4:0] n3616;
wire            n3617;
wire            n3618;
wire            n3619;
wire            n362;
wire            n3620;
wire            n3621;
wire            n3622;
wire            n3623;
wire            n3624;
wire            n3625;
wire            n3626;
wire            n3627;
wire            n3628;
wire            n3629;
wire            n363;
wire            n3630;
wire            n3631;
wire            n3632;
wire            n3633;
wire            n3634;
wire            n3635;
wire            n3636;
wire            n3637;
wire            n3638;
wire            n3639;
wire            n364;
wire            n3640;
wire            n3641;
wire            n3642;
wire            n3643;
wire            n3644;
wire            n3645;
wire            n3646;
wire            n3647;
wire            n3648;
wire            n3649;
wire            n365;
wire            n3650;
wire            n3651;
wire            n3652;
wire            n3653;
wire            n3654;
wire            n3655;
wire            n3656;
wire            n3657;
wire            n3658;
wire            n3659;
wire            n366;
wire            n3660;
wire            n3661;
wire            n3662;
wire            n3663;
wire            n3664;
wire            n3665;
wire            n3666;
wire            n3667;
wire            n3668;
wire            n3669;
wire            n367;
wire            n3670;
wire            n3671;
wire            n3672;
wire            n3673;
wire            n3674;
wire            n3675;
wire            n3676;
wire            n3677;
wire            n3678;
wire            n3679;
wire            n368;
wire            n3680;
wire            n3681;
wire            n3682;
wire            n3683;
wire            n3684;
wire            n3685;
wire            n3686;
wire            n3687;
wire            n3688;
wire            n3689;
wire            n369;
wire            n3690;
wire            n3691;
wire            n3692;
wire            n3693;
wire            n3694;
wire            n3695;
wire            n3696;
wire            n3697;
wire            n3698;
wire            n3699;
wire            n37;
wire            n370;
wire            n3700;
wire            n3701;
wire            n3702;
wire            n3703;
wire            n3704;
wire            n3705;
wire            n3706;
wire            n3707;
wire            n3708;
wire            n3709;
wire            n371;
wire            n3710;
wire            n3711;
wire            n3712;
wire            n3713;
wire            n3714;
wire            n3715;
wire            n3716;
wire            n3717;
wire            n3718;
wire            n3719;
wire            n372;
wire            n3720;
wire            n3721;
wire            n3722;
wire            n3723;
wire            n3724;
wire            n3725;
wire            n3726;
wire            n3727;
wire            n3728;
wire            n3729;
wire            n373;
wire            n3730;
wire            n3731;
wire            n3732;
wire            n3733;
wire            n3734;
wire            n3735;
wire            n3736;
wire            n3737;
wire            n3738;
wire            n3739;
wire            n374;
wire            n3740;
wire            n3741;
wire            n3742;
wire            n3743;
wire            n3744;
wire            n3745;
wire            n3746;
wire            n3747;
wire            n3748;
wire            n3749;
wire            n375;
wire            n3750;
wire            n3751;
wire            n3752;
wire            n3753;
wire            n3754;
wire            n3755;
wire            n3756;
wire            n3757;
wire            n3758;
wire            n3759;
wire            n376;
wire            n3760;
wire            n3761;
wire      [5:0] n3762;
wire            n3763;
wire            n3764;
wire            n3765;
wire            n3766;
wire            n3767;
wire            n3768;
wire      [6:0] n3769;
wire            n377;
wire            n3770;
wire            n3771;
wire            n3772;
wire            n3773;
wire            n3774;
wire            n3775;
wire            n3776;
wire            n3777;
wire            n3778;
wire            n3779;
wire            n378;
wire            n3780;
wire            n3781;
wire            n3782;
wire            n3783;
wire            n3784;
wire            n3785;
wire            n3786;
wire            n3787;
wire            n3788;
wire            n3789;
wire            n379;
wire            n3790;
wire            n3791;
wire            n3792;
wire            n3793;
wire            n3794;
wire            n3795;
wire            n3796;
wire            n3797;
wire            n3798;
wire            n3799;
wire            n38;
wire            n380;
wire            n3800;
wire            n3801;
wire            n3802;
wire            n3803;
wire            n3804;
wire            n3805;
wire            n3806;
wire            n3807;
wire            n3808;
wire            n3809;
wire            n381;
wire            n3810;
wire            n3811;
wire            n3812;
wire            n3813;
wire            n3814;
wire            n3815;
wire            n3816;
wire            n3817;
wire            n3818;
wire            n3819;
wire            n382;
wire            n3820;
wire            n3821;
wire            n3822;
wire            n3823;
wire            n3824;
wire            n3825;
wire            n3826;
wire            n3827;
wire            n3828;
wire            n3829;
wire            n383;
wire            n3830;
wire            n3831;
wire            n3832;
wire            n3833;
wire            n3834;
wire            n3835;
wire            n3836;
wire            n3837;
wire            n3838;
wire            n3839;
wire            n384;
wire            n3840;
wire            n3841;
wire            n3842;
wire            n3843;
wire            n3844;
wire            n3845;
wire            n3846;
wire            n3847;
wire            n3848;
wire      [7:0] n3849;
wire            n385;
wire            n3850;
wire            n3851;
wire            n3852;
wire            n3853;
wire            n3854;
wire            n3855;
wire      [8:0] n3856;
wire            n3857;
wire            n3858;
wire            n3859;
wire            n386;
wire            n3860;
wire            n3861;
wire            n3862;
wire            n3863;
wire            n3864;
wire            n3865;
wire            n3866;
wire            n3867;
wire            n3868;
wire            n3869;
wire            n387;
wire            n3870;
wire            n3871;
wire            n3872;
wire            n3873;
wire            n3874;
wire            n3875;
wire            n3876;
wire            n3877;
wire            n3878;
wire            n3879;
wire            n388;
wire            n3880;
wire            n3881;
wire            n3882;
wire            n3883;
wire            n3884;
wire            n3885;
wire            n3886;
wire            n3887;
wire            n3888;
wire            n3889;
wire            n389;
wire            n3890;
wire            n3891;
wire            n3892;
wire            n3893;
wire            n3894;
wire            n3895;
wire            n3896;
wire            n3897;
wire            n3898;
wire            n3899;
wire            n39;
wire            n390;
wire            n3900;
wire            n3901;
wire            n3902;
wire            n3903;
wire            n3904;
wire            n3905;
wire            n3906;
wire            n3907;
wire            n3908;
wire            n3909;
wire            n391;
wire            n3910;
wire            n3911;
wire            n3912;
wire            n3913;
wire            n3914;
wire            n3915;
wire            n3916;
wire            n3917;
wire            n3918;
wire            n3919;
wire            n392;
wire            n3920;
wire            n3921;
wire            n3922;
wire            n3923;
wire            n3924;
wire            n3925;
wire            n3926;
wire            n3927;
wire            n3928;
wire            n3929;
wire            n393;
wire            n3930;
wire            n3931;
wire            n3932;
wire            n3933;
wire            n3934;
wire            n3935;
wire            n3936;
wire            n3937;
wire            n3938;
wire            n3939;
wire            n394;
wire            n3940;
wire            n3941;
wire            n3942;
wire            n3943;
wire      [9:0] n3944;
wire            n3945;
wire            n3946;
wire            n3947;
wire            n3948;
wire            n3949;
wire            n395;
wire            n3950;
wire     [10:0] n3951;
wire            n3952;
wire            n3953;
wire            n3954;
wire            n3955;
wire            n3956;
wire            n3957;
wire            n3958;
wire            n3959;
wire            n396;
wire            n3960;
wire            n3961;
wire            n3962;
wire            n3963;
wire            n3964;
wire            n3965;
wire            n3966;
wire            n3967;
wire            n3968;
wire            n3969;
wire            n397;
wire            n3970;
wire            n3971;
wire            n3972;
wire            n3973;
wire            n3974;
wire            n3975;
wire            n3976;
wire            n3977;
wire            n3978;
wire            n3979;
wire            n398;
wire            n3980;
wire            n3981;
wire            n3982;
wire            n3983;
wire            n3984;
wire            n3985;
wire            n3986;
wire            n3987;
wire            n3988;
wire            n3989;
wire            n399;
wire            n3990;
wire            n3991;
wire            n3992;
wire            n3993;
wire            n3994;
wire            n3995;
wire            n3996;
wire            n3997;
wire            n3998;
wire            n3999;
wire            n4;
wire            n40;
wire            n400;
wire            n4000;
wire            n4001;
wire            n4002;
wire            n4003;
wire            n4004;
wire            n4005;
wire            n4006;
wire            n4007;
wire            n4008;
wire            n4009;
wire            n401;
wire            n4010;
wire            n4011;
wire            n4012;
wire            n4013;
wire            n4014;
wire            n4015;
wire            n4016;
wire            n4017;
wire            n4018;
wire            n4019;
wire            n402;
wire            n4020;
wire            n4021;
wire            n4022;
wire            n4023;
wire            n4024;
wire            n4025;
wire            n4026;
wire            n4027;
wire            n4028;
wire            n4029;
wire            n403;
wire            n4030;
wire            n4031;
wire            n4032;
wire     [11:0] n4033;
wire            n4034;
wire            n4035;
wire            n4036;
wire            n4037;
wire            n4038;
wire            n4039;
wire            n404;
wire            n4040;
wire            n4041;
wire            n4042;
wire            n4043;
wire            n4044;
wire            n4045;
wire            n4046;
wire            n4047;
wire            n4048;
wire            n4049;
wire            n405;
wire            n4050;
wire     [12:0] n4051;
wire            n4052;
wire            n4053;
wire            n4054;
wire            n4055;
wire            n4056;
wire            n4057;
wire            n4058;
wire            n4059;
wire            n406;
wire            n4060;
wire            n4061;
wire            n4062;
wire            n4063;
wire            n4064;
wire            n4065;
wire            n4066;
wire            n4067;
wire            n4068;
wire            n4069;
wire            n407;
wire            n4070;
wire            n4071;
wire            n4072;
wire            n4073;
wire            n4074;
wire            n4075;
wire            n4076;
wire            n4077;
wire            n4078;
wire            n4079;
wire            n408;
wire            n4080;
wire            n4081;
wire            n4082;
wire            n4083;
wire            n4084;
wire            n4085;
wire            n4086;
wire            n4087;
wire            n4088;
wire            n4089;
wire            n409;
wire            n4090;
wire            n4091;
wire            n4092;
wire            n4093;
wire            n4094;
wire            n4095;
wire            n4096;
wire            n4097;
wire            n4098;
wire            n4099;
wire            n41;
wire            n410;
wire            n4100;
wire            n4101;
wire            n4102;
wire            n4103;
wire            n4104;
wire            n4105;
wire            n4106;
wire            n4107;
wire            n4108;
wire            n4109;
wire            n411;
wire            n4110;
wire            n4111;
wire            n4112;
wire            n4113;
wire            n4114;
wire            n4115;
wire            n4116;
wire            n4117;
wire            n4118;
wire            n4119;
wire            n412;
wire            n4120;
wire            n4121;
wire            n4122;
wire            n4123;
wire            n4124;
wire            n4125;
wire            n4126;
wire            n4127;
wire            n4128;
wire            n4129;
wire            n413;
wire            n4130;
wire            n4131;
wire            n4132;
wire            n4133;
wire            n4134;
wire            n4135;
wire            n4136;
wire            n4137;
wire            n4138;
wire            n4139;
wire            n414;
wire            n4140;
wire            n4141;
wire            n4142;
wire            n4143;
wire            n4144;
wire            n4145;
wire            n4146;
wire     [13:0] n4147;
wire            n4148;
wire            n4149;
wire            n415;
wire            n4150;
wire            n4151;
wire            n4152;
wire            n4153;
wire            n4154;
wire            n4155;
wire            n4156;
wire            n4157;
wire            n4158;
wire            n4159;
wire            n416;
wire            n4160;
wire            n4161;
wire            n4162;
wire            n4163;
wire            n4164;
wire            n4165;
wire            n4166;
wire            n4167;
wire            n4168;
wire            n4169;
wire            n417;
wire            n4170;
wire            n4171;
wire            n4172;
wire     [14:0] n4173;
wire            n4174;
wire            n4175;
wire            n4176;
wire            n4177;
wire            n4178;
wire            n4179;
wire            n418;
wire            n4180;
wire            n4181;
wire            n4182;
wire            n4183;
wire            n4184;
wire            n4185;
wire            n4186;
wire            n4187;
wire            n4188;
wire            n4189;
wire            n419;
wire            n4190;
wire            n4191;
wire            n4192;
wire            n4193;
wire            n4194;
wire            n4195;
wire            n4196;
wire            n4197;
wire            n4198;
wire            n4199;
wire            n42;
wire            n420;
wire            n4200;
wire            n4201;
wire            n4202;
wire            n4203;
wire            n4204;
wire     [15:0] n4205;
wire            n4206;
wire            n4207;
wire            n4208;
wire            n4209;
wire            n421;
wire            n4210;
wire            n4211;
wire            n4212;
wire            n4213;
wire            n4214;
wire            n4215;
wire            n4216;
wire            n4217;
wire            n4218;
wire            n4219;
wire            n422;
wire            n4220;
wire            n4221;
wire            n4222;
wire            n4223;
wire            n4224;
wire            n4225;
wire            n4226;
wire            n4227;
wire     [16:0] n4228;
wire            n4229;
wire            n423;
wire            n4230;
wire            n4231;
wire            n4232;
wire            n4233;
wire            n4234;
wire            n4235;
wire            n4236;
wire            n4237;
wire            n4238;
wire            n4239;
wire            n424;
wire            n4240;
wire            n4241;
wire            n4242;
wire            n4243;
wire            n4244;
wire            n4245;
wire            n4246;
wire            n4247;
wire            n4248;
wire            n4249;
wire            n425;
wire            n4250;
wire            n4251;
wire            n4252;
wire            n4253;
wire            n4254;
wire            n4255;
wire            n4256;
wire            n4257;
wire     [17:0] n4258;
wire            n4259;
wire            n426;
wire            n4260;
wire            n4261;
wire            n4262;
wire            n4263;
wire            n4264;
wire            n4265;
wire            n4266;
wire            n4267;
wire            n4268;
wire            n4269;
wire            n427;
wire            n4270;
wire            n4271;
wire            n4272;
wire            n4273;
wire            n4274;
wire            n4275;
wire            n4276;
wire            n4277;
wire            n4278;
wire            n4279;
wire            n428;
wire     [18:0] n4280;
wire            n4281;
wire            n4282;
wire            n4283;
wire            n4284;
wire            n4285;
wire            n4286;
wire            n4287;
wire            n4288;
wire            n4289;
wire            n429;
wire            n4290;
wire            n4291;
wire            n4292;
wire            n4293;
wire            n4294;
wire            n4295;
wire            n4296;
wire            n4297;
wire            n4298;
wire            n4299;
wire            n43;
wire            n430;
wire            n4300;
wire            n4301;
wire            n4302;
wire            n4303;
wire            n4304;
wire            n4305;
wire            n4306;
wire            n4307;
wire            n4308;
wire     [19:0] n4309;
wire            n431;
wire            n4310;
wire            n4311;
wire            n4312;
wire            n4313;
wire            n4314;
wire            n4315;
wire            n4316;
wire            n4317;
wire            n4318;
wire            n4319;
wire            n432;
wire            n4320;
wire            n4321;
wire            n4322;
wire            n4323;
wire            n4324;
wire            n4325;
wire            n4326;
wire            n4327;
wire            n4328;
wire            n4329;
wire            n433;
wire            n4330;
wire     [20:0] n4331;
wire            n4332;
wire            n4333;
wire            n4334;
wire            n4335;
wire            n4336;
wire            n4337;
wire            n4338;
wire            n4339;
wire            n434;
wire            n4340;
wire            n4341;
wire            n4342;
wire            n4343;
wire            n4344;
wire            n4345;
wire            n4346;
wire            n4347;
wire            n4348;
wire            n4349;
wire            n435;
wire            n4350;
wire            n4351;
wire            n4352;
wire            n4353;
wire            n4354;
wire            n4355;
wire            n4356;
wire            n4357;
wire            n4358;
wire            n4359;
wire            n436;
wire     [21:0] n4360;
wire            n4361;
wire            n4362;
wire            n4363;
wire            n4364;
wire            n4365;
wire            n4366;
wire            n4367;
wire            n4368;
wire            n4369;
wire            n437;
wire            n4370;
wire            n4371;
wire            n4372;
wire            n4373;
wire            n4374;
wire            n4375;
wire            n4376;
wire            n4377;
wire            n4378;
wire            n4379;
wire            n438;
wire            n4380;
wire     [22:0] n4381;
wire            n4382;
wire            n4383;
wire            n4384;
wire            n4385;
wire            n4386;
wire            n4387;
wire            n4388;
wire            n4389;
wire            n439;
wire            n4390;
wire            n4391;
wire            n4392;
wire            n4393;
wire            n4394;
wire            n4395;
wire            n4396;
wire            n4397;
wire            n4398;
wire            n4399;
wire            n44;
wire            n440;
wire            n4400;
wire            n4401;
wire            n4402;
wire            n4403;
wire            n4404;
wire            n4405;
wire            n4406;
wire            n4407;
wire     [23:0] n4408;
wire            n4409;
wire            n441;
wire            n4410;
wire            n4411;
wire            n4412;
wire            n4413;
wire            n4414;
wire            n4415;
wire            n4416;
wire            n4417;
wire            n4418;
wire            n4419;
wire            n442;
wire            n4420;
wire            n4421;
wire            n4422;
wire            n4423;
wire            n4424;
wire            n4425;
wire     [24:0] n4426;
wire            n4427;
wire            n4428;
wire            n4429;
wire            n443;
wire            n4430;
wire            n4431;
wire            n4432;
wire            n4433;
wire            n4434;
wire            n4435;
wire            n4436;
wire            n4437;
wire            n4438;
wire            n4439;
wire            n444;
wire            n4440;
wire            n4441;
wire            n4442;
wire            n4443;
wire            n4444;
wire            n4445;
wire            n4446;
wire            n4447;
wire            n4448;
wire            n4449;
wire            n445;
wire            n4450;
wire            n4451;
wire     [25:0] n4452;
wire            n4453;
wire            n4454;
wire            n4455;
wire            n4456;
wire            n4457;
wire            n4458;
wire            n4459;
wire            n446;
wire            n4460;
wire            n4461;
wire            n4462;
wire            n4463;
wire            n4464;
wire            n4465;
wire            n4466;
wire            n4467;
wire            n4468;
wire     [26:0] n4469;
wire            n447;
wire            n4470;
wire            n4471;
wire            n4472;
wire            n4473;
wire            n4474;
wire            n4475;
wire            n4476;
wire            n4477;
wire            n4478;
wire            n4479;
wire            n448;
wire            n4480;
wire            n4481;
wire            n4482;
wire            n4483;
wire            n4484;
wire            n4485;
wire            n4486;
wire            n4487;
wire            n4488;
wire            n4489;
wire            n449;
wire            n4490;
wire            n4491;
wire            n4492;
wire            n4493;
wire     [27:0] n4494;
wire            n4495;
wire            n4496;
wire            n4497;
wire            n4498;
wire            n4499;
wire            n45;
wire            n450;
wire            n4500;
wire            n4501;
wire            n4502;
wire            n4503;
wire            n4504;
wire            n4505;
wire            n4506;
wire            n4507;
wire     [28:0] n4508;
wire            n4509;
wire            n451;
wire            n4510;
wire            n4511;
wire            n4512;
wire            n4513;
wire            n4514;
wire            n4515;
wire            n4516;
wire            n4517;
wire            n4518;
wire            n4519;
wire            n452;
wire            n4520;
wire            n4521;
wire            n4522;
wire            n4523;
wire            n4524;
wire            n4525;
wire            n4526;
wire            n4527;
wire            n4528;
wire            n4529;
wire            n453;
wire            n4530;
wire            n4531;
wire            n4532;
wire            n4533;
wire     [29:0] n4534;
wire            n4535;
wire            n4536;
wire            n4537;
wire            n4538;
wire            n4539;
wire            n454;
wire            n4540;
wire            n4541;
wire            n4542;
wire            n4543;
wire            n4544;
wire            n4545;
wire            n4546;
wire     [30:0] n4547;
wire            n4548;
wire            n4549;
wire            n455;
wire            n4550;
wire            n4551;
wire            n4552;
wire     [31:0] n4553;
wire            n456;
wire            n457;
wire            n458;
wire            n459;
wire            n46;
wire            n460;
wire            n461;
wire            n462;
wire            n463;
wire            n464;
wire            n465;
wire            n466;
wire            n467;
wire            n468;
wire            n469;
wire            n47;
wire            n470;
wire            n471;
wire            n472;
wire            n473;
wire            n474;
wire            n475;
wire            n476;
wire            n477;
wire            n478;
wire            n479;
wire            n48;
wire            n480;
wire            n481;
wire            n482;
wire            n483;
wire            n484;
wire            n485;
wire            n486;
wire            n487;
wire            n488;
wire            n489;
wire            n49;
wire            n490;
wire            n491;
wire            n492;
wire            n493;
wire            n494;
wire            n495;
wire            n496;
wire            n497;
wire            n498;
wire            n499;
wire            n5;
wire            n50;
wire            n500;
wire            n501;
wire            n502;
wire            n503;
wire            n504;
wire            n505;
wire            n506;
wire            n507;
wire            n508;
wire            n509;
wire            n51;
wire            n510;
wire            n511;
wire            n512;
wire            n513;
wire            n514;
wire            n515;
wire            n516;
wire            n517;
wire            n518;
wire            n519;
wire            n52;
wire            n520;
wire            n521;
wire            n522;
wire            n523;
wire            n524;
wire            n525;
wire            n526;
wire            n527;
wire            n528;
wire            n529;
wire            n53;
wire            n530;
wire            n531;
wire            n532;
wire            n533;
wire            n534;
wire            n535;
wire            n536;
wire            n537;
wire            n538;
wire            n539;
wire            n54;
wire            n540;
wire            n541;
wire            n542;
wire            n543;
wire            n544;
wire            n545;
wire            n546;
wire            n547;
wire            n548;
wire            n549;
wire            n55;
wire            n550;
wire            n551;
wire            n552;
wire            n553;
wire            n554;
wire            n555;
wire            n556;
wire            n557;
wire            n558;
wire            n559;
wire            n56;
wire            n560;
wire            n561;
wire            n562;
wire            n563;
wire            n564;
wire            n565;
wire            n566;
wire            n567;
wire            n568;
wire            n569;
wire            n57;
wire            n570;
wire            n571;
wire            n572;
wire            n573;
wire            n574;
wire            n575;
wire            n576;
wire            n577;
wire            n578;
wire            n579;
wire            n58;
wire            n580;
wire            n581;
wire            n582;
wire            n583;
wire            n584;
wire            n585;
wire            n586;
wire            n587;
wire            n588;
wire            n589;
wire            n59;
wire            n590;
wire            n591;
wire            n592;
wire            n593;
wire            n594;
wire            n595;
wire            n596;
wire            n597;
wire            n598;
wire            n599;
wire            n6;
wire            n60;
wire            n600;
wire            n601;
wire            n602;
wire            n603;
wire            n604;
wire            n605;
wire            n606;
wire            n607;
wire            n608;
wire            n609;
wire            n61;
wire            n610;
wire            n611;
wire            n612;
wire            n613;
wire            n614;
wire            n615;
wire            n616;
wire            n617;
wire            n618;
wire            n619;
wire            n62;
wire            n620;
wire            n621;
wire            n622;
wire            n623;
wire            n624;
wire            n625;
wire            n626;
wire            n627;
wire            n628;
wire            n629;
wire            n63;
wire            n630;
wire            n631;
wire            n632;
wire            n633;
wire            n634;
wire            n635;
wire            n636;
wire            n637;
wire            n638;
wire            n639;
wire            n64;
wire            n640;
wire            n641;
wire            n642;
wire            n643;
wire            n644;
wire            n645;
wire            n646;
wire            n647;
wire            n648;
wire            n649;
wire            n65;
wire            n650;
wire            n651;
wire            n652;
wire            n653;
wire            n654;
wire            n655;
wire            n656;
wire            n657;
wire            n658;
wire            n659;
wire            n66;
wire            n660;
wire            n661;
wire            n662;
wire            n663;
wire            n664;
wire            n665;
wire            n666;
wire            n667;
wire            n668;
wire            n669;
wire            n67;
wire            n670;
wire            n671;
wire            n672;
wire            n673;
wire            n674;
wire            n675;
wire            n676;
wire            n677;
wire            n678;
wire            n679;
wire            n68;
wire            n680;
wire            n681;
wire            n682;
wire            n683;
wire            n684;
wire            n685;
wire            n686;
wire            n687;
wire            n688;
wire            n689;
wire            n69;
wire            n690;
wire            n691;
wire            n692;
wire            n693;
wire            n694;
wire            n695;
wire            n696;
wire            n697;
wire            n698;
wire            n699;
wire            n7;
wire            n70;
wire            n700;
wire            n701;
wire            n702;
wire            n703;
wire            n704;
wire            n705;
wire            n706;
wire            n707;
wire            n708;
wire            n709;
wire            n71;
wire            n710;
wire            n711;
wire            n712;
wire            n713;
wire            n714;
wire            n715;
wire            n716;
wire            n717;
wire            n718;
wire            n719;
wire            n72;
wire            n720;
wire            n721;
wire            n722;
wire            n723;
wire            n724;
wire            n725;
wire            n726;
wire            n727;
wire            n728;
wire            n729;
wire            n73;
wire            n730;
wire            n731;
wire            n732;
wire            n733;
wire            n734;
wire            n735;
wire            n736;
wire            n737;
wire            n738;
wire            n739;
wire            n740;
wire            n741;
wire            n742;
wire            n743;
wire            n744;
wire            n745;
wire            n746;
wire            n747;
wire            n748;
wire            n749;
wire            n75;
wire            n750;
wire            n751;
wire            n752;
wire            n753;
wire            n754;
wire            n755;
wire            n756;
wire            n757;
wire            n758;
wire            n759;
wire            n76;
wire            n760;
wire            n761;
wire            n762;
wire            n763;
wire            n764;
wire            n765;
wire            n766;
wire            n767;
wire            n768;
wire            n769;
wire            n77;
wire            n770;
wire            n771;
wire            n772;
wire            n773;
wire            n774;
wire            n775;
wire            n776;
wire            n777;
wire            n778;
wire            n779;
wire            n78;
wire            n780;
wire            n781;
wire            n782;
wire            n783;
wire            n784;
wire            n785;
wire            n786;
wire            n787;
wire            n788;
wire            n789;
wire            n79;
wire            n790;
wire            n791;
wire            n792;
wire            n793;
wire            n794;
wire            n795;
wire            n796;
wire            n797;
wire            n798;
wire            n799;
wire            n8;
wire            n80;
wire            n800;
wire            n801;
wire            n802;
wire            n803;
wire            n804;
wire            n805;
wire            n806;
wire            n807;
wire            n808;
wire            n809;
wire            n81;
wire            n810;
wire            n811;
wire            n812;
wire            n813;
wire            n814;
wire            n815;
wire            n816;
wire            n817;
wire            n818;
wire            n819;
wire            n82;
wire            n820;
wire            n821;
wire            n822;
wire            n823;
wire            n824;
wire            n825;
wire            n826;
wire            n827;
wire            n828;
wire            n829;
wire            n83;
wire            n830;
wire            n831;
wire            n832;
wire            n833;
wire            n834;
wire            n835;
wire            n836;
wire            n837;
wire            n838;
wire            n839;
wire            n84;
wire            n840;
wire            n841;
wire            n842;
wire            n843;
wire            n844;
wire            n845;
wire            n846;
wire            n847;
wire            n848;
wire            n849;
wire            n85;
wire            n850;
wire            n851;
wire            n852;
wire            n853;
wire            n854;
wire            n855;
wire            n856;
wire            n857;
wire            n858;
wire            n859;
wire            n86;
wire            n860;
wire            n861;
wire            n862;
wire            n863;
wire            n864;
wire            n865;
wire            n866;
wire            n867;
wire            n868;
wire            n869;
wire            n87;
wire            n870;
wire            n871;
wire            n872;
wire            n873;
wire            n874;
wire            n875;
wire            n876;
wire            n877;
wire            n878;
wire            n879;
wire            n88;
wire            n880;
wire            n881;
wire            n882;
wire            n883;
wire            n884;
wire            n885;
wire            n886;
wire            n887;
wire            n888;
wire            n889;
wire            n89;
wire            n890;
wire            n891;
wire            n892;
wire            n893;
wire            n894;
wire            n895;
wire            n896;
wire            n897;
wire            n898;
wire            n899;
wire            n9;
wire            n90;
wire            n900;
wire            n901;
wire            n902;
wire            n903;
wire            n904;
wire            n905;
wire            n906;
wire            n907;
wire            n908;
wire            n909;
wire            n91;
wire            n910;
wire            n911;
wire            n912;
wire            n913;
wire            n914;
wire            n915;
wire            n916;
wire            n917;
wire            n918;
wire            n919;
wire            n92;
wire            n920;
wire            n921;
wire            n922;
wire            n923;
wire            n924;
wire            n925;
wire            n926;
wire            n927;
wire            n928;
wire            n929;
wire            n93;
wire            n930;
wire            n931;
wire            n932;
wire            n933;
wire            n934;
wire            n935;
wire            n936;
wire            n937;
wire            n938;
wire            n939;
wire            n94;
wire            n940;
wire            n941;
wire            n942;
wire            n943;
wire            n944;
wire            n945;
wire            n946;
wire            n947;
wire            n948;
wire            n949;
wire            n95;
wire            n950;
wire            n951;
wire            n952;
wire            n953;
wire            n954;
wire            n955;
wire            n956;
wire            n957;
wire            n958;
wire            n959;
wire            n96;
wire            n960;
wire            n961;
wire            n962;
wire            n963;
wire            n964;
wire            n965;
wire            n966;
wire            n967;
wire            n968;
wire            n969;
wire            n97;
wire            n970;
wire            n971;
wire            n972;
wire            n973;
wire            n974;
wire            n975;
wire            n976;
wire            n977;
wire            n978;
wire            n979;
wire            n98;
wire            n980;
wire            n981;
wire            n982;
wire            n983;
wire            n984;
wire            n985;
wire            n986;
wire            n987;
wire            n988;
wire            n989;
wire            n99;
wire            n990;
wire            n991;
wire            n992;
wire            n993;
wire            n994;
wire            n995;
wire            n996;
wire            n997;
wire            n998;
wire            n999;
wire            rst;
assign __ILA_bar_valid__ = 1'b1 ;
assign __ILA_bar_decode_of_i1__ = 1'b1 ;
assign n1 = ki[1:1] ;
assign bv_1_1_n2 = 1'h1 ;
assign n3 =  ( n1 ) == ( bv_1_1_n2 )  ;
assign n4 = ki[0:0] ;
assign n5 =  ( n4 ) == ( bv_1_1_n2 )  ;
assign n6 =  ( n3 ) | ( n5 )  ;
assign n7 = ki[1:1] ;
assign n8 =  ( n7 ) == ( bv_1_1_n2 )  ;
assign n9 = i_wb_data[1:1] ;
assign n10 = ~ ( n9 ) ;
assign n11 = sp[1:1] ;
assign n12 =  ( n10 ) ^ ( n11 )  ;
assign n13 = i_wb_data[1:1] ;
assign n14 = sp[1:1] ;
assign n15 = ~ ( n14 ) ;
assign n16 =  ( n13 ) | ( n15 )  ;
assign n17 = ~ ( n16 ) ;
assign n18 = i_wb_data[1:1] ;
assign n19 = ~ ( n18 ) ;
assign n20 = sp[1:1] ;
assign n21 =  ( n19 ) ^ ( n20 )  ;
assign n22 = ~ ( n21 ) ;
assign n23 = i_wb_data[1:1] ;
assign n24 =  ( n22 ) | ( n23 )  ;
assign n25 = sp[1:1] ;
assign n26 = ~ ( n25 ) ;
assign n27 =  ( n24 ) | ( n26 )  ;
assign n28 = ~ ( n27 ) ;
assign n29 =  ( n17 ) | ( n28 )  ;
assign n30 =  ( n17 ) | ( n28 )  ;
assign n31 = ~ ( n30 ) ;
assign n32 =  ( n22 ) | ( n31 )  ;
assign n33 = ~ ( n32 ) ;
assign n34 =  ( n29 ) | ( n33 )  ;
assign n35 =  ( n17 ) | ( n28 )  ;
assign n36 =  ( n35 ) | ( n33 )  ;
assign n37 = ~ ( n36 ) ;
assign n38 =  ( n22 ) | ( n37 )  ;
assign n39 = ~ ( n38 ) ;
assign n40 =  ( n34 ) | ( n39 )  ;
assign n41 =  ( n17 ) | ( n28 )  ;
assign n42 =  ( n41 ) | ( n33 )  ;
assign n43 =  ( n17 ) | ( n28 )  ;
assign n44 = i_wb_data[0:0] ;
assign n45 = sp[0:0] ;
assign n46 = ~ ( n45 ) ;
assign n47 =  ( n44 ) | ( n46 )  ;
assign n48 = ~ ( n47 ) ;
assign n49 = i_wb_data[0:0] ;
assign n50 = ~ ( n49 ) ;
assign n51 = sp[0:0] ;
assign n52 =  ( n50 ) ^ ( n51 )  ;
assign n53 =  ( n48 ) | ( n52 )  ;
assign n54 = ~ ( n53 ) ;
assign n55 =  ( n22 ) | ( n54 )  ;
assign n56 = ~ ( n55 ) ;
assign n57 =  ( n43 ) | ( n56 )  ;
assign n58 = ~ ( n57 ) ;
assign n59 =  ( n22 ) | ( n58 )  ;
assign n60 = ~ ( n59 ) ;
assign n61 =  ( n42 ) | ( n60 )  ;
assign n62 = ~ ( n61 ) ;
assign n63 =  ( n22 ) | ( n62 )  ;
assign n64 = ~ ( n63 ) ;
assign n65 =  ( n40 ) | ( n64 )  ;
assign n66 =  ( n12 ) ^ ( n65 )  ;
assign n67 = ~ ( n66 ) ;
assign n68 = i_wb_data[1:1] ;
assign n69 = ~ ( n68 ) ;
assign n70 = sp[1:1] ;
assign n71 =  ( n69 ) ^ ( n70 )  ;
assign n72 =  ( n71 ) ^ ( n65 )  ;
assign n73 =  ( n8 ) ? ( n67 ) : ( n72 ) ;
assign bv_1_0_n74 = 1'h0 ;
assign n75 =  ( n6 ) ? ( n73 ) : ( bv_1_0_n74 ) ;
assign n76 = ki[1:1] ;
assign n77 =  ( n76 ) == ( bv_1_0_n74 )  ;
assign n78 = i_wb_data[1:1] ;
assign n79 = ~ ( n78 ) ;
assign n80 = sp[1:1] ;
assign n81 =  ( n79 ) ^ ( n80 )  ;
assign n82 =  ( n17 ) | ( n28 )  ;
assign n83 =  ( n82 ) | ( n33 )  ;
assign n84 =  ( n83 ) | ( n39 )  ;
assign n85 =  ( n17 ) | ( n28 )  ;
assign n86 =  ( n85 ) | ( n33 )  ;
assign n87 = ~ ( n53 ) ;
assign n88 =  ( n22 ) | ( n87 )  ;
assign n89 = ~ ( n88 ) ;
assign n90 =  ( n86 ) | ( n89 )  ;
assign n91 = ~ ( n90 ) ;
assign n92 =  ( n22 ) | ( n91 )  ;
assign n93 = ~ ( n92 ) ;
assign n94 =  ( n84 ) | ( n93 )  ;
assign n95 = ~ ( n94 ) ;
assign n96 =  ( n22 ) | ( n95 )  ;
assign n97 = ~ ( n96 ) ;
assign n98 =  ( n17 ) | ( n97 )  ;
assign n99 =  ( n81 ) ^ ( n98 )  ;
assign n100 =  ( n77 ) ? ( bv_1_0_n74 ) : ( n99 ) ;
assign n101 = ~ ( n100 ) ;
assign n102 =  ( n75 ) | ( n101 )  ;
assign n103 = ki[1:1] ;
assign n104 =  ( n103 ) == ( bv_1_0_n74 )  ;
assign n105 = i_wb_data[1:1] ;
assign n106 = ~ ( n105 ) ;
assign n107 = sp[1:1] ;
assign n108 =  ( n106 ) ^ ( n107 )  ;
assign n109 =  ( n108 ) ^ ( n65 )  ;
assign n110 =  ( n104 ) ? ( bv_1_0_n74 ) : ( n109 ) ;
assign n111 = ~ ( n110 ) ;
assign n112 =  ( n102 ) | ( n111 )  ;
assign n113 = ~ ( n112 ) ;
assign n114 = ~ ( n100 ) ;
assign n115 =  ( n75 ) | ( n114 )  ;
assign n116 = ~ ( n115 ) ;
assign n117 =  ( n116 ) ^ ( n110 )  ;
assign n118 =  ( n113 ) | ( n117 )  ;
assign n119 = ~ ( n118 ) ;
assign n120 =  ( n119 ) | ( n110 )  ;
assign n121 = ~ ( n120 ) ;
assign n122 = ~ ( n118 ) ;
assign n123 =  ( n122 ) | ( n110 )  ;
assign n124 = ~ ( n123 ) ;
assign n125 = ki[0:0] ;
assign n126 =  ( n125 ) == ( bv_1_1_n2 )  ;
assign n127 = ki[1:1] ;
assign n128 =  ( n127 ) == ( bv_1_0_n74 )  ;
assign n129 =  ( n126 ) | ( n128 )  ;
assign n130 = ki[1:1] ;
assign n131 =  ( n130 ) == ( bv_1_1_n2 )  ;
assign n132 = ki[0:0] ;
assign n133 =  ( n132 ) == ( bv_1_1_n2 )  ;
assign n134 =  ( n131 ) | ( n133 )  ;
assign n135 = ki[1:1] ;
assign n136 =  ( n135 ) == ( bv_1_1_n2 )  ;
assign n137 = i_wb_data[1:1] ;
assign n138 = ~ ( n137 ) ;
assign n139 = sp[1:1] ;
assign n140 =  ( n138 ) ^ ( n139 )  ;
assign n141 =  ( n140 ) ^ ( n98 )  ;
assign n142 = ~ ( n141 ) ;
assign n143 = i_wb_data[1:1] ;
assign n144 = ~ ( n143 ) ;
assign n145 = sp[1:1] ;
assign n146 =  ( n144 ) ^ ( n145 )  ;
assign n147 =  ( n146 ) ^ ( n98 )  ;
assign n148 =  ( n136 ) ? ( n142 ) : ( n147 ) ;
assign n149 =  ( n134 ) ? ( n148 ) : ( bv_1_0_n74 ) ;
assign n150 =  ( n129 ) ? ( n75 ) : ( n149 ) ;
assign n151 = ~ ( n150 ) ;
assign n152 =  ( n124 ) | ( n151 )  ;
assign n153 = ki[1:1] ;
assign n154 =  ( n153 ) == ( bv_1_0_n74 )  ;
assign n155 = i_wb_data[1:1] ;
assign n156 = ~ ( n155 ) ;
assign n157 = sp[1:1] ;
assign n158 =  ( n156 ) ^ ( n157 )  ;
assign n159 =  ( n158 ) ^ ( n94 )  ;
assign n160 =  ( n154 ) ? ( bv_1_0_n74 ) : ( n159 ) ;
assign n161 = ~ ( n160 ) ;
assign n162 =  ( n152 ) | ( n161 )  ;
assign n163 = ~ ( n75 ) ;
assign n164 =  ( n163 ) ^ ( n100 )  ;
assign n165 = ~ ( n164 ) ;
assign n166 =  ( n162 ) | ( n165 )  ;
assign n167 = ~ ( n100 ) ;
assign n168 =  ( n75 ) | ( n167 )  ;
assign n169 = ~ ( n168 ) ;
assign n170 =  ( bv_1_1_n2 ) ^ ( n169 )  ;
assign n171 =  ( n170 ) ^ ( n110 )  ;
assign n172 = ~ ( n171 ) ;
assign n173 =  ( n166 ) | ( n172 )  ;
assign n174 = ~ ( n110 ) ;
assign n175 =  ( n118 ) ^ ( n174 )  ;
assign n176 = ~ ( n175 ) ;
assign n177 =  ( n173 ) | ( n176 )  ;
assign n178 = ~ ( n177 ) ;
assign n179 =  ( n121 ) | ( n178 )  ;
assign n180 = ~ ( n118 ) ;
assign n181 =  ( n180 ) | ( n110 )  ;
assign n182 = ~ ( n181 ) ;
assign n183 = ~ ( n150 ) ;
assign n184 = ~ ( n160 ) ;
assign n185 =  ( n183 ) | ( n184 )  ;
assign n186 = ~ ( n75 ) ;
assign n187 =  ( n186 ) ^ ( n100 )  ;
assign n188 = ~ ( n187 ) ;
assign n189 =  ( n185 ) | ( n188 )  ;
assign n190 = ~ ( n171 ) ;
assign n191 =  ( n189 ) | ( n190 )  ;
assign n192 = ~ ( n110 ) ;
assign n193 =  ( n118 ) ^ ( n192 )  ;
assign n194 = ~ ( n193 ) ;
assign n195 =  ( n191 ) | ( n194 )  ;
assign n196 = ~ ( n195 ) ;
assign n197 = ~ ( n118 ) ;
assign n198 =  ( n197 ) | ( n110 )  ;
assign n199 =  ( n196 ) ^ ( n198 )  ;
assign n200 = ~ ( n199 ) ;
assign n201 =  ( n182 ) | ( n200 )  ;
assign n202 = ki[0:0] ;
assign n203 =  ( n202 ) == ( bv_1_1_n2 )  ;
assign n204 = ki[1:1] ;
assign n205 =  ( n204 ) == ( bv_1_0_n74 )  ;
assign n206 =  ( n203 ) | ( n205 )  ;
assign n207 = ki[1:1] ;
assign n208 =  ( n207 ) == ( bv_1_1_n2 )  ;
assign n209 = ki[0:0] ;
assign n210 =  ( n209 ) == ( bv_1_1_n2 )  ;
assign n211 =  ( n208 ) | ( n210 )  ;
assign n212 = ki[1:1] ;
assign n213 =  ( n212 ) == ( bv_1_1_n2 )  ;
assign n214 = i_wb_data[1:1] ;
assign n215 = ~ ( n214 ) ;
assign n216 = sp[1:1] ;
assign n217 =  ( n215 ) ^ ( n216 )  ;
assign n218 =  ( n217 ) ^ ( n94 )  ;
assign n219 = ~ ( n218 ) ;
assign n220 = i_wb_data[1:1] ;
assign n221 = ~ ( n220 ) ;
assign n222 = sp[1:1] ;
assign n223 =  ( n221 ) ^ ( n222 )  ;
assign n224 =  ( n223 ) ^ ( n94 )  ;
assign n225 =  ( n213 ) ? ( n219 ) : ( n224 ) ;
assign n226 =  ( n211 ) ? ( n225 ) : ( bv_1_0_n74 ) ;
assign n227 =  ( n206 ) ? ( n149 ) : ( n226 ) ;
assign n228 = ~ ( n227 ) ;
assign n229 = ki[1:1] ;
assign n230 =  ( n229 ) == ( bv_1_0_n74 )  ;
assign n231 = i_wb_data[1:1] ;
assign n232 = ~ ( n231 ) ;
assign n233 = sp[1:1] ;
assign n234 =  ( n232 ) ^ ( n233 )  ;
assign n235 =  ( n17 ) | ( n28 )  ;
assign n236 =  ( n235 ) | ( n33 )  ;
assign n237 =  ( n236 ) | ( n39 )  ;
assign n238 = ~ ( n57 ) ;
assign n239 =  ( n22 ) | ( n238 )  ;
assign n240 = ~ ( n239 ) ;
assign n241 =  ( n237 ) | ( n240 )  ;
assign n242 = ~ ( n241 ) ;
assign n243 =  ( n22 ) | ( n242 )  ;
assign n244 = ~ ( n243 ) ;
assign n245 =  ( n17 ) | ( n244 )  ;
assign n246 =  ( n234 ) ^ ( n245 )  ;
assign n247 =  ( n230 ) ? ( bv_1_0_n74 ) : ( n246 ) ;
assign n248 = ~ ( n247 ) ;
assign n249 =  ( n228 ) | ( n248 )  ;
assign n250 =  ( n150 ) ^ ( n160 )  ;
assign n251 = ~ ( n250 ) ;
assign n252 =  ( n249 ) | ( n251 )  ;
assign n253 = ~ ( n150 ) ;
assign n254 = ~ ( n160 ) ;
assign n255 =  ( n253 ) | ( n254 )  ;
assign n256 = ~ ( n255 ) ;
assign n257 = ~ ( n75 ) ;
assign n258 =  ( n256 ) ^ ( n257 )  ;
assign n259 =  ( n258 ) ^ ( n100 )  ;
assign n260 = ~ ( n259 ) ;
assign n261 =  ( n252 ) | ( n260 )  ;
assign n262 = ~ ( n150 ) ;
assign n263 = ~ ( n160 ) ;
assign n264 =  ( n262 ) | ( n263 )  ;
assign n265 = ~ ( n75 ) ;
assign n266 =  ( n265 ) ^ ( n100 )  ;
assign n267 = ~ ( n266 ) ;
assign n268 =  ( n264 ) | ( n267 )  ;
assign n269 = ~ ( n268 ) ;
assign n270 =  ( bv_1_1_n2 ) ^ ( n269 )  ;
assign n271 = ~ ( n100 ) ;
assign n272 =  ( n75 ) | ( n271 )  ;
assign n273 = ~ ( n272 ) ;
assign n274 =  ( n270 ) ^ ( n273 )  ;
assign n275 =  ( n274 ) ^ ( n110 )  ;
assign n276 = ~ ( n275 ) ;
assign n277 =  ( n261 ) | ( n276 )  ;
assign n278 = ~ ( n150 ) ;
assign n279 = ~ ( n160 ) ;
assign n280 =  ( n278 ) | ( n279 )  ;
assign n281 = ~ ( n75 ) ;
assign n282 =  ( n281 ) ^ ( n100 )  ;
assign n283 = ~ ( n282 ) ;
assign n284 =  ( n280 ) | ( n283 )  ;
assign n285 = ~ ( n171 ) ;
assign n286 =  ( n284 ) | ( n285 )  ;
assign n287 = ~ ( n286 ) ;
assign n288 =  ( n287 ) ^ ( n118 )  ;
assign n289 = ~ ( n110 ) ;
assign n290 =  ( n288 ) ^ ( n289 )  ;
assign n291 = ~ ( n290 ) ;
assign n292 =  ( n277 ) | ( n291 )  ;
assign n293 = ~ ( n292 ) ;
assign n294 = ~ ( n227 ) ;
assign n295 = ~ ( n247 ) ;
assign n296 =  ( n294 ) | ( n295 )  ;
assign n297 =  ( n150 ) ^ ( n160 )  ;
assign n298 = ~ ( n297 ) ;
assign n299 =  ( n296 ) | ( n298 )  ;
assign n300 = ~ ( n259 ) ;
assign n301 =  ( n299 ) | ( n300 )  ;
assign n302 = ~ ( n275 ) ;
assign n303 =  ( n301 ) | ( n302 )  ;
assign n304 = ~ ( n303 ) ;
assign n305 = ~ ( n286 ) ;
assign n306 =  ( n304 ) ^ ( n305 )  ;
assign n307 =  ( n306 ) ^ ( n118 )  ;
assign n308 = ~ ( n110 ) ;
assign n309 =  ( n307 ) ^ ( n308 )  ;
assign n310 = ~ ( n309 ) ;
assign n311 = ki[0:0] ;
assign n312 =  ( n311 ) == ( bv_1_1_n2 )  ;
assign n313 = ki[1:1] ;
assign n314 =  ( n313 ) == ( bv_1_0_n74 )  ;
assign n315 =  ( n312 ) | ( n314 )  ;
assign n316 = ki[1:1] ;
assign n317 =  ( n316 ) == ( bv_1_1_n2 )  ;
assign n318 = ki[0:0] ;
assign n319 =  ( n318 ) == ( bv_1_1_n2 )  ;
assign n320 =  ( n317 ) | ( n319 )  ;
assign n321 = ki[1:1] ;
assign n322 =  ( n321 ) == ( bv_1_1_n2 )  ;
assign n323 = i_wb_data[1:1] ;
assign n324 = ~ ( n323 ) ;
assign n325 = sp[1:1] ;
assign n326 =  ( n324 ) ^ ( n325 )  ;
assign n327 =  ( n326 ) ^ ( n245 )  ;
assign n328 = ~ ( n327 ) ;
assign n329 = i_wb_data[1:1] ;
assign n330 = ~ ( n329 ) ;
assign n331 = sp[1:1] ;
assign n332 =  ( n330 ) ^ ( n331 )  ;
assign n333 =  ( n332 ) ^ ( n245 )  ;
assign n334 =  ( n322 ) ? ( n328 ) : ( n333 ) ;
assign n335 =  ( n320 ) ? ( n334 ) : ( bv_1_0_n74 ) ;
assign n336 =  ( n315 ) ? ( n226 ) : ( n335 ) ;
assign n337 = ~ ( n336 ) ;
assign n338 = ki[1:1] ;
assign n339 =  ( n338 ) == ( bv_1_0_n74 )  ;
assign n340 = i_wb_data[1:1] ;
assign n341 = ~ ( n340 ) ;
assign n342 = sp[1:1] ;
assign n343 =  ( n341 ) ^ ( n342 )  ;
assign n344 =  ( n343 ) ^ ( n241 )  ;
assign n345 =  ( n339 ) ? ( bv_1_0_n74 ) : ( n344 ) ;
assign n346 = ~ ( n345 ) ;
assign n347 =  ( n337 ) | ( n346 )  ;
assign n348 =  ( n227 ) ^ ( n247 )  ;
assign n349 = ~ ( n348 ) ;
assign n350 =  ( n347 ) | ( n349 )  ;
assign n351 = ~ ( n227 ) ;
assign n352 = ~ ( n247 ) ;
assign n353 =  ( n351 ) | ( n352 )  ;
assign n354 = ~ ( n353 ) ;
assign n355 =  ( n354 ) ^ ( n150 )  ;
assign n356 =  ( n355 ) ^ ( n160 )  ;
assign n357 = ~ ( n356 ) ;
assign n358 =  ( n350 ) | ( n357 )  ;
assign n359 = ~ ( n227 ) ;
assign n360 = ~ ( n247 ) ;
assign n361 =  ( n359 ) | ( n360 )  ;
assign n362 =  ( n150 ) ^ ( n160 )  ;
assign n363 = ~ ( n362 ) ;
assign n364 =  ( n361 ) | ( n363 )  ;
assign n365 = ~ ( n364 ) ;
assign n366 = ~ ( n150 ) ;
assign n367 = ~ ( n160 ) ;
assign n368 =  ( n366 ) | ( n367 )  ;
assign n369 = ~ ( n368 ) ;
assign n370 =  ( n365 ) ^ ( n369 )  ;
assign n371 = ~ ( n75 ) ;
assign n372 =  ( n370 ) ^ ( n371 )  ;
assign n373 =  ( n372 ) ^ ( n100 )  ;
assign n374 = ~ ( n373 ) ;
assign n375 =  ( n358 ) | ( n374 )  ;
assign n376 = ~ ( n375 ) ;
assign n377 = ~ ( n336 ) ;
assign n378 = ~ ( n345 ) ;
assign n379 =  ( n377 ) | ( n378 )  ;
assign n380 =  ( n227 ) ^ ( n247 )  ;
assign n381 = ~ ( n380 ) ;
assign n382 =  ( n379 ) | ( n381 )  ;
assign n383 = ~ ( n356 ) ;
assign n384 =  ( n382 ) | ( n383 )  ;
assign n385 = ~ ( n384 ) ;
assign n386 =  ( n385 ) ^ ( n365 )  ;
assign n387 = ~ ( n150 ) ;
assign n388 = ~ ( n160 ) ;
assign n389 =  ( n387 ) | ( n388 )  ;
assign n390 = ~ ( n389 ) ;
assign n391 =  ( n386 ) ^ ( n390 )  ;
assign n392 = ~ ( n75 ) ;
assign n393 =  ( n391 ) ^ ( n392 )  ;
assign n394 =  ( n393 ) ^ ( n100 )  ;
assign n395 =  ( n376 ) | ( n394 )  ;
assign n396 = ~ ( n395 ) ;
assign n397 =  ( n310 ) | ( n396 )  ;
assign n398 = ~ ( n227 ) ;
assign n399 = ~ ( n247 ) ;
assign n400 =  ( n398 ) | ( n399 )  ;
assign n401 =  ( n150 ) ^ ( n160 )  ;
assign n402 = ~ ( n401 ) ;
assign n403 =  ( n400 ) | ( n402 )  ;
assign n404 = ~ ( n259 ) ;
assign n405 =  ( n403 ) | ( n404 )  ;
assign n406 = ~ ( n405 ) ;
assign n407 =  ( bv_1_1_n2 ) ^ ( n406 )  ;
assign n408 = ~ ( n268 ) ;
assign n409 =  ( n407 ) ^ ( n408 )  ;
assign n410 = ~ ( n100 ) ;
assign n411 =  ( n75 ) | ( n410 )  ;
assign n412 = ~ ( n411 ) ;
assign n413 =  ( n409 ) ^ ( n412 )  ;
assign n414 =  ( n413 ) ^ ( n110 )  ;
assign n415 = ~ ( n414 ) ;
assign n416 =  ( n397 ) | ( n415 )  ;
assign n417 = ~ ( n416 ) ;
assign n418 =  ( n293 ) | ( n417 )  ;
assign n419 = ~ ( n286 ) ;
assign n420 =  ( n304 ) ^ ( n419 )  ;
assign n421 =  ( n420 ) ^ ( n118 )  ;
assign n422 = ~ ( n110 ) ;
assign n423 =  ( n421 ) ^ ( n422 )  ;
assign n424 = ~ ( n423 ) ;
assign n425 =  ( n376 ) | ( n394 )  ;
assign n426 =  ( bv_1_1_n2 ) ^ ( n425 )  ;
assign n427 =  ( n426 ) ^ ( n406 )  ;
assign n428 = ~ ( n268 ) ;
assign n429 =  ( n427 ) ^ ( n428 )  ;
assign n430 = ~ ( n100 ) ;
assign n431 =  ( n75 ) | ( n430 )  ;
assign n432 = ~ ( n431 ) ;
assign n433 =  ( n429 ) ^ ( n432 )  ;
assign n434 =  ( n433 ) ^ ( n110 )  ;
assign n435 = ~ ( n434 ) ;
assign n436 =  ( n424 ) | ( n435 )  ;
assign n437 = ki[0:0] ;
assign n438 =  ( n437 ) == ( bv_1_1_n2 )  ;
assign n439 = ki[1:1] ;
assign n440 =  ( n439 ) == ( bv_1_0_n74 )  ;
assign n441 =  ( n438 ) | ( n440 )  ;
assign n442 = ki[1:1] ;
assign n443 =  ( n442 ) == ( bv_1_1_n2 )  ;
assign n444 = ki[0:0] ;
assign n445 =  ( n444 ) == ( bv_1_1_n2 )  ;
assign n446 =  ( n443 ) | ( n445 )  ;
assign n447 = ki[1:1] ;
assign n448 =  ( n447 ) == ( bv_1_1_n2 )  ;
assign n449 = i_wb_data[1:1] ;
assign n450 = ~ ( n449 ) ;
assign n451 = sp[1:1] ;
assign n452 =  ( n450 ) ^ ( n451 )  ;
assign n453 =  ( n452 ) ^ ( n241 )  ;
assign n454 = ~ ( n453 ) ;
assign n455 = i_wb_data[1:1] ;
assign n456 = ~ ( n455 ) ;
assign n457 = sp[1:1] ;
assign n458 =  ( n456 ) ^ ( n457 )  ;
assign n459 =  ( n458 ) ^ ( n241 )  ;
assign n460 =  ( n448 ) ? ( n454 ) : ( n459 ) ;
assign n461 =  ( n446 ) ? ( n460 ) : ( bv_1_0_n74 ) ;
assign n462 =  ( n441 ) ? ( n335 ) : ( n461 ) ;
assign n463 = ~ ( n462 ) ;
assign n464 = ki[1:1] ;
assign n465 =  ( n464 ) == ( bv_1_0_n74 )  ;
assign n466 = i_wb_data[1:1] ;
assign n467 = ~ ( n466 ) ;
assign n468 = sp[1:1] ;
assign n469 =  ( n467 ) ^ ( n468 )  ;
assign n470 =  ( n17 ) | ( n28 )  ;
assign n471 =  ( n470 ) | ( n33 )  ;
assign n472 =  ( n471 ) | ( n39 )  ;
assign n473 = ~ ( n53 ) ;
assign n474 =  ( n22 ) | ( n473 )  ;
assign n475 = ~ ( n474 ) ;
assign n476 =  ( n472 ) | ( n475 )  ;
assign n477 = ~ ( n476 ) ;
assign n478 =  ( n22 ) | ( n477 )  ;
assign n479 = ~ ( n478 ) ;
assign n480 =  ( n17 ) | ( n479 )  ;
assign n481 =  ( n469 ) ^ ( n480 )  ;
assign n482 =  ( n465 ) ? ( bv_1_0_n74 ) : ( n481 ) ;
assign n483 = ~ ( n482 ) ;
assign n484 =  ( n463 ) | ( n483 )  ;
assign n485 =  ( n336 ) ^ ( n345 )  ;
assign n486 = ~ ( n485 ) ;
assign n487 =  ( n484 ) | ( n486 )  ;
assign n488 = ~ ( n336 ) ;
assign n489 = ~ ( n345 ) ;
assign n490 =  ( n488 ) | ( n489 )  ;
assign n491 = ~ ( n490 ) ;
assign n492 =  ( n491 ) ^ ( n227 )  ;
assign n493 =  ( n492 ) ^ ( n247 )  ;
assign n494 = ~ ( n493 ) ;
assign n495 =  ( n487 ) | ( n494 )  ;
assign n496 = ~ ( n336 ) ;
assign n497 = ~ ( n345 ) ;
assign n498 =  ( n496 ) | ( n497 )  ;
assign n499 =  ( n227 ) ^ ( n247 )  ;
assign n500 = ~ ( n499 ) ;
assign n501 =  ( n498 ) | ( n500 )  ;
assign n502 = ~ ( n501 ) ;
assign n503 = ~ ( n227 ) ;
assign n504 = ~ ( n247 ) ;
assign n505 =  ( n503 ) | ( n504 )  ;
assign n506 = ~ ( n505 ) ;
assign n507 =  ( n502 ) ^ ( n506 )  ;
assign n508 =  ( n507 ) ^ ( n150 )  ;
assign n509 =  ( n508 ) ^ ( n160 )  ;
assign n510 = ~ ( n509 ) ;
assign n511 =  ( n495 ) | ( n510 )  ;
assign n512 =  ( bv_1_1_n2 ) ^ ( n385 )  ;
assign n513 =  ( n512 ) ^ ( n365 )  ;
assign n514 = ~ ( n150 ) ;
assign n515 = ~ ( n160 ) ;
assign n516 =  ( n514 ) | ( n515 )  ;
assign n517 = ~ ( n516 ) ;
assign n518 =  ( n513 ) ^ ( n517 )  ;
assign n519 = ~ ( n75 ) ;
assign n520 =  ( n518 ) ^ ( n519 )  ;
assign n521 =  ( n520 ) ^ ( n100 )  ;
assign n522 = ~ ( n521 ) ;
assign n523 =  ( n511 ) | ( n522 )  ;
assign n524 = ~ ( n523 ) ;
assign n525 = ~ ( n462 ) ;
assign n526 = ~ ( n482 ) ;
assign n527 =  ( n525 ) | ( n526 )  ;
assign n528 =  ( n336 ) ^ ( n345 )  ;
assign n529 = ~ ( n528 ) ;
assign n530 =  ( n527 ) | ( n529 )  ;
assign n531 = ~ ( n493 ) ;
assign n532 =  ( n530 ) | ( n531 )  ;
assign n533 = ~ ( n509 ) ;
assign n534 =  ( n532 ) | ( n533 )  ;
assign n535 = ~ ( n534 ) ;
assign n536 =  ( bv_1_1_n2 ) ^ ( n535 )  ;
assign n537 =  ( n536 ) ^ ( n385 )  ;
assign n538 =  ( n537 ) ^ ( n365 )  ;
assign n539 = ~ ( n150 ) ;
assign n540 = ~ ( n160 ) ;
assign n541 =  ( n539 ) | ( n540 )  ;
assign n542 = ~ ( n541 ) ;
assign n543 =  ( n538 ) ^ ( n542 )  ;
assign n544 = ~ ( n75 ) ;
assign n545 =  ( n543 ) ^ ( n544 )  ;
assign n546 =  ( n545 ) ^ ( n100 )  ;
assign n547 = ~ ( n546 ) ;
assign n548 = ki[0:0] ;
assign n549 =  ( n548 ) == ( bv_1_1_n2 )  ;
assign n550 = ki[1:1] ;
assign n551 =  ( n550 ) == ( bv_1_0_n74 )  ;
assign n552 =  ( n549 ) | ( n551 )  ;
assign n553 = ki[1:1] ;
assign n554 =  ( n553 ) == ( bv_1_1_n2 )  ;
assign n555 = ki[0:0] ;
assign n556 =  ( n555 ) == ( bv_1_1_n2 )  ;
assign n557 =  ( n554 ) | ( n556 )  ;
assign n558 = ki[1:1] ;
assign n559 =  ( n558 ) == ( bv_1_1_n2 )  ;
assign n560 = i_wb_data[1:1] ;
assign n561 = ~ ( n560 ) ;
assign n562 = sp[1:1] ;
assign n563 =  ( n561 ) ^ ( n562 )  ;
assign n564 =  ( n563 ) ^ ( n480 )  ;
assign n565 = ~ ( n564 ) ;
assign n566 = i_wb_data[1:1] ;
assign n567 = ~ ( n566 ) ;
assign n568 = sp[1:1] ;
assign n569 =  ( n567 ) ^ ( n568 )  ;
assign n570 =  ( n569 ) ^ ( n480 )  ;
assign n571 =  ( n559 ) ? ( n565 ) : ( n570 ) ;
assign n572 =  ( n557 ) ? ( n571 ) : ( bv_1_0_n74 ) ;
assign n573 =  ( n552 ) ? ( n461 ) : ( n572 ) ;
assign n574 = ~ ( n573 ) ;
assign n575 =  ( n547 ) | ( n574 )  ;
assign n576 = ki[1:1] ;
assign n577 =  ( n576 ) == ( bv_1_0_n74 )  ;
assign n578 = i_wb_data[1:1] ;
assign n579 = ~ ( n578 ) ;
assign n580 = sp[1:1] ;
assign n581 =  ( n579 ) ^ ( n580 )  ;
assign n582 =  ( n581 ) ^ ( n476 )  ;
assign n583 =  ( n577 ) ? ( bv_1_0_n74 ) : ( n582 ) ;
assign n584 = ~ ( n583 ) ;
assign n585 =  ( n575 ) | ( n584 )  ;
assign n586 =  ( n462 ) ^ ( n482 )  ;
assign n587 = ~ ( n586 ) ;
assign n588 =  ( n585 ) | ( n587 )  ;
assign n589 = ~ ( n462 ) ;
assign n590 = ~ ( n482 ) ;
assign n591 =  ( n589 ) | ( n590 )  ;
assign n592 = ~ ( n591 ) ;
assign n593 =  ( n592 ) ^ ( n336 )  ;
assign n594 =  ( n593 ) ^ ( n345 )  ;
assign n595 = ~ ( n594 ) ;
assign n596 =  ( n588 ) | ( n595 )  ;
assign n597 = ~ ( n462 ) ;
assign n598 = ~ ( n482 ) ;
assign n599 =  ( n597 ) | ( n598 )  ;
assign n600 =  ( n336 ) ^ ( n345 )  ;
assign n601 = ~ ( n600 ) ;
assign n602 =  ( n599 ) | ( n601 )  ;
assign n603 = ~ ( n602 ) ;
assign n604 = ~ ( n336 ) ;
assign n605 = ~ ( n345 ) ;
assign n606 =  ( n604 ) | ( n605 )  ;
assign n607 = ~ ( n606 ) ;
assign n608 =  ( n603 ) ^ ( n607 )  ;
assign n609 =  ( n608 ) ^ ( n227 )  ;
assign n610 =  ( n609 ) ^ ( n247 )  ;
assign n611 = ~ ( n610 ) ;
assign n612 =  ( n596 ) | ( n611 )  ;
assign n613 = ~ ( n462 ) ;
assign n614 = ~ ( n482 ) ;
assign n615 =  ( n613 ) | ( n614 )  ;
assign n616 =  ( n336 ) ^ ( n345 )  ;
assign n617 = ~ ( n616 ) ;
assign n618 =  ( n615 ) | ( n617 )  ;
assign n619 = ~ ( n493 ) ;
assign n620 =  ( n618 ) | ( n619 )  ;
assign n621 = ~ ( n620 ) ;
assign n622 =  ( n621 ) ^ ( n502 )  ;
assign n623 = ~ ( n227 ) ;
assign n624 = ~ ( n247 ) ;
assign n625 =  ( n623 ) | ( n624 )  ;
assign n626 = ~ ( n625 ) ;
assign n627 =  ( n622 ) ^ ( n626 )  ;
assign n628 =  ( n627 ) ^ ( n150 )  ;
assign n629 =  ( n628 ) ^ ( n160 )  ;
assign n630 = ~ ( n629 ) ;
assign n631 =  ( n612 ) | ( n630 )  ;
assign n632 = ~ ( n631 ) ;
assign n633 =  ( n524 ) | ( n632 )  ;
assign n634 = ~ ( n633 ) ;
assign n635 =  ( n436 ) | ( n634 )  ;
assign n636 = ~ ( n635 ) ;
assign n637 =  ( n418 ) | ( n636 )  ;
assign n638 = ~ ( n637 ) ;
assign n639 =  ( n201 ) | ( n638 )  ;
assign n640 = ~ ( n639 ) ;
assign n641 =  ( n179 ) | ( n640 )  ;
assign n642 = ~ ( n118 ) ;
assign n643 =  ( n642 ) | ( n110 )  ;
assign n644 = ~ ( n643 ) ;
assign n645 =  ( n644 ) | ( n200 )  ;
assign n646 = ~ ( n286 ) ;
assign n647 =  ( n304 ) ^ ( n646 )  ;
assign n648 =  ( n647 ) ^ ( n118 )  ;
assign n649 = ~ ( n110 ) ;
assign n650 =  ( n648 ) ^ ( n649 )  ;
assign n651 = ~ ( n650 ) ;
assign n652 =  ( n645 ) | ( n651 )  ;
assign n653 = ~ ( n434 ) ;
assign n654 =  ( n652 ) | ( n653 )  ;
assign n655 = ~ ( n546 ) ;
assign n656 =  ( n654 ) | ( n655 )  ;
assign n657 = ~ ( n573 ) ;
assign n658 = ~ ( n583 ) ;
assign n659 =  ( n657 ) | ( n658 )  ;
assign n660 =  ( n462 ) ^ ( n482 )  ;
assign n661 = ~ ( n660 ) ;
assign n662 =  ( n659 ) | ( n661 )  ;
assign n663 = ~ ( n594 ) ;
assign n664 =  ( n662 ) | ( n663 )  ;
assign n665 = ~ ( n610 ) ;
assign n666 =  ( n664 ) | ( n665 )  ;
assign n667 = ~ ( n666 ) ;
assign n668 =  ( n667 ) ^ ( n621 )  ;
assign n669 =  ( n668 ) ^ ( n502 )  ;
assign n670 = ~ ( n227 ) ;
assign n671 = ~ ( n247 ) ;
assign n672 =  ( n670 ) | ( n671 )  ;
assign n673 = ~ ( n672 ) ;
assign n674 =  ( n669 ) ^ ( n673 )  ;
assign n675 =  ( n674 ) ^ ( n150 )  ;
assign n676 =  ( n675 ) ^ ( n160 )  ;
assign n677 = ~ ( n676 ) ;
assign n678 =  ( n656 ) | ( n677 )  ;
assign n679 = ki[0:0] ;
assign n680 =  ( n679 ) == ( bv_1_1_n2 )  ;
assign n681 = ki[1:1] ;
assign n682 =  ( n681 ) == ( bv_1_0_n74 )  ;
assign n683 =  ( n680 ) | ( n682 )  ;
assign n684 = ki[1:1] ;
assign n685 =  ( n684 ) == ( bv_1_1_n2 )  ;
assign n686 = ki[0:0] ;
assign n687 =  ( n686 ) == ( bv_1_1_n2 )  ;
assign n688 =  ( n685 ) | ( n687 )  ;
assign n689 = ki[1:1] ;
assign n690 =  ( n689 ) == ( bv_1_1_n2 )  ;
assign n691 = i_wb_data[1:1] ;
assign n692 = ~ ( n691 ) ;
assign n693 = sp[1:1] ;
assign n694 =  ( n692 ) ^ ( n693 )  ;
assign n695 =  ( n694 ) ^ ( n476 )  ;
assign n696 = ~ ( n695 ) ;
assign n697 = i_wb_data[1:1] ;
assign n698 = ~ ( n697 ) ;
assign n699 = sp[1:1] ;
assign n700 =  ( n698 ) ^ ( n699 )  ;
assign n701 =  ( n700 ) ^ ( n476 )  ;
assign n702 =  ( n690 ) ? ( n696 ) : ( n701 ) ;
assign n703 =  ( n688 ) ? ( n702 ) : ( bv_1_0_n74 ) ;
assign n704 =  ( n683 ) ? ( n572 ) : ( n703 ) ;
assign n705 = ~ ( n704 ) ;
assign n706 = ki[1:1] ;
assign n707 =  ( n706 ) == ( bv_1_0_n74 )  ;
assign n708 = i_wb_data[1:1] ;
assign n709 = ~ ( n708 ) ;
assign n710 = sp[1:1] ;
assign n711 =  ( n709 ) ^ ( n710 )  ;
assign n712 = ~ ( n61 ) ;
assign n713 =  ( n22 ) | ( n712 )  ;
assign n714 = ~ ( n713 ) ;
assign n715 =  ( n17 ) | ( n714 )  ;
assign n716 =  ( n711 ) ^ ( n715 )  ;
assign n717 =  ( n707 ) ? ( bv_1_0_n74 ) : ( n716 ) ;
assign n718 = ~ ( n717 ) ;
assign n719 =  ( n705 ) | ( n718 )  ;
assign n720 =  ( n573 ) ^ ( n583 )  ;
assign n721 = ~ ( n720 ) ;
assign n722 =  ( n719 ) | ( n721 )  ;
assign n723 = ~ ( n573 ) ;
assign n724 = ~ ( n583 ) ;
assign n725 =  ( n723 ) | ( n724 )  ;
assign n726 = ~ ( n725 ) ;
assign n727 =  ( n726 ) ^ ( n462 )  ;
assign n728 =  ( n727 ) ^ ( n482 )  ;
assign n729 = ~ ( n728 ) ;
assign n730 =  ( n722 ) | ( n729 )  ;
assign n731 = ~ ( n573 ) ;
assign n732 = ~ ( n583 ) ;
assign n733 =  ( n731 ) | ( n732 )  ;
assign n734 =  ( n462 ) ^ ( n482 )  ;
assign n735 = ~ ( n734 ) ;
assign n736 =  ( n733 ) | ( n735 )  ;
assign n737 = ~ ( n736 ) ;
assign n738 = ~ ( n462 ) ;
assign n739 = ~ ( n482 ) ;
assign n740 =  ( n738 ) | ( n739 )  ;
assign n741 = ~ ( n740 ) ;
assign n742 =  ( n737 ) ^ ( n741 )  ;
assign n743 =  ( n742 ) ^ ( n336 )  ;
assign n744 =  ( n743 ) ^ ( n345 )  ;
assign n745 = ~ ( n744 ) ;
assign n746 =  ( n730 ) | ( n745 )  ;
assign n747 = ~ ( n573 ) ;
assign n748 = ~ ( n583 ) ;
assign n749 =  ( n747 ) | ( n748 )  ;
assign n750 =  ( n462 ) ^ ( n482 )  ;
assign n751 = ~ ( n750 ) ;
assign n752 =  ( n749 ) | ( n751 )  ;
assign n753 = ~ ( n594 ) ;
assign n754 =  ( n752 ) | ( n753 )  ;
assign n755 = ~ ( n754 ) ;
assign n756 =  ( n755 ) ^ ( n603 )  ;
assign n757 = ~ ( n336 ) ;
assign n758 = ~ ( n345 ) ;
assign n759 =  ( n757 ) | ( n758 )  ;
assign n760 = ~ ( n759 ) ;
assign n761 =  ( n756 ) ^ ( n760 )  ;
assign n762 =  ( n761 ) ^ ( n227 )  ;
assign n763 =  ( n762 ) ^ ( n247 )  ;
assign n764 = ~ ( n763 ) ;
assign n765 =  ( n746 ) | ( n764 )  ;
assign n766 = ~ ( n765 ) ;
assign n767 = ~ ( n704 ) ;
assign n768 = ~ ( n717 ) ;
assign n769 =  ( n767 ) | ( n768 )  ;
assign n770 =  ( n573 ) ^ ( n583 )  ;
assign n771 = ~ ( n770 ) ;
assign n772 =  ( n769 ) | ( n771 )  ;
assign n773 = ~ ( n728 ) ;
assign n774 =  ( n772 ) | ( n773 )  ;
assign n775 = ~ ( n744 ) ;
assign n776 =  ( n774 ) | ( n775 )  ;
assign n777 = ~ ( n776 ) ;
assign n778 =  ( n777 ) ^ ( n755 )  ;
assign n779 =  ( n778 ) ^ ( n603 )  ;
assign n780 = ~ ( n336 ) ;
assign n781 = ~ ( n345 ) ;
assign n782 =  ( n780 ) | ( n781 )  ;
assign n783 = ~ ( n782 ) ;
assign n784 =  ( n779 ) ^ ( n783 )  ;
assign n785 =  ( n784 ) ^ ( n227 )  ;
assign n786 =  ( n785 ) ^ ( n247 )  ;
assign n787 = ~ ( n786 ) ;
assign n788 = ki[0:0] ;
assign n789 =  ( n788 ) == ( bv_1_1_n2 )  ;
assign n790 = ki[1:1] ;
assign n791 =  ( n790 ) == ( bv_1_0_n74 )  ;
assign n792 =  ( n789 ) | ( n791 )  ;
assign n793 = ki[1:1] ;
assign n794 =  ( n793 ) == ( bv_1_1_n2 )  ;
assign n795 = ki[0:0] ;
assign n796 =  ( n795 ) == ( bv_1_1_n2 )  ;
assign n797 =  ( n794 ) | ( n796 )  ;
assign n798 = ki[1:1] ;
assign n799 =  ( n798 ) == ( bv_1_1_n2 )  ;
assign n800 = i_wb_data[1:1] ;
assign n801 = ~ ( n800 ) ;
assign n802 = sp[1:1] ;
assign n803 =  ( n801 ) ^ ( n802 )  ;
assign n804 =  ( n803 ) ^ ( n715 )  ;
assign n805 = ~ ( n804 ) ;
assign n806 = i_wb_data[1:1] ;
assign n807 = ~ ( n806 ) ;
assign n808 = sp[1:1] ;
assign n809 =  ( n807 ) ^ ( n808 )  ;
assign n810 =  ( n809 ) ^ ( n715 )  ;
assign n811 =  ( n799 ) ? ( n805 ) : ( n810 ) ;
assign n812 =  ( n797 ) ? ( n811 ) : ( bv_1_0_n74 ) ;
assign n813 =  ( n792 ) ? ( n703 ) : ( n812 ) ;
assign n814 = ~ ( n813 ) ;
assign n815 =  ( n787 ) | ( n814 )  ;
assign n816 = ki[1:1] ;
assign n817 =  ( n816 ) == ( bv_1_0_n74 )  ;
assign n818 = i_wb_data[1:1] ;
assign n819 = ~ ( n818 ) ;
assign n820 = sp[1:1] ;
assign n821 =  ( n819 ) ^ ( n820 )  ;
assign n822 =  ( n821 ) ^ ( n61 )  ;
assign n823 =  ( n817 ) ? ( bv_1_0_n74 ) : ( n822 ) ;
assign n824 = ~ ( n823 ) ;
assign n825 =  ( n815 ) | ( n824 )  ;
assign n826 =  ( n704 ) ^ ( n717 )  ;
assign n827 = ~ ( n826 ) ;
assign n828 =  ( n825 ) | ( n827 )  ;
assign n829 = ~ ( n704 ) ;
assign n830 = ~ ( n717 ) ;
assign n831 =  ( n829 ) | ( n830 )  ;
assign n832 = ~ ( n831 ) ;
assign n833 =  ( n832 ) ^ ( n573 )  ;
assign n834 =  ( n833 ) ^ ( n583 )  ;
assign n835 = ~ ( n834 ) ;
assign n836 =  ( n828 ) | ( n835 )  ;
assign n837 = ~ ( n704 ) ;
assign n838 = ~ ( n717 ) ;
assign n839 =  ( n837 ) | ( n838 )  ;
assign n840 =  ( n573 ) ^ ( n583 )  ;
assign n841 = ~ ( n840 ) ;
assign n842 =  ( n839 ) | ( n841 )  ;
assign n843 = ~ ( n842 ) ;
assign n844 = ~ ( n573 ) ;
assign n845 = ~ ( n583 ) ;
assign n846 =  ( n844 ) | ( n845 )  ;
assign n847 = ~ ( n846 ) ;
assign n848 =  ( n843 ) ^ ( n847 )  ;
assign n849 =  ( n848 ) ^ ( n462 )  ;
assign n850 =  ( n849 ) ^ ( n482 )  ;
assign n851 = ~ ( n850 ) ;
assign n852 =  ( n836 ) | ( n851 )  ;
assign n853 = ~ ( n704 ) ;
assign n854 = ~ ( n717 ) ;
assign n855 =  ( n853 ) | ( n854 )  ;
assign n856 =  ( n573 ) ^ ( n583 )  ;
assign n857 = ~ ( n856 ) ;
assign n858 =  ( n855 ) | ( n857 )  ;
assign n859 = ~ ( n728 ) ;
assign n860 =  ( n858 ) | ( n859 )  ;
assign n861 = ~ ( n860 ) ;
assign n862 =  ( n861 ) ^ ( n737 )  ;
assign n863 = ~ ( n462 ) ;
assign n864 = ~ ( n482 ) ;
assign n865 =  ( n863 ) | ( n864 )  ;
assign n866 = ~ ( n865 ) ;
assign n867 =  ( n862 ) ^ ( n866 )  ;
assign n868 =  ( n867 ) ^ ( n336 )  ;
assign n869 =  ( n868 ) ^ ( n345 )  ;
assign n870 = ~ ( n869 ) ;
assign n871 =  ( n852 ) | ( n870 )  ;
assign n872 = ~ ( n871 ) ;
assign n873 =  ( n766 ) | ( n872 )  ;
assign n874 = ~ ( n786 ) ;
assign n875 = ~ ( n813 ) ;
assign n876 = ~ ( n823 ) ;
assign n877 =  ( n875 ) | ( n876 )  ;
assign n878 =  ( n704 ) ^ ( n717 )  ;
assign n879 = ~ ( n878 ) ;
assign n880 =  ( n877 ) | ( n879 )  ;
assign n881 = ~ ( n834 ) ;
assign n882 =  ( n880 ) | ( n881 )  ;
assign n883 = ~ ( n850 ) ;
assign n884 =  ( n882 ) | ( n883 )  ;
assign n885 = ~ ( n884 ) ;
assign n886 =  ( n885 ) ^ ( n861 )  ;
assign n887 =  ( n886 ) ^ ( n737 )  ;
assign n888 = ~ ( n462 ) ;
assign n889 = ~ ( n482 ) ;
assign n890 =  ( n888 ) | ( n889 )  ;
assign n891 = ~ ( n890 ) ;
assign n892 =  ( n887 ) ^ ( n891 )  ;
assign n893 =  ( n892 ) ^ ( n336 )  ;
assign n894 =  ( n893 ) ^ ( n345 )  ;
assign n895 = ~ ( n894 ) ;
assign n896 =  ( n874 ) | ( n895 )  ;
assign n897 = ~ ( n813 ) ;
assign n898 = ~ ( n823 ) ;
assign n899 =  ( n897 ) | ( n898 )  ;
assign n900 =  ( n704 ) ^ ( n717 )  ;
assign n901 = ~ ( n900 ) ;
assign n902 =  ( n899 ) | ( n901 )  ;
assign n903 = ~ ( n834 ) ;
assign n904 =  ( n902 ) | ( n903 )  ;
assign n905 = ~ ( n904 ) ;
assign n906 =  ( n905 ) ^ ( n843 )  ;
assign n907 = ~ ( n573 ) ;
assign n908 = ~ ( n583 ) ;
assign n909 =  ( n907 ) | ( n908 )  ;
assign n910 = ~ ( n909 ) ;
assign n911 =  ( n906 ) ^ ( n910 )  ;
assign n912 =  ( n911 ) ^ ( n462 )  ;
assign n913 =  ( n912 ) ^ ( n482 )  ;
assign n914 = ~ ( n913 ) ;
assign n915 =  ( n896 ) | ( n914 )  ;
assign n916 = ki[0:0] ;
assign n917 =  ( n916 ) == ( bv_1_1_n2 )  ;
assign n918 = ki[1:1] ;
assign n919 =  ( n918 ) == ( bv_1_0_n74 )  ;
assign n920 =  ( n917 ) | ( n919 )  ;
assign n921 = ki[1:1] ;
assign n922 =  ( n921 ) == ( bv_1_1_n2 )  ;
assign n923 = ki[0:0] ;
assign n924 =  ( n923 ) == ( bv_1_1_n2 )  ;
assign n925 =  ( n922 ) | ( n924 )  ;
assign n926 = ki[1:1] ;
assign n927 =  ( n926 ) == ( bv_1_1_n2 )  ;
assign n928 = i_wb_data[1:1] ;
assign n929 = ~ ( n928 ) ;
assign n930 = sp[1:1] ;
assign n931 =  ( n929 ) ^ ( n930 )  ;
assign n932 =  ( n931 ) ^ ( n61 )  ;
assign n933 = ~ ( n932 ) ;
assign n934 = i_wb_data[1:1] ;
assign n935 = ~ ( n934 ) ;
assign n936 = sp[1:1] ;
assign n937 =  ( n935 ) ^ ( n936 )  ;
assign n938 =  ( n937 ) ^ ( n61 )  ;
assign n939 =  ( n927 ) ? ( n933 ) : ( n938 ) ;
assign n940 =  ( n925 ) ? ( n939 ) : ( bv_1_0_n74 ) ;
assign n941 =  ( n920 ) ? ( n812 ) : ( n940 ) ;
assign n942 = ~ ( n941 ) ;
assign n943 =  ( n915 ) | ( n942 )  ;
assign n944 = ki[1:1] ;
assign n945 =  ( n944 ) == ( bv_1_0_n74 )  ;
assign n946 = i_wb_data[1:1] ;
assign n947 = ~ ( n946 ) ;
assign n948 = sp[1:1] ;
assign n949 =  ( n947 ) ^ ( n948 )  ;
assign n950 = ~ ( n90 ) ;
assign n951 =  ( n22 ) | ( n950 )  ;
assign n952 = ~ ( n951 ) ;
assign n953 =  ( n17 ) | ( n952 )  ;
assign n954 =  ( n949 ) ^ ( n953 )  ;
assign n955 =  ( n945 ) ? ( bv_1_0_n74 ) : ( n954 ) ;
assign n956 = ~ ( n955 ) ;
assign n957 =  ( n943 ) | ( n956 )  ;
assign n958 =  ( n813 ) ^ ( n823 )  ;
assign n959 = ~ ( n958 ) ;
assign n960 =  ( n957 ) | ( n959 )  ;
assign n961 = ~ ( n813 ) ;
assign n962 = ~ ( n823 ) ;
assign n963 =  ( n961 ) | ( n962 )  ;
assign n964 = ~ ( n963 ) ;
assign n965 =  ( n964 ) ^ ( n704 )  ;
assign n966 =  ( n965 ) ^ ( n717 )  ;
assign n967 = ~ ( n966 ) ;
assign n968 =  ( n960 ) | ( n967 )  ;
assign n969 = ~ ( n813 ) ;
assign n970 = ~ ( n823 ) ;
assign n971 =  ( n969 ) | ( n970 )  ;
assign n972 =  ( n704 ) ^ ( n717 )  ;
assign n973 = ~ ( n972 ) ;
assign n974 =  ( n971 ) | ( n973 )  ;
assign n975 = ~ ( n974 ) ;
assign n976 = ~ ( n704 ) ;
assign n977 = ~ ( n717 ) ;
assign n978 =  ( n976 ) | ( n977 )  ;
assign n979 = ~ ( n978 ) ;
assign n980 =  ( n975 ) ^ ( n979 )  ;
assign n981 =  ( n980 ) ^ ( n573 )  ;
assign n982 =  ( n981 ) ^ ( n583 )  ;
assign n983 = ~ ( n982 ) ;
assign n984 =  ( n968 ) | ( n983 )  ;
assign n985 = ~ ( n984 ) ;
assign n986 =  ( n873 ) | ( n985 )  ;
assign n987 = ~ ( n786 ) ;
assign n988 = ~ ( n894 ) ;
assign n989 =  ( n987 ) | ( n988 )  ;
assign n990 = ~ ( n913 ) ;
assign n991 =  ( n989 ) | ( n990 )  ;
assign n992 = ~ ( n941 ) ;
assign n993 = ~ ( n955 ) ;
assign n994 =  ( n992 ) | ( n993 )  ;
assign n995 =  ( n813 ) ^ ( n823 )  ;
assign n996 = ~ ( n995 ) ;
assign n997 =  ( n994 ) | ( n996 )  ;
assign n998 = ~ ( n966 ) ;
assign n999 =  ( n997 ) | ( n998 )  ;
assign n1000 = ~ ( n999 ) ;
assign n1001 =  ( n1000 ) ^ ( n975 )  ;
assign n1002 = ~ ( n704 ) ;
assign n1003 = ~ ( n717 ) ;
assign n1004 =  ( n1002 ) | ( n1003 )  ;
assign n1005 = ~ ( n1004 ) ;
assign n1006 =  ( n1001 ) ^ ( n1005 )  ;
assign n1007 =  ( n1006 ) ^ ( n573 )  ;
assign n1008 =  ( n1007 ) ^ ( n583 )  ;
assign n1009 = ~ ( n1008 ) ;
assign n1010 =  ( n991 ) | ( n1009 )  ;
assign n1011 = ki[0:0] ;
assign n1012 =  ( n1011 ) == ( bv_1_1_n2 )  ;
assign n1013 = ki[1:1] ;
assign n1014 =  ( n1013 ) == ( bv_1_0_n74 )  ;
assign n1015 =  ( n1012 ) | ( n1014 )  ;
assign n1016 = ki[1:1] ;
assign n1017 =  ( n1016 ) == ( bv_1_1_n2 )  ;
assign n1018 = ki[0:0] ;
assign n1019 =  ( n1018 ) == ( bv_1_1_n2 )  ;
assign n1020 =  ( n1017 ) | ( n1019 )  ;
assign n1021 = ki[1:1] ;
assign n1022 =  ( n1021 ) == ( bv_1_1_n2 )  ;
assign n1023 = i_wb_data[1:1] ;
assign n1024 = ~ ( n1023 ) ;
assign n1025 = sp[1:1] ;
assign n1026 =  ( n1024 ) ^ ( n1025 )  ;
assign n1027 =  ( n1026 ) ^ ( n953 )  ;
assign n1028 = ~ ( n1027 ) ;
assign n1029 = i_wb_data[1:1] ;
assign n1030 = ~ ( n1029 ) ;
assign n1031 = sp[1:1] ;
assign n1032 =  ( n1030 ) ^ ( n1031 )  ;
assign n1033 =  ( n1032 ) ^ ( n953 )  ;
assign n1034 =  ( n1022 ) ? ( n1028 ) : ( n1033 ) ;
assign n1035 =  ( n1020 ) ? ( n1034 ) : ( bv_1_0_n74 ) ;
assign n1036 =  ( n1015 ) ? ( n940 ) : ( n1035 ) ;
assign n1037 = ~ ( n1036 ) ;
assign n1038 = ki[1:1] ;
assign n1039 =  ( n1038 ) == ( bv_1_0_n74 )  ;
assign n1040 = i_wb_data[1:1] ;
assign n1041 = ~ ( n1040 ) ;
assign n1042 = sp[1:1] ;
assign n1043 =  ( n1041 ) ^ ( n1042 )  ;
assign n1044 =  ( n1043 ) ^ ( n90 )  ;
assign n1045 =  ( n1039 ) ? ( bv_1_0_n74 ) : ( n1044 ) ;
assign n1046 = ~ ( n1045 ) ;
assign n1047 =  ( n1037 ) | ( n1046 )  ;
assign n1048 =  ( n941 ) ^ ( n955 )  ;
assign n1049 = ~ ( n1048 ) ;
assign n1050 =  ( n1047 ) | ( n1049 )  ;
assign n1051 = ~ ( n941 ) ;
assign n1052 = ~ ( n955 ) ;
assign n1053 =  ( n1051 ) | ( n1052 )  ;
assign n1054 = ~ ( n1053 ) ;
assign n1055 =  ( n1054 ) ^ ( n813 )  ;
assign n1056 =  ( n1055 ) ^ ( n823 )  ;
assign n1057 = ~ ( n1056 ) ;
assign n1058 =  ( n1050 ) | ( n1057 )  ;
assign n1059 = ~ ( n941 ) ;
assign n1060 = ~ ( n955 ) ;
assign n1061 =  ( n1059 ) | ( n1060 )  ;
assign n1062 =  ( n813 ) ^ ( n823 )  ;
assign n1063 = ~ ( n1062 ) ;
assign n1064 =  ( n1061 ) | ( n1063 )  ;
assign n1065 = ~ ( n1064 ) ;
assign n1066 = ~ ( n813 ) ;
assign n1067 = ~ ( n823 ) ;
assign n1068 =  ( n1066 ) | ( n1067 )  ;
assign n1069 = ~ ( n1068 ) ;
assign n1070 =  ( n1065 ) ^ ( n1069 )  ;
assign n1071 =  ( n1070 ) ^ ( n704 )  ;
assign n1072 =  ( n1071 ) ^ ( n717 )  ;
assign n1073 = ~ ( n1072 ) ;
assign n1074 =  ( n1058 ) | ( n1073 )  ;
assign n1075 = ~ ( n1074 ) ;
assign n1076 = ~ ( n1036 ) ;
assign n1077 = ~ ( n1045 ) ;
assign n1078 =  ( n1076 ) | ( n1077 )  ;
assign n1079 =  ( n941 ) ^ ( n955 )  ;
assign n1080 = ~ ( n1079 ) ;
assign n1081 =  ( n1078 ) | ( n1080 )  ;
assign n1082 = ~ ( n1056 ) ;
assign n1083 =  ( n1081 ) | ( n1082 )  ;
assign n1084 = ~ ( n1083 ) ;
assign n1085 =  ( n1084 ) ^ ( n1065 )  ;
assign n1086 = ~ ( n813 ) ;
assign n1087 = ~ ( n823 ) ;
assign n1088 =  ( n1086 ) | ( n1087 )  ;
assign n1089 = ~ ( n1088 ) ;
assign n1090 =  ( n1085 ) ^ ( n1089 )  ;
assign n1091 =  ( n1090 ) ^ ( n704 )  ;
assign n1092 =  ( n1091 ) ^ ( n717 )  ;
assign n1093 = ~ ( n1092 ) ;
assign n1094 = ki[0:0] ;
assign n1095 =  ( n1094 ) == ( bv_1_1_n2 )  ;
assign n1096 = ki[1:1] ;
assign n1097 =  ( n1096 ) == ( bv_1_0_n74 )  ;
assign n1098 =  ( n1095 ) | ( n1097 )  ;
assign n1099 = ki[1:1] ;
assign n1100 =  ( n1099 ) == ( bv_1_1_n2 )  ;
assign n1101 = ki[0:0] ;
assign n1102 =  ( n1101 ) == ( bv_1_1_n2 )  ;
assign n1103 =  ( n1100 ) | ( n1102 )  ;
assign n1104 = ki[1:1] ;
assign n1105 =  ( n1104 ) == ( bv_1_1_n2 )  ;
assign n1106 = i_wb_data[1:1] ;
assign n1107 = ~ ( n1106 ) ;
assign n1108 = sp[1:1] ;
assign n1109 =  ( n1107 ) ^ ( n1108 )  ;
assign n1110 =  ( n1109 ) ^ ( n90 )  ;
assign n1111 = ~ ( n1110 ) ;
assign n1112 = i_wb_data[1:1] ;
assign n1113 = ~ ( n1112 ) ;
assign n1114 = sp[1:1] ;
assign n1115 =  ( n1113 ) ^ ( n1114 )  ;
assign n1116 =  ( n1115 ) ^ ( n90 )  ;
assign n1117 =  ( n1105 ) ? ( n1111 ) : ( n1116 ) ;
assign n1118 =  ( n1103 ) ? ( n1117 ) : ( bv_1_0_n74 ) ;
assign n1119 =  ( n1098 ) ? ( n1035 ) : ( n1118 ) ;
assign n1120 = ~ ( n1119 ) ;
assign n1121 =  ( n1093 ) | ( n1120 )  ;
assign n1122 = ki[1:1] ;
assign n1123 =  ( n1122 ) == ( bv_1_0_n74 )  ;
assign n1124 = i_wb_data[1:1] ;
assign n1125 = ~ ( n1124 ) ;
assign n1126 = sp[1:1] ;
assign n1127 =  ( n1125 ) ^ ( n1126 )  ;
assign n1128 = ~ ( n57 ) ;
assign n1129 =  ( n22 ) | ( n1128 )  ;
assign n1130 = ~ ( n1129 ) ;
assign n1131 =  ( n17 ) | ( n1130 )  ;
assign n1132 =  ( n1127 ) ^ ( n1131 )  ;
assign n1133 =  ( n1123 ) ? ( bv_1_0_n74 ) : ( n1132 ) ;
assign n1134 = ~ ( n1133 ) ;
assign n1135 =  ( n1121 ) | ( n1134 )  ;
assign n1136 =  ( n1036 ) ^ ( n1045 )  ;
assign n1137 = ~ ( n1136 ) ;
assign n1138 =  ( n1135 ) | ( n1137 )  ;
assign n1139 = ~ ( n1036 ) ;
assign n1140 = ~ ( n1045 ) ;
assign n1141 =  ( n1139 ) | ( n1140 )  ;
assign n1142 = ~ ( n1141 ) ;
assign n1143 =  ( n1142 ) ^ ( n941 )  ;
assign n1144 =  ( n1143 ) ^ ( n955 )  ;
assign n1145 = ~ ( n1144 ) ;
assign n1146 =  ( n1138 ) | ( n1145 )  ;
assign n1147 = ~ ( n1036 ) ;
assign n1148 = ~ ( n1045 ) ;
assign n1149 =  ( n1147 ) | ( n1148 )  ;
assign n1150 =  ( n941 ) ^ ( n955 )  ;
assign n1151 = ~ ( n1150 ) ;
assign n1152 =  ( n1149 ) | ( n1151 )  ;
assign n1153 = ~ ( n1152 ) ;
assign n1154 = ~ ( n941 ) ;
assign n1155 = ~ ( n955 ) ;
assign n1156 =  ( n1154 ) | ( n1155 )  ;
assign n1157 = ~ ( n1156 ) ;
assign n1158 =  ( n1153 ) ^ ( n1157 )  ;
assign n1159 =  ( n1158 ) ^ ( n813 )  ;
assign n1160 =  ( n1159 ) ^ ( n823 )  ;
assign n1161 = ~ ( n1160 ) ;
assign n1162 =  ( n1146 ) | ( n1161 )  ;
assign n1163 = ~ ( n1162 ) ;
assign n1164 =  ( n1075 ) | ( n1163 )  ;
assign n1165 = ~ ( n1092 ) ;
assign n1166 = ~ ( n1119 ) ;
assign n1167 = ~ ( n1133 ) ;
assign n1168 =  ( n1166 ) | ( n1167 )  ;
assign n1169 =  ( n1036 ) ^ ( n1045 )  ;
assign n1170 = ~ ( n1169 ) ;
assign n1171 =  ( n1168 ) | ( n1170 )  ;
assign n1172 = ~ ( n1144 ) ;
assign n1173 =  ( n1171 ) | ( n1172 )  ;
assign n1174 = ~ ( n1173 ) ;
assign n1175 =  ( n1174 ) ^ ( n1153 )  ;
assign n1176 = ~ ( n941 ) ;
assign n1177 = ~ ( n955 ) ;
assign n1178 =  ( n1176 ) | ( n1177 )  ;
assign n1179 = ~ ( n1178 ) ;
assign n1180 =  ( n1175 ) ^ ( n1179 )  ;
assign n1181 =  ( n1180 ) ^ ( n813 )  ;
assign n1182 =  ( n1181 ) ^ ( n823 )  ;
assign n1183 = ~ ( n1182 ) ;
assign n1184 =  ( n1165 ) | ( n1183 )  ;
assign n1185 = ~ ( n1119 ) ;
assign n1186 = ~ ( n1133 ) ;
assign n1187 =  ( n1185 ) | ( n1186 )  ;
assign n1188 =  ( n1036 ) ^ ( n1045 )  ;
assign n1189 = ~ ( n1188 ) ;
assign n1190 =  ( n1187 ) | ( n1189 )  ;
assign n1191 = ~ ( n1190 ) ;
assign n1192 = ~ ( n1036 ) ;
assign n1193 = ~ ( n1045 ) ;
assign n1194 =  ( n1192 ) | ( n1193 )  ;
assign n1195 = ~ ( n1194 ) ;
assign n1196 =  ( n1191 ) ^ ( n1195 )  ;
assign n1197 =  ( n1196 ) ^ ( n941 )  ;
assign n1198 =  ( n1197 ) ^ ( n955 )  ;
assign n1199 = ~ ( n1198 ) ;
assign n1200 =  ( n1184 ) | ( n1199 )  ;
assign n1201 = ki[0:0] ;
assign n1202 =  ( n1201 ) == ( bv_1_1_n2 )  ;
assign n1203 = ki[1:1] ;
assign n1204 =  ( n1203 ) == ( bv_1_0_n74 )  ;
assign n1205 =  ( n1202 ) | ( n1204 )  ;
assign n1206 = ki[1:1] ;
assign n1207 =  ( n1206 ) == ( bv_1_1_n2 )  ;
assign n1208 = ki[0:0] ;
assign n1209 =  ( n1208 ) == ( bv_1_1_n2 )  ;
assign n1210 =  ( n1207 ) | ( n1209 )  ;
assign n1211 = ki[1:1] ;
assign n1212 =  ( n1211 ) == ( bv_1_1_n2 )  ;
assign n1213 = i_wb_data[1:1] ;
assign n1214 = ~ ( n1213 ) ;
assign n1215 = sp[1:1] ;
assign n1216 =  ( n1214 ) ^ ( n1215 )  ;
assign n1217 =  ( n1216 ) ^ ( n1131 )  ;
assign n1218 = ~ ( n1217 ) ;
assign n1219 = i_wb_data[1:1] ;
assign n1220 = ~ ( n1219 ) ;
assign n1221 = sp[1:1] ;
assign n1222 =  ( n1220 ) ^ ( n1221 )  ;
assign n1223 =  ( n1222 ) ^ ( n1131 )  ;
assign n1224 =  ( n1212 ) ? ( n1218 ) : ( n1223 ) ;
assign n1225 =  ( n1210 ) ? ( n1224 ) : ( bv_1_0_n74 ) ;
assign n1226 =  ( n1205 ) ? ( n1118 ) : ( n1225 ) ;
assign n1227 = ~ ( n1226 ) ;
assign n1228 =  ( n1200 ) | ( n1227 )  ;
assign n1229 = ki[1:1] ;
assign n1230 =  ( n1229 ) == ( bv_1_0_n74 )  ;
assign n1231 = i_wb_data[1:1] ;
assign n1232 = ~ ( n1231 ) ;
assign n1233 = sp[1:1] ;
assign n1234 =  ( n1232 ) ^ ( n1233 )  ;
assign n1235 =  ( n1234 ) ^ ( n57 )  ;
assign n1236 =  ( n1230 ) ? ( bv_1_0_n74 ) : ( n1235 ) ;
assign n1237 = ~ ( n1236 ) ;
assign n1238 =  ( n1228 ) | ( n1237 )  ;
assign n1239 =  ( n1119 ) ^ ( n1133 )  ;
assign n1240 = ~ ( n1239 ) ;
assign n1241 =  ( n1238 ) | ( n1240 )  ;
assign n1242 = ~ ( n1119 ) ;
assign n1243 = ~ ( n1133 ) ;
assign n1244 =  ( n1242 ) | ( n1243 )  ;
assign n1245 = ~ ( n1244 ) ;
assign n1246 =  ( n1245 ) ^ ( n1036 )  ;
assign n1247 =  ( n1246 ) ^ ( n1045 )  ;
assign n1248 = ~ ( n1247 ) ;
assign n1249 =  ( n1241 ) | ( n1248 )  ;
assign n1250 = ~ ( n1249 ) ;
assign n1251 =  ( n1164 ) | ( n1250 )  ;
assign n1252 = ~ ( n1251 ) ;
assign n1253 =  ( n1010 ) | ( n1252 )  ;
assign n1254 = ~ ( n1253 ) ;
assign n1255 =  ( n986 ) | ( n1254 )  ;
assign n1256 = ~ ( n786 ) ;
assign n1257 = ~ ( n894 ) ;
assign n1258 =  ( n1256 ) | ( n1257 )  ;
assign n1259 = ~ ( n913 ) ;
assign n1260 =  ( n1258 ) | ( n1259 )  ;
assign n1261 = ~ ( n1008 ) ;
assign n1262 =  ( n1260 ) | ( n1261 )  ;
assign n1263 = ~ ( n1092 ) ;
assign n1264 =  ( n1262 ) | ( n1263 )  ;
assign n1265 = ~ ( n1182 ) ;
assign n1266 =  ( n1264 ) | ( n1265 )  ;
assign n1267 = ~ ( n1198 ) ;
assign n1268 =  ( n1266 ) | ( n1267 )  ;
assign n1269 = ~ ( n1226 ) ;
assign n1270 = ~ ( n1236 ) ;
assign n1271 =  ( n1269 ) | ( n1270 )  ;
assign n1272 =  ( n1119 ) ^ ( n1133 )  ;
assign n1273 = ~ ( n1272 ) ;
assign n1274 =  ( n1271 ) | ( n1273 )  ;
assign n1275 = ~ ( n1274 ) ;
assign n1276 = ~ ( n1119 ) ;
assign n1277 = ~ ( n1133 ) ;
assign n1278 =  ( n1276 ) | ( n1277 )  ;
assign n1279 = ~ ( n1278 ) ;
assign n1280 =  ( n1275 ) ^ ( n1279 )  ;
assign n1281 =  ( n1280 ) ^ ( n1036 )  ;
assign n1282 =  ( n1281 ) ^ ( n1045 )  ;
assign n1283 = ~ ( n1282 ) ;
assign n1284 =  ( n1268 ) | ( n1283 )  ;
assign n1285 = ki[0:0] ;
assign n1286 =  ( n1285 ) == ( bv_1_1_n2 )  ;
assign n1287 = ki[1:1] ;
assign n1288 =  ( n1287 ) == ( bv_1_0_n74 )  ;
assign n1289 =  ( n1286 ) | ( n1288 )  ;
assign n1290 = ki[1:1] ;
assign n1291 =  ( n1290 ) == ( bv_1_1_n2 )  ;
assign n1292 = ki[0:0] ;
assign n1293 =  ( n1292 ) == ( bv_1_1_n2 )  ;
assign n1294 =  ( n1291 ) | ( n1293 )  ;
assign n1295 = ki[1:1] ;
assign n1296 =  ( n1295 ) == ( bv_1_1_n2 )  ;
assign n1297 = i_wb_data[1:1] ;
assign n1298 = ~ ( n1297 ) ;
assign n1299 = sp[1:1] ;
assign n1300 =  ( n1298 ) ^ ( n1299 )  ;
assign n1301 =  ( n1300 ) ^ ( n57 )  ;
assign n1302 = ~ ( n1301 ) ;
assign n1303 = i_wb_data[1:1] ;
assign n1304 = ~ ( n1303 ) ;
assign n1305 = sp[1:1] ;
assign n1306 =  ( n1304 ) ^ ( n1305 )  ;
assign n1307 =  ( n1306 ) ^ ( n57 )  ;
assign n1308 =  ( n1296 ) ? ( n1302 ) : ( n1307 ) ;
assign n1309 =  ( n1294 ) ? ( n1308 ) : ( bv_1_0_n74 ) ;
assign n1310 =  ( n1289 ) ? ( n1225 ) : ( n1309 ) ;
assign n1311 = ~ ( n1310 ) ;
assign n1312 = ki[1:1] ;
assign n1313 =  ( n1312 ) == ( bv_1_0_n74 )  ;
assign n1314 = i_wb_data[1:1] ;
assign n1315 = ~ ( n1314 ) ;
assign n1316 = sp[1:1] ;
assign n1317 =  ( n1315 ) ^ ( n1316 )  ;
assign n1318 = ~ ( n53 ) ;
assign n1319 =  ( n22 ) | ( n1318 )  ;
assign n1320 = ~ ( n1319 ) ;
assign n1321 =  ( n17 ) | ( n1320 )  ;
assign n1322 =  ( n1317 ) ^ ( n1321 )  ;
assign n1323 =  ( n1313 ) ? ( bv_1_0_n74 ) : ( n1322 ) ;
assign n1324 = ~ ( n1323 ) ;
assign n1325 =  ( n1311 ) | ( n1324 )  ;
assign n1326 =  ( n1226 ) ^ ( n1236 )  ;
assign n1327 = ~ ( n1326 ) ;
assign n1328 =  ( n1325 ) | ( n1327 )  ;
assign n1329 = ~ ( n1226 ) ;
assign n1330 = ~ ( n1236 ) ;
assign n1331 =  ( n1329 ) | ( n1330 )  ;
assign n1332 = ~ ( n1331 ) ;
assign n1333 =  ( n1332 ) ^ ( n1119 )  ;
assign n1334 =  ( n1333 ) ^ ( n1133 )  ;
assign n1335 = ~ ( n1334 ) ;
assign n1336 =  ( n1328 ) | ( n1335 )  ;
assign n1337 = ~ ( n1336 ) ;
assign n1338 = ~ ( n1310 ) ;
assign n1339 = ~ ( n1323 ) ;
assign n1340 =  ( n1338 ) | ( n1339 )  ;
assign n1341 =  ( n1226 ) ^ ( n1236 )  ;
assign n1342 = ~ ( n1341 ) ;
assign n1343 =  ( n1340 ) | ( n1342 )  ;
assign n1344 = ~ ( n1343 ) ;
assign n1345 = ~ ( n1226 ) ;
assign n1346 = ~ ( n1236 ) ;
assign n1347 =  ( n1345 ) | ( n1346 )  ;
assign n1348 = ~ ( n1347 ) ;
assign n1349 =  ( n1344 ) ^ ( n1348 )  ;
assign n1350 =  ( n1349 ) ^ ( n1119 )  ;
assign n1351 =  ( n1350 ) ^ ( n1133 )  ;
assign n1352 = ~ ( n1351 ) ;
assign n1353 = ~ ( n1310 ) ;
assign n1354 = ~ ( n1323 ) ;
assign n1355 =  ( n1353 ) | ( n1354 )  ;
assign n1356 = ~ ( n1355 ) ;
assign n1357 =  ( n1356 ) ^ ( n1226 )  ;
assign n1358 =  ( n1357 ) ^ ( n1236 )  ;
assign n1359 = ~ ( n1358 ) ;
assign n1360 =  ( n1352 ) | ( n1359 )  ;
assign n1361 = ki[0:0] ;
assign n1362 =  ( n1361 ) == ( bv_1_1_n2 )  ;
assign n1363 = ki[1:1] ;
assign n1364 =  ( n1363 ) == ( bv_1_0_n74 )  ;
assign n1365 =  ( n1362 ) | ( n1364 )  ;
assign n1366 = ki[1:1] ;
assign n1367 =  ( n1366 ) == ( bv_1_1_n2 )  ;
assign n1368 = ki[0:0] ;
assign n1369 =  ( n1368 ) == ( bv_1_1_n2 )  ;
assign n1370 =  ( n1367 ) | ( n1369 )  ;
assign n1371 = ki[1:1] ;
assign n1372 =  ( n1371 ) == ( bv_1_1_n2 )  ;
assign n1373 = i_wb_data[1:1] ;
assign n1374 = ~ ( n1373 ) ;
assign n1375 = sp[1:1] ;
assign n1376 =  ( n1374 ) ^ ( n1375 )  ;
assign n1377 =  ( n1376 ) ^ ( n1321 )  ;
assign n1378 = ~ ( n1377 ) ;
assign n1379 = i_wb_data[1:1] ;
assign n1380 = ~ ( n1379 ) ;
assign n1381 = sp[1:1] ;
assign n1382 =  ( n1380 ) ^ ( n1381 )  ;
assign n1383 =  ( n1382 ) ^ ( n1321 )  ;
assign n1384 =  ( n1372 ) ? ( n1378 ) : ( n1383 ) ;
assign n1385 =  ( n1370 ) ? ( n1384 ) : ( bv_1_0_n74 ) ;
assign n1386 =  ( n1365 ) ? ( n1309 ) : ( n1385 ) ;
assign n1387 = ~ ( n1386 ) ;
assign n1388 = ki[1:1] ;
assign n1389 =  ( n1388 ) == ( bv_1_0_n74 )  ;
assign n1390 = i_wb_data[1:1] ;
assign n1391 = ~ ( n1390 ) ;
assign n1392 = sp[1:1] ;
assign n1393 =  ( n1391 ) ^ ( n1392 )  ;
assign n1394 =  ( n1393 ) ^ ( n53 )  ;
assign n1395 =  ( n1389 ) ? ( bv_1_0_n74 ) : ( n1394 ) ;
assign n1396 = ~ ( n1395 ) ;
assign n1397 =  ( n1387 ) | ( n1396 )  ;
assign n1398 =  ( n1310 ) ^ ( n1323 )  ;
assign n1399 = ~ ( n1398 ) ;
assign n1400 =  ( n1397 ) | ( n1399 )  ;
assign n1401 = ~ ( n1400 ) ;
assign n1402 = ~ ( n1386 ) ;
assign n1403 = ~ ( n1395 ) ;
assign n1404 =  ( n1402 ) | ( n1403 )  ;
assign n1405 = ~ ( n1404 ) ;
assign n1406 =  ( n1405 ) ^ ( n1310 )  ;
assign n1407 =  ( n1406 ) ^ ( n1323 )  ;
assign n1408 = ~ ( n1407 ) ;
assign n1409 = ki[0:0] ;
assign n1410 =  ( n1409 ) == ( bv_1_1_n2 )  ;
assign n1411 = ki[1:1] ;
assign n1412 =  ( n1411 ) == ( bv_1_0_n74 )  ;
assign n1413 =  ( n1410 ) | ( n1412 )  ;
assign n1414 = ki[1:1] ;
assign n1415 =  ( n1414 ) == ( bv_1_1_n2 )  ;
assign n1416 = ki[0:0] ;
assign n1417 =  ( n1416 ) == ( bv_1_1_n2 )  ;
assign n1418 =  ( n1415 ) | ( n1417 )  ;
assign n1419 = ki[1:1] ;
assign n1420 =  ( n1419 ) == ( bv_1_1_n2 )  ;
assign n1421 = i_wb_data[1:1] ;
assign n1422 = ~ ( n1421 ) ;
assign n1423 = sp[1:1] ;
assign n1424 =  ( n1422 ) ^ ( n1423 )  ;
assign n1425 =  ( n1424 ) ^ ( n53 )  ;
assign n1426 = ~ ( n1425 ) ;
assign n1427 = i_wb_data[1:1] ;
assign n1428 = ~ ( n1427 ) ;
assign n1429 = sp[1:1] ;
assign n1430 =  ( n1428 ) ^ ( n1429 )  ;
assign n1431 =  ( n1430 ) ^ ( n53 )  ;
assign n1432 =  ( n1420 ) ? ( n1426 ) : ( n1431 ) ;
assign n1433 =  ( n1418 ) ? ( n1432 ) : ( bv_1_0_n74 ) ;
assign n1434 =  ( n1413 ) ? ( n1385 ) : ( n1433 ) ;
assign n1435 = ~ ( n1434 ) ;
assign n1436 =  ( n1408 ) | ( n1435 )  ;
assign n1437 = ki[1:1] ;
assign n1438 =  ( n1437 ) == ( bv_1_0_n74 )  ;
assign n1439 = i_wb_data[0:0] ;
assign n1440 = ~ ( n1439 ) ;
assign n1441 =  ( bv_1_1_n2 ) ^ ( n1440 )  ;
assign n1442 = sp[0:0] ;
assign n1443 =  ( n1441 ) ^ ( n1442 )  ;
assign n1444 =  ( n1438 ) ? ( bv_1_0_n74 ) : ( n1443 ) ;
assign n1445 = ~ ( n1444 ) ;
assign n1446 =  ( n1436 ) | ( n1445 )  ;
assign n1447 =  ( n1386 ) ^ ( n1395 )  ;
assign n1448 = ~ ( n1447 ) ;
assign n1449 =  ( n1446 ) | ( n1448 )  ;
assign n1450 = ~ ( n1449 ) ;
assign n1451 =  ( n1401 ) | ( n1450 )  ;
assign n1452 = ~ ( n1451 ) ;
assign n1453 =  ( n1360 ) | ( n1452 )  ;
assign n1454 = ~ ( n1453 ) ;
assign n1455 =  ( n1337 ) | ( n1454 )  ;
assign n1456 = ~ ( n1351 ) ;
assign n1457 = ~ ( n1358 ) ;
assign n1458 =  ( n1456 ) | ( n1457 )  ;
assign n1459 = ~ ( n1407 ) ;
assign n1460 =  ( n1458 ) | ( n1459 )  ;
assign n1461 = ~ ( n1434 ) ;
assign n1462 = ~ ( n1444 ) ;
assign n1463 =  ( n1461 ) | ( n1462 )  ;
assign n1464 = ~ ( n1463 ) ;
assign n1465 =  ( n1464 ) ^ ( n1386 )  ;
assign n1466 =  ( n1465 ) ^ ( n1395 )  ;
assign n1467 = ~ ( n1466 ) ;
assign n1468 =  ( n1460 ) | ( n1467 )  ;
assign n1469 =  ( n1434 ) ^ ( n1444 )  ;
assign n1470 = ~ ( n1469 ) ;
assign n1471 =  ( n1468 ) | ( n1470 )  ;
assign n1472 = ki[0:0] ;
assign n1473 =  ( n1472 ) == ( bv_1_1_n2 )  ;
assign n1474 = ki[1:1] ;
assign n1475 =  ( n1474 ) == ( bv_1_0_n74 )  ;
assign n1476 =  ( n1473 ) | ( n1475 )  ;
assign n1477 = ki[1:1] ;
assign n1478 =  ( n1477 ) == ( bv_1_1_n2 )  ;
assign n1479 = ki[0:0] ;
assign n1480 =  ( n1479 ) == ( bv_1_1_n2 )  ;
assign n1481 =  ( n1478 ) | ( n1480 )  ;
assign n1482 = ki[1:1] ;
assign n1483 =  ( n1482 ) == ( bv_1_1_n2 )  ;
assign n1484 = i_wb_data[0:0] ;
assign n1485 = ~ ( n1484 ) ;
assign n1486 =  ( bv_1_1_n2 ) ^ ( n1485 )  ;
assign n1487 = sp[0:0] ;
assign n1488 =  ( n1486 ) ^ ( n1487 )  ;
assign n1489 = ~ ( n1488 ) ;
assign n1490 = i_wb_data[0:0] ;
assign n1491 = ~ ( n1490 ) ;
assign n1492 =  ( bv_1_1_n2 ) ^ ( n1491 )  ;
assign n1493 = sp[0:0] ;
assign n1494 =  ( n1492 ) ^ ( n1493 )  ;
assign n1495 =  ( n1483 ) ? ( n1489 ) : ( n1494 ) ;
assign n1496 =  ( n1481 ) ? ( n1495 ) : ( bv_1_0_n74 ) ;
assign n1497 =  ( n1476 ) ? ( n1433 ) : ( n1496 ) ;
assign n1498 = ~ ( n1497 ) ;
assign n1499 =  ( n1471 ) | ( n1498 )  ;
assign n1500 = ki[0:0] ;
assign n1501 =  ( n1500 ) == ( bv_1_1_n2 )  ;
assign n1502 = ki[1:1] ;
assign n1503 =  ( n1502 ) == ( bv_1_0_n74 )  ;
assign n1504 =  ( n1501 ) | ( n1503 )  ;
assign n1505 = ki[1:1] ;
assign n1506 =  ( n1504 ) ? ( n1496 ) : ( n1505 ) ;
assign n1507 = ~ ( n1506 ) ;
assign n1508 =  ( n1499 ) | ( n1507 )  ;
assign n1509 = ki[1:1] ;
assign n1510 = ~ ( n1509 ) ;
assign n1511 =  ( n1508 ) | ( n1510 )  ;
assign n1512 = ~ ( n1511 ) ;
assign n1513 =  ( n1455 ) | ( n1512 )  ;
assign n1514 = ~ ( n1513 ) ;
assign n1515 =  ( n1284 ) | ( n1514 )  ;
assign n1516 = ~ ( n1515 ) ;
assign n1517 =  ( n1255 ) | ( n1516 )  ;
assign n1518 = ~ ( n1517 ) ;
assign n1519 =  ( n678 ) | ( n1518 )  ;
assign n1520 = ~ ( n1519 ) ;
assign n1521 =  ( n641 ) | ( n1520 )  ;
assign n1522 = ~ ( n1521 ) ;
assign n1523 = kd[1:1] ;
assign n1524 =  ( n1523 ) == ( bv_1_1_n2 )  ;
assign n1525 = kd[0:0] ;
assign n1526 =  ( n1525 ) == ( bv_1_1_n2 )  ;
assign n1527 =  ( n1524 ) | ( n1526 )  ;
assign n1528 = kd[1:1] ;
assign n1529 =  ( n1528 ) == ( bv_1_1_n2 )  ;
assign n1530 =  ( n1529 ) ? ( bv_1_1_n2 ) : ( bv_1_0_n74 ) ;
assign n1531 =  ( n1527 ) ? ( n1530 ) : ( bv_1_0_n74 ) ;
assign n1532 = ~ ( n1531 ) ;
assign n1533 = ~ ( n1531 ) ;
assign n1534 = kd[0:0] ;
assign n1535 =  ( n1534 ) == ( bv_1_1_n2 )  ;
assign n1536 = kd[1:1] ;
assign n1537 =  ( n1536 ) == ( bv_1_0_n74 )  ;
assign n1538 =  ( n1535 ) | ( n1537 )  ;
assign n1539 = kd[1:1] ;
assign n1540 =  ( n1538 ) ? ( n1531 ) : ( n1539 ) ;
assign n1541 = ~ ( n1540 ) ;
assign n1542 =  ( n1533 ) | ( n1541 )  ;
assign n1543 = kd[1:1] ;
assign n1544 = ~ ( n1543 ) ;
assign n1545 =  ( n1542 ) | ( n1544 )  ;
assign n1546 = ~ ( n1545 ) ;
assign n1547 =  ( n1532 ) | ( n1546 )  ;
assign n1548 = ~ ( n1547 ) ;
assign n1549 =  ( n1522 ) ^ ( n1548 )  ;
assign n1550 = ~ ( n118 ) ;
assign n1551 =  ( n1550 ) | ( n110 )  ;
assign n1552 = ~ ( n1551 ) ;
assign n1553 = ~ ( n177 ) ;
assign n1554 =  ( n1552 ) | ( n1553 )  ;
assign n1555 = ~ ( n118 ) ;
assign n1556 =  ( n1555 ) | ( n110 )  ;
assign n1557 = ~ ( n1556 ) ;
assign n1558 =  ( n1557 ) | ( n200 )  ;
assign n1559 = ~ ( n292 ) ;
assign n1560 = ~ ( n416 ) ;
assign n1561 =  ( n1559 ) | ( n1560 )  ;
assign n1562 = ~ ( n1561 ) ;
assign n1563 =  ( n1558 ) | ( n1562 )  ;
assign n1564 = ~ ( n1563 ) ;
assign n1565 =  ( n1554 ) | ( n1564 )  ;
assign n1566 = ~ ( n118 ) ;
assign n1567 =  ( n1566 ) | ( n110 )  ;
assign n1568 = ~ ( n1567 ) ;
assign n1569 =  ( n1568 ) | ( n200 )  ;
assign n1570 = ~ ( n286 ) ;
assign n1571 =  ( n304 ) ^ ( n1570 )  ;
assign n1572 =  ( n1571 ) ^ ( n118 )  ;
assign n1573 = ~ ( n110 ) ;
assign n1574 =  ( n1572 ) ^ ( n1573 )  ;
assign n1575 = ~ ( n1574 ) ;
assign n1576 =  ( n1569 ) | ( n1575 )  ;
assign n1577 = ~ ( n434 ) ;
assign n1578 =  ( n1576 ) | ( n1577 )  ;
assign n1579 =  ( n524 ) | ( n632 )  ;
assign n1580 = ~ ( n546 ) ;
assign n1581 = ~ ( n676 ) ;
assign n1582 =  ( n1580 ) | ( n1581 )  ;
assign n1583 =  ( n766 ) | ( n872 )  ;
assign n1584 = ~ ( n1583 ) ;
assign n1585 =  ( n1582 ) | ( n1584 )  ;
assign n1586 = ~ ( n1585 ) ;
assign n1587 =  ( n1579 ) | ( n1586 )  ;
assign n1588 = ~ ( n1587 ) ;
assign n1589 =  ( n1578 ) | ( n1588 )  ;
assign n1590 = ~ ( n1589 ) ;
assign n1591 =  ( n1565 ) | ( n1590 )  ;
assign n1592 = ~ ( n118 ) ;
assign n1593 =  ( n1592 ) | ( n110 )  ;
assign n1594 = ~ ( n1593 ) ;
assign n1595 =  ( n1594 ) | ( n200 )  ;
assign n1596 = ~ ( n286 ) ;
assign n1597 =  ( n304 ) ^ ( n1596 )  ;
assign n1598 =  ( n1597 ) ^ ( n118 )  ;
assign n1599 = ~ ( n110 ) ;
assign n1600 =  ( n1598 ) ^ ( n1599 )  ;
assign n1601 = ~ ( n1600 ) ;
assign n1602 =  ( n1595 ) | ( n1601 )  ;
assign n1603 = ~ ( n434 ) ;
assign n1604 =  ( n1602 ) | ( n1603 )  ;
assign n1605 = ~ ( n546 ) ;
assign n1606 =  ( n1604 ) | ( n1605 )  ;
assign n1607 = ~ ( n676 ) ;
assign n1608 =  ( n1606 ) | ( n1607 )  ;
assign n1609 = ~ ( n786 ) ;
assign n1610 =  ( n1608 ) | ( n1609 )  ;
assign n1611 = ~ ( n894 ) ;
assign n1612 =  ( n1610 ) | ( n1611 )  ;
assign n1613 = ~ ( n913 ) ;
assign n1614 = ~ ( n941 ) ;
assign n1615 =  ( n1613 ) | ( n1614 )  ;
assign n1616 = ~ ( n955 ) ;
assign n1617 =  ( n1615 ) | ( n1616 )  ;
assign n1618 =  ( n813 ) ^ ( n823 )  ;
assign n1619 = ~ ( n1618 ) ;
assign n1620 =  ( n1617 ) | ( n1619 )  ;
assign n1621 = ~ ( n966 ) ;
assign n1622 =  ( n1620 ) | ( n1621 )  ;
assign n1623 = ~ ( n982 ) ;
assign n1624 =  ( n1622 ) | ( n1623 )  ;
assign n1625 = ~ ( n1624 ) ;
assign n1626 = ~ ( n913 ) ;
assign n1627 = ~ ( n1008 ) ;
assign n1628 =  ( n1626 ) | ( n1627 )  ;
assign n1629 =  ( n1075 ) | ( n1163 )  ;
assign n1630 = ~ ( n1629 ) ;
assign n1631 =  ( n1628 ) | ( n1630 )  ;
assign n1632 = ~ ( n1631 ) ;
assign n1633 =  ( n1625 ) | ( n1632 )  ;
assign n1634 = ~ ( n913 ) ;
assign n1635 = ~ ( n1008 ) ;
assign n1636 =  ( n1634 ) | ( n1635 )  ;
assign n1637 = ~ ( n1092 ) ;
assign n1638 =  ( n1636 ) | ( n1637 )  ;
assign n1639 = ~ ( n1182 ) ;
assign n1640 =  ( n1638 ) | ( n1639 )  ;
assign n1641 = ~ ( n1198 ) ;
assign n1642 = ~ ( n1226 ) ;
assign n1643 =  ( n1641 ) | ( n1642 )  ;
assign n1644 = ~ ( n1236 ) ;
assign n1645 =  ( n1643 ) | ( n1644 )  ;
assign n1646 =  ( n1119 ) ^ ( n1133 )  ;
assign n1647 = ~ ( n1646 ) ;
assign n1648 =  ( n1645 ) | ( n1647 )  ;
assign n1649 = ~ ( n1247 ) ;
assign n1650 =  ( n1648 ) | ( n1649 )  ;
assign n1651 = ~ ( n1650 ) ;
assign n1652 = ~ ( n1198 ) ;
assign n1653 = ~ ( n1282 ) ;
assign n1654 =  ( n1652 ) | ( n1653 )  ;
assign n1655 = ~ ( n1310 ) ;
assign n1656 =  ( n1654 ) | ( n1655 )  ;
assign n1657 = ~ ( n1323 ) ;
assign n1658 =  ( n1656 ) | ( n1657 )  ;
assign n1659 =  ( n1226 ) ^ ( n1236 )  ;
assign n1660 = ~ ( n1659 ) ;
assign n1661 =  ( n1658 ) | ( n1660 )  ;
assign n1662 = ~ ( n1334 ) ;
assign n1663 =  ( n1661 ) | ( n1662 )  ;
assign n1664 = ~ ( n1663 ) ;
assign n1665 =  ( n1651 ) | ( n1664 )  ;
assign n1666 = ~ ( n1665 ) ;
assign n1667 =  ( n1640 ) | ( n1666 )  ;
assign n1668 = ~ ( n1667 ) ;
assign n1669 =  ( n1633 ) | ( n1668 )  ;
assign n1670 = ~ ( n913 ) ;
assign n1671 = ~ ( n1008 ) ;
assign n1672 =  ( n1670 ) | ( n1671 )  ;
assign n1673 = ~ ( n1092 ) ;
assign n1674 =  ( n1672 ) | ( n1673 )  ;
assign n1675 = ~ ( n1182 ) ;
assign n1676 =  ( n1674 ) | ( n1675 )  ;
assign n1677 = ~ ( n1198 ) ;
assign n1678 =  ( n1676 ) | ( n1677 )  ;
assign n1679 = ~ ( n1282 ) ;
assign n1680 =  ( n1678 ) | ( n1679 )  ;
assign n1681 = ~ ( n1351 ) ;
assign n1682 =  ( n1680 ) | ( n1681 )  ;
assign n1683 = ~ ( n1358 ) ;
assign n1684 =  ( n1682 ) | ( n1683 )  ;
assign n1685 =  ( n1401 ) | ( n1450 )  ;
assign n1686 = ~ ( n1407 ) ;
assign n1687 = ~ ( n1466 ) ;
assign n1688 =  ( n1686 ) | ( n1687 )  ;
assign n1689 =  ( n1434 ) ^ ( n1444 )  ;
assign n1690 = ~ ( n1689 ) ;
assign n1691 =  ( n1688 ) | ( n1690 )  ;
assign n1692 = ~ ( n1497 ) ;
assign n1693 =  ( n1691 ) | ( n1692 )  ;
assign n1694 = ~ ( n1506 ) ;
assign n1695 =  ( n1693 ) | ( n1694 )  ;
assign n1696 = ki[1:1] ;
assign n1697 = ~ ( n1696 ) ;
assign n1698 =  ( n1695 ) | ( n1697 )  ;
assign n1699 = ~ ( n1698 ) ;
assign n1700 =  ( n1685 ) | ( n1699 )  ;
assign n1701 = ~ ( n1700 ) ;
assign n1702 =  ( n1684 ) | ( n1701 )  ;
assign n1703 = ~ ( n1702 ) ;
assign n1704 =  ( n1669 ) | ( n1703 )  ;
assign n1705 = ~ ( n1704 ) ;
assign n1706 =  ( n1612 ) | ( n1705 )  ;
assign n1707 = ~ ( n1706 ) ;
assign n1708 =  ( n1591 ) | ( n1707 )  ;
assign n1709 = ~ ( n1531 ) ;
assign n1710 =  ( n1708 ) | ( n1709 )  ;
assign n1711 =  ( n1710 ) | ( n1546 )  ;
assign n1712 = ~ ( n1711 ) ;
assign n1713 = ~ ( n118 ) ;
assign n1714 =  ( n1713 ) | ( n110 )  ;
assign n1715 = ~ ( n1714 ) ;
assign n1716 = ~ ( n177 ) ;
assign n1717 =  ( n1715 ) | ( n1716 )  ;
assign n1718 = ~ ( n1563 ) ;
assign n1719 =  ( n1717 ) | ( n1718 )  ;
assign n1720 = ~ ( n1589 ) ;
assign n1721 =  ( n1719 ) | ( n1720 )  ;
assign n1722 = ~ ( n1706 ) ;
assign n1723 =  ( n1721 ) | ( n1722 )  ;
assign n1724 = ~ ( n1723 ) ;
assign n1725 = ~ ( n1531 ) ;
assign n1726 =  ( n1725 ) | ( n1546 )  ;
assign n1727 = ~ ( n1726 ) ;
assign n1728 =  ( n1724 ) ^ ( n1727 )  ;
assign n1729 = ~ ( n1728 ) ;
assign n1730 = ~ ( n118 ) ;
assign n1731 =  ( n1730 ) | ( n110 )  ;
assign n1732 = ~ ( n1731 ) ;
assign n1733 =  ( n1729 ) | ( n1732 )  ;
assign n1734 = ~ ( n177 ) ;
assign n1735 =  ( n1733 ) | ( n1734 )  ;
assign n1736 = ~ ( n1563 ) ;
assign n1737 =  ( n1735 ) | ( n1736 )  ;
assign n1738 = ~ ( n1589 ) ;
assign n1739 =  ( n1737 ) | ( n1738 )  ;
assign n1740 = ~ ( n1706 ) ;
assign n1741 =  ( n1739 ) | ( n1740 )  ;
assign n1742 = ~ ( n1531 ) ;
assign n1743 =  ( n1741 ) | ( n1742 )  ;
assign n1744 =  ( n1743 ) | ( n1546 )  ;
assign n1745 = ~ ( n1744 ) ;
assign n1746 =  ( n1712 ) | ( n1745 )  ;
assign n1747 = ~ ( n1728 ) ;
assign n1748 = ~ ( n118 ) ;
assign n1749 =  ( n1748 ) | ( n110 )  ;
assign n1750 = ~ ( n1749 ) ;
assign n1751 = ~ ( n177 ) ;
assign n1752 =  ( n1750 ) | ( n1751 )  ;
assign n1753 = ~ ( n118 ) ;
assign n1754 =  ( n1753 ) | ( n110 )  ;
assign n1755 = ~ ( n1754 ) ;
assign n1756 =  ( n1755 ) | ( n200 )  ;
assign n1757 = ~ ( n292 ) ;
assign n1758 = ~ ( n416 ) ;
assign n1759 =  ( n1757 ) | ( n1758 )  ;
assign n1760 = ~ ( n635 ) ;
assign n1761 =  ( n1759 ) | ( n1760 )  ;
assign n1762 = ~ ( n286 ) ;
assign n1763 =  ( n304 ) ^ ( n1762 )  ;
assign n1764 =  ( n1763 ) ^ ( n118 )  ;
assign n1765 = ~ ( n110 ) ;
assign n1766 =  ( n1764 ) ^ ( n1765 )  ;
assign n1767 = ~ ( n1766 ) ;
assign n1768 = ~ ( n434 ) ;
assign n1769 =  ( n1767 ) | ( n1768 )  ;
assign n1770 = ~ ( n546 ) ;
assign n1771 =  ( n1769 ) | ( n1770 )  ;
assign n1772 = ~ ( n676 ) ;
assign n1773 =  ( n1771 ) | ( n1772 )  ;
assign n1774 =  ( n766 ) | ( n872 )  ;
assign n1775 =  ( n1774 ) | ( n985 )  ;
assign n1776 = ~ ( n1775 ) ;
assign n1777 =  ( n1773 ) | ( n1776 )  ;
assign n1778 = ~ ( n1777 ) ;
assign n1779 =  ( n1761 ) | ( n1778 )  ;
assign n1780 = ~ ( n1779 ) ;
assign n1781 =  ( n1756 ) | ( n1780 )  ;
assign n1782 = ~ ( n1781 ) ;
assign n1783 =  ( n1752 ) | ( n1782 )  ;
assign n1784 = ~ ( n118 ) ;
assign n1785 =  ( n1784 ) | ( n110 )  ;
assign n1786 = ~ ( n1785 ) ;
assign n1787 =  ( n1786 ) | ( n200 )  ;
assign n1788 = ~ ( n286 ) ;
assign n1789 =  ( n304 ) ^ ( n1788 )  ;
assign n1790 =  ( n1789 ) ^ ( n118 )  ;
assign n1791 = ~ ( n110 ) ;
assign n1792 =  ( n1790 ) ^ ( n1791 )  ;
assign n1793 = ~ ( n1792 ) ;
assign n1794 =  ( n1787 ) | ( n1793 )  ;
assign n1795 = ~ ( n434 ) ;
assign n1796 =  ( n1794 ) | ( n1795 )  ;
assign n1797 = ~ ( n546 ) ;
assign n1798 =  ( n1796 ) | ( n1797 )  ;
assign n1799 = ~ ( n676 ) ;
assign n1800 =  ( n1798 ) | ( n1799 )  ;
assign n1801 = ~ ( n786 ) ;
assign n1802 =  ( n1800 ) | ( n1801 )  ;
assign n1803 = ~ ( n894 ) ;
assign n1804 =  ( n1802 ) | ( n1803 )  ;
assign n1805 = ~ ( n913 ) ;
assign n1806 =  ( n1804 ) | ( n1805 )  ;
assign n1807 = ~ ( n1008 ) ;
assign n1808 =  ( n1806 ) | ( n1807 )  ;
assign n1809 =  ( n1075 ) | ( n1163 )  ;
assign n1810 =  ( n1809 ) | ( n1250 )  ;
assign n1811 = ~ ( n1092 ) ;
assign n1812 = ~ ( n1182 ) ;
assign n1813 =  ( n1811 ) | ( n1812 )  ;
assign n1814 = ~ ( n1198 ) ;
assign n1815 =  ( n1813 ) | ( n1814 )  ;
assign n1816 = ~ ( n1282 ) ;
assign n1817 =  ( n1815 ) | ( n1816 )  ;
assign n1818 =  ( n1337 ) | ( n1454 )  ;
assign n1819 = ~ ( n1818 ) ;
assign n1820 =  ( n1817 ) | ( n1819 )  ;
assign n1821 = ~ ( n1820 ) ;
assign n1822 =  ( n1810 ) | ( n1821 )  ;
assign n1823 = ~ ( n1092 ) ;
assign n1824 = ~ ( n1182 ) ;
assign n1825 =  ( n1823 ) | ( n1824 )  ;
assign n1826 = ~ ( n1198 ) ;
assign n1827 =  ( n1825 ) | ( n1826 )  ;
assign n1828 = ~ ( n1282 ) ;
assign n1829 =  ( n1827 ) | ( n1828 )  ;
assign n1830 = ~ ( n1351 ) ;
assign n1831 =  ( n1829 ) | ( n1830 )  ;
assign n1832 = ~ ( n1358 ) ;
assign n1833 =  ( n1831 ) | ( n1832 )  ;
assign n1834 = ~ ( n1407 ) ;
assign n1835 =  ( n1833 ) | ( n1834 )  ;
assign n1836 = ~ ( n1466 ) ;
assign n1837 =  ( n1835 ) | ( n1836 )  ;
assign n1838 =  ( n1434 ) ^ ( n1444 )  ;
assign n1839 = ~ ( n1838 ) ;
assign n1840 =  ( n1837 ) | ( n1839 )  ;
assign n1841 = ~ ( n1497 ) ;
assign n1842 =  ( n1840 ) | ( n1841 )  ;
assign n1843 = ~ ( n1506 ) ;
assign n1844 =  ( n1842 ) | ( n1843 )  ;
assign n1845 = ki[1:1] ;
assign n1846 = ~ ( n1845 ) ;
assign n1847 =  ( n1844 ) | ( n1846 )  ;
assign n1848 = ~ ( n1847 ) ;
assign n1849 =  ( n1822 ) | ( n1848 )  ;
assign n1850 = ~ ( n1849 ) ;
assign n1851 =  ( n1808 ) | ( n1850 )  ;
assign n1852 = ~ ( n1851 ) ;
assign n1853 =  ( n1783 ) | ( n1852 )  ;
assign n1854 = ~ ( n1531 ) ;
assign n1855 =  ( n1853 ) | ( n1854 )  ;
assign n1856 =  ( n1855 ) | ( n1546 )  ;
assign n1857 = ~ ( n1856 ) ;
assign n1858 = ~ ( n118 ) ;
assign n1859 =  ( n1858 ) | ( n110 )  ;
assign n1860 = ~ ( n1859 ) ;
assign n1861 = ~ ( n177 ) ;
assign n1862 =  ( n1860 ) | ( n1861 )  ;
assign n1863 = ~ ( n1781 ) ;
assign n1864 =  ( n1862 ) | ( n1863 )  ;
assign n1865 = ~ ( n1851 ) ;
assign n1866 =  ( n1864 ) | ( n1865 )  ;
assign n1867 = ~ ( n1866 ) ;
assign n1868 = ~ ( n1531 ) ;
assign n1869 =  ( n1868 ) | ( n1546 )  ;
assign n1870 = ~ ( n1869 ) ;
assign n1871 =  ( n1867 ) ^ ( n1870 )  ;
assign n1872 = ~ ( n1871 ) ;
assign n1873 = ~ ( n118 ) ;
assign n1874 =  ( n1873 ) | ( n110 )  ;
assign n1875 = ~ ( n1874 ) ;
assign n1876 =  ( n1872 ) | ( n1875 )  ;
assign n1877 = ~ ( n177 ) ;
assign n1878 =  ( n1876 ) | ( n1877 )  ;
assign n1879 = ~ ( n1781 ) ;
assign n1880 =  ( n1878 ) | ( n1879 )  ;
assign n1881 = ~ ( n1851 ) ;
assign n1882 =  ( n1880 ) | ( n1881 )  ;
assign n1883 = ~ ( n1531 ) ;
assign n1884 =  ( n1882 ) | ( n1883 )  ;
assign n1885 =  ( n1884 ) | ( n1546 )  ;
assign n1886 = ~ ( n1885 ) ;
assign n1887 =  ( n1857 ) | ( n1886 )  ;
assign n1888 = ~ ( n1887 ) ;
assign n1889 =  ( n1747 ) | ( n1888 )  ;
assign n1890 = ~ ( n1889 ) ;
assign n1891 =  ( n1746 ) | ( n1890 )  ;
assign n1892 = ~ ( n1728 ) ;
assign n1893 = ~ ( n1871 ) ;
assign n1894 =  ( n1892 ) | ( n1893 )  ;
assign n1895 = ~ ( n118 ) ;
assign n1896 =  ( n1895 ) | ( n110 )  ;
assign n1897 = ~ ( n1896 ) ;
assign n1898 = ~ ( n177 ) ;
assign n1899 =  ( n1897 ) | ( n1898 )  ;
assign n1900 = ~ ( n1563 ) ;
assign n1901 =  ( n1899 ) | ( n1900 )  ;
assign n1902 = ~ ( n118 ) ;
assign n1903 =  ( n1902 ) | ( n110 )  ;
assign n1904 = ~ ( n1903 ) ;
assign n1905 =  ( n1904 ) | ( n200 )  ;
assign n1906 = ~ ( n286 ) ;
assign n1907 =  ( n304 ) ^ ( n1906 )  ;
assign n1908 =  ( n1907 ) ^ ( n118 )  ;
assign n1909 = ~ ( n110 ) ;
assign n1910 =  ( n1908 ) ^ ( n1909 )  ;
assign n1911 = ~ ( n1910 ) ;
assign n1912 =  ( n1905 ) | ( n1911 )  ;
assign n1913 = ~ ( n434 ) ;
assign n1914 =  ( n1912 ) | ( n1913 )  ;
assign n1915 =  ( n524 ) | ( n632 )  ;
assign n1916 =  ( n1915 ) | ( n1586 )  ;
assign n1917 = ~ ( n546 ) ;
assign n1918 = ~ ( n676 ) ;
assign n1919 =  ( n1917 ) | ( n1918 )  ;
assign n1920 = ~ ( n786 ) ;
assign n1921 =  ( n1919 ) | ( n1920 )  ;
assign n1922 = ~ ( n894 ) ;
assign n1923 =  ( n1921 ) | ( n1922 )  ;
assign n1924 =  ( n1625 ) | ( n1632 )  ;
assign n1925 = ~ ( n1924 ) ;
assign n1926 =  ( n1923 ) | ( n1925 )  ;
assign n1927 = ~ ( n1926 ) ;
assign n1928 =  ( n1916 ) | ( n1927 )  ;
assign n1929 = ~ ( n1928 ) ;
assign n1930 =  ( n1914 ) | ( n1929 )  ;
assign n1931 = ~ ( n1930 ) ;
assign n1932 =  ( n1901 ) | ( n1931 )  ;
assign n1933 = ~ ( n118 ) ;
assign n1934 =  ( n1933 ) | ( n110 )  ;
assign n1935 = ~ ( n1934 ) ;
assign n1936 =  ( n1935 ) | ( n200 )  ;
assign n1937 = ~ ( n286 ) ;
assign n1938 =  ( n304 ) ^ ( n1937 )  ;
assign n1939 =  ( n1938 ) ^ ( n118 )  ;
assign n1940 = ~ ( n110 ) ;
assign n1941 =  ( n1939 ) ^ ( n1940 )  ;
assign n1942 = ~ ( n1941 ) ;
assign n1943 =  ( n1936 ) | ( n1942 )  ;
assign n1944 = ~ ( n434 ) ;
assign n1945 =  ( n1943 ) | ( n1944 )  ;
assign n1946 = ~ ( n546 ) ;
assign n1947 =  ( n1945 ) | ( n1946 )  ;
assign n1948 = ~ ( n676 ) ;
assign n1949 =  ( n1947 ) | ( n1948 )  ;
assign n1950 = ~ ( n786 ) ;
assign n1951 =  ( n1949 ) | ( n1950 )  ;
assign n1952 = ~ ( n894 ) ;
assign n1953 =  ( n1951 ) | ( n1952 )  ;
assign n1954 = ~ ( n913 ) ;
assign n1955 =  ( n1953 ) | ( n1954 )  ;
assign n1956 = ~ ( n1008 ) ;
assign n1957 =  ( n1955 ) | ( n1956 )  ;
assign n1958 = ~ ( n1092 ) ;
assign n1959 =  ( n1957 ) | ( n1958 )  ;
assign n1960 = ~ ( n1182 ) ;
assign n1961 =  ( n1959 ) | ( n1960 )  ;
assign n1962 =  ( n1651 ) | ( n1664 )  ;
assign n1963 = ~ ( n1198 ) ;
assign n1964 = ~ ( n1282 ) ;
assign n1965 =  ( n1963 ) | ( n1964 )  ;
assign n1966 = ~ ( n1351 ) ;
assign n1967 =  ( n1965 ) | ( n1966 )  ;
assign n1968 = ~ ( n1358 ) ;
assign n1969 =  ( n1967 ) | ( n1968 )  ;
assign n1970 =  ( n1401 ) | ( n1450 )  ;
assign n1971 = ~ ( n1970 ) ;
assign n1972 =  ( n1969 ) | ( n1971 )  ;
assign n1973 = ~ ( n1972 ) ;
assign n1974 =  ( n1962 ) | ( n1973 )  ;
assign n1975 = ~ ( n1198 ) ;
assign n1976 = ~ ( n1282 ) ;
assign n1977 =  ( n1975 ) | ( n1976 )  ;
assign n1978 = ~ ( n1351 ) ;
assign n1979 =  ( n1977 ) | ( n1978 )  ;
assign n1980 = ~ ( n1358 ) ;
assign n1981 =  ( n1979 ) | ( n1980 )  ;
assign n1982 = ~ ( n1407 ) ;
assign n1983 =  ( n1981 ) | ( n1982 )  ;
assign n1984 = ~ ( n1466 ) ;
assign n1985 =  ( n1983 ) | ( n1984 )  ;
assign n1986 =  ( n1434 ) ^ ( n1444 )  ;
assign n1987 = ~ ( n1986 ) ;
assign n1988 =  ( n1985 ) | ( n1987 )  ;
assign n1989 = ~ ( n1497 ) ;
assign n1990 =  ( n1988 ) | ( n1989 )  ;
assign n1991 = ~ ( n1506 ) ;
assign n1992 =  ( n1990 ) | ( n1991 )  ;
assign n1993 = ki[1:1] ;
assign n1994 = ~ ( n1993 ) ;
assign n1995 =  ( n1992 ) | ( n1994 )  ;
assign n1996 = ~ ( n1995 ) ;
assign n1997 =  ( n1974 ) | ( n1996 )  ;
assign n1998 = ~ ( n1997 ) ;
assign n1999 =  ( n1961 ) | ( n1998 )  ;
assign n2000 = ~ ( n1999 ) ;
assign n2001 =  ( n1932 ) | ( n2000 )  ;
assign n2002 = ~ ( n1531 ) ;
assign n2003 =  ( n2001 ) | ( n2002 )  ;
assign n2004 =  ( n2003 ) | ( n1546 )  ;
assign n2005 = ~ ( n2004 ) ;
assign n2006 = ~ ( n118 ) ;
assign n2007 =  ( n2006 ) | ( n110 )  ;
assign n2008 = ~ ( n2007 ) ;
assign n2009 = ~ ( n177 ) ;
assign n2010 =  ( n2008 ) | ( n2009 )  ;
assign n2011 = ~ ( n1563 ) ;
assign n2012 =  ( n2010 ) | ( n2011 )  ;
assign n2013 = ~ ( n1930 ) ;
assign n2014 =  ( n2012 ) | ( n2013 )  ;
assign n2015 = ~ ( n1999 ) ;
assign n2016 =  ( n2014 ) | ( n2015 )  ;
assign n2017 = ~ ( n2016 ) ;
assign n2018 = ~ ( n1531 ) ;
assign n2019 =  ( n2018 ) | ( n1546 )  ;
assign n2020 = ~ ( n2019 ) ;
assign n2021 =  ( n2017 ) ^ ( n2020 )  ;
assign n2022 = ~ ( n2021 ) ;
assign n2023 = ~ ( n118 ) ;
assign n2024 =  ( n2023 ) | ( n110 )  ;
assign n2025 = ~ ( n2024 ) ;
assign n2026 =  ( n2022 ) | ( n2025 )  ;
assign n2027 = ~ ( n177 ) ;
assign n2028 =  ( n2026 ) | ( n2027 )  ;
assign n2029 = ~ ( n1563 ) ;
assign n2030 =  ( n2028 ) | ( n2029 )  ;
assign n2031 = ~ ( n1930 ) ;
assign n2032 =  ( n2030 ) | ( n2031 )  ;
assign n2033 = ~ ( n1999 ) ;
assign n2034 =  ( n2032 ) | ( n2033 )  ;
assign n2035 = ~ ( n1531 ) ;
assign n2036 =  ( n2034 ) | ( n2035 )  ;
assign n2037 =  ( n2036 ) | ( n1546 )  ;
assign n2038 = ~ ( n2037 ) ;
assign n2039 =  ( n2005 ) | ( n2038 )  ;
assign n2040 = ~ ( n2021 ) ;
assign n2041 = ~ ( n118 ) ;
assign n2042 =  ( n2041 ) | ( n110 )  ;
assign n2043 = ~ ( n2042 ) ;
assign n2044 = ~ ( n177 ) ;
assign n2045 =  ( n2043 ) | ( n2044 )  ;
assign n2046 = ~ ( n639 ) ;
assign n2047 =  ( n2045 ) | ( n2046 )  ;
assign n2048 = ~ ( n118 ) ;
assign n2049 =  ( n2048 ) | ( n110 )  ;
assign n2050 = ~ ( n2049 ) ;
assign n2051 =  ( n2050 ) | ( n200 )  ;
assign n2052 = ~ ( n286 ) ;
assign n2053 =  ( n304 ) ^ ( n2052 )  ;
assign n2054 =  ( n2053 ) ^ ( n118 )  ;
assign n2055 = ~ ( n110 ) ;
assign n2056 =  ( n2054 ) ^ ( n2055 )  ;
assign n2057 = ~ ( n2056 ) ;
assign n2058 =  ( n2051 ) | ( n2057 )  ;
assign n2059 = ~ ( n434 ) ;
assign n2060 =  ( n2058 ) | ( n2059 )  ;
assign n2061 = ~ ( n546 ) ;
assign n2062 =  ( n2060 ) | ( n2061 )  ;
assign n2063 = ~ ( n676 ) ;
assign n2064 =  ( n2062 ) | ( n2063 )  ;
assign n2065 =  ( n766 ) | ( n872 )  ;
assign n2066 =  ( n2065 ) | ( n985 )  ;
assign n2067 =  ( n2066 ) | ( n1254 )  ;
assign n2068 = ~ ( n2067 ) ;
assign n2069 =  ( n2064 ) | ( n2068 )  ;
assign n2070 = ~ ( n2069 ) ;
assign n2071 =  ( n2047 ) | ( n2070 )  ;
assign n2072 = ~ ( n118 ) ;
assign n2073 =  ( n2072 ) | ( n110 )  ;
assign n2074 = ~ ( n2073 ) ;
assign n2075 =  ( n2074 ) | ( n200 )  ;
assign n2076 = ~ ( n286 ) ;
assign n2077 =  ( n304 ) ^ ( n2076 )  ;
assign n2078 =  ( n2077 ) ^ ( n118 )  ;
assign n2079 = ~ ( n110 ) ;
assign n2080 =  ( n2078 ) ^ ( n2079 )  ;
assign n2081 = ~ ( n2080 ) ;
assign n2082 =  ( n2075 ) | ( n2081 )  ;
assign n2083 = ~ ( n434 ) ;
assign n2084 =  ( n2082 ) | ( n2083 )  ;
assign n2085 = ~ ( n546 ) ;
assign n2086 =  ( n2084 ) | ( n2085 )  ;
assign n2087 = ~ ( n676 ) ;
assign n2088 =  ( n2086 ) | ( n2087 )  ;
assign n2089 = ~ ( n786 ) ;
assign n2090 =  ( n2088 ) | ( n2089 )  ;
assign n2091 = ~ ( n894 ) ;
assign n2092 =  ( n2090 ) | ( n2091 )  ;
assign n2093 = ~ ( n913 ) ;
assign n2094 =  ( n2092 ) | ( n2093 )  ;
assign n2095 = ~ ( n1008 ) ;
assign n2096 =  ( n2094 ) | ( n2095 )  ;
assign n2097 = ~ ( n1092 ) ;
assign n2098 =  ( n2096 ) | ( n2097 )  ;
assign n2099 = ~ ( n1182 ) ;
assign n2100 =  ( n2098 ) | ( n2099 )  ;
assign n2101 = ~ ( n1198 ) ;
assign n2102 =  ( n2100 ) | ( n2101 )  ;
assign n2103 = ~ ( n1282 ) ;
assign n2104 =  ( n2102 ) | ( n2103 )  ;
assign n2105 =  ( n1337 ) | ( n1454 )  ;
assign n2106 =  ( n2105 ) | ( n1512 )  ;
assign n2107 = ~ ( n2106 ) ;
assign n2108 =  ( n2104 ) | ( n2107 )  ;
assign n2109 = ~ ( n2108 ) ;
assign n2110 =  ( n2071 ) | ( n2109 )  ;
assign n2111 = ~ ( n1531 ) ;
assign n2112 =  ( n2110 ) | ( n2111 )  ;
assign n2113 =  ( n2112 ) | ( n1546 )  ;
assign n2114 = ~ ( n2113 ) ;
assign n2115 = ~ ( n118 ) ;
assign n2116 =  ( n2115 ) | ( n110 )  ;
assign n2117 = ~ ( n2116 ) ;
assign n2118 = ~ ( n177 ) ;
assign n2119 =  ( n2117 ) | ( n2118 )  ;
assign n2120 = ~ ( n639 ) ;
assign n2121 =  ( n2119 ) | ( n2120 )  ;
assign n2122 = ~ ( n2069 ) ;
assign n2123 =  ( n2121 ) | ( n2122 )  ;
assign n2124 = ~ ( n2108 ) ;
assign n2125 =  ( n2123 ) | ( n2124 )  ;
assign n2126 = ~ ( n2125 ) ;
assign n2127 = ~ ( n1531 ) ;
assign n2128 =  ( n2127 ) | ( n1546 )  ;
assign n2129 = ~ ( n2128 ) ;
assign n2130 =  ( n2126 ) ^ ( n2129 )  ;
assign n2131 = ~ ( n2130 ) ;
assign n2132 = ~ ( n118 ) ;
assign n2133 =  ( n2132 ) | ( n110 )  ;
assign n2134 = ~ ( n2133 ) ;
assign n2135 =  ( n2131 ) | ( n2134 )  ;
assign n2136 = ~ ( n177 ) ;
assign n2137 =  ( n2135 ) | ( n2136 )  ;
assign n2138 = ~ ( n639 ) ;
assign n2139 =  ( n2137 ) | ( n2138 )  ;
assign n2140 = ~ ( n2069 ) ;
assign n2141 =  ( n2139 ) | ( n2140 )  ;
assign n2142 = ~ ( n2108 ) ;
assign n2143 =  ( n2141 ) | ( n2142 )  ;
assign n2144 = ~ ( n1531 ) ;
assign n2145 =  ( n2143 ) | ( n2144 )  ;
assign n2146 =  ( n2145 ) | ( n1546 )  ;
assign n2147 = ~ ( n2146 ) ;
assign n2148 =  ( n2114 ) | ( n2147 )  ;
assign n2149 = ~ ( n2148 ) ;
assign n2150 =  ( n2040 ) | ( n2149 )  ;
assign n2151 = ~ ( n2150 ) ;
assign n2152 =  ( n2039 ) | ( n2151 )  ;
assign n2153 = ~ ( n2152 ) ;
assign n2154 =  ( n1894 ) | ( n2153 )  ;
assign n2155 = ~ ( n2154 ) ;
assign n2156 =  ( n1891 ) | ( n2155 )  ;
assign n2157 = ~ ( n1728 ) ;
assign n2158 = ~ ( n1871 ) ;
assign n2159 =  ( n2157 ) | ( n2158 )  ;
assign n2160 = ~ ( n2021 ) ;
assign n2161 =  ( n2159 ) | ( n2160 )  ;
assign n2162 = ~ ( n2130 ) ;
assign n2163 =  ( n2161 ) | ( n2162 )  ;
assign n2164 = ~ ( n118 ) ;
assign n2165 =  ( n2164 ) | ( n110 )  ;
assign n2166 = ~ ( n2165 ) ;
assign n2167 = ~ ( n177 ) ;
assign n2168 =  ( n2166 ) | ( n2167 )  ;
assign n2169 = ~ ( n1563 ) ;
assign n2170 =  ( n2168 ) | ( n2169 )  ;
assign n2171 = ~ ( n1589 ) ;
assign n2172 =  ( n2170 ) | ( n2171 )  ;
assign n2173 = ~ ( n118 ) ;
assign n2174 =  ( n2173 ) | ( n110 )  ;
assign n2175 = ~ ( n2174 ) ;
assign n2176 =  ( n2175 ) | ( n200 )  ;
assign n2177 = ~ ( n286 ) ;
assign n2178 =  ( n304 ) ^ ( n2177 )  ;
assign n2179 =  ( n2178 ) ^ ( n118 )  ;
assign n2180 = ~ ( n110 ) ;
assign n2181 =  ( n2179 ) ^ ( n2180 )  ;
assign n2182 = ~ ( n2181 ) ;
assign n2183 =  ( n2176 ) | ( n2182 )  ;
assign n2184 = ~ ( n434 ) ;
assign n2185 =  ( n2183 ) | ( n2184 )  ;
assign n2186 = ~ ( n546 ) ;
assign n2187 =  ( n2185 ) | ( n2186 )  ;
assign n2188 = ~ ( n676 ) ;
assign n2189 =  ( n2187 ) | ( n2188 )  ;
assign n2190 = ~ ( n786 ) ;
assign n2191 =  ( n2189 ) | ( n2190 )  ;
assign n2192 = ~ ( n894 ) ;
assign n2193 =  ( n2191 ) | ( n2192 )  ;
assign n2194 =  ( n1625 ) | ( n1632 )  ;
assign n2195 =  ( n2194 ) | ( n1668 )  ;
assign n2196 = ~ ( n2195 ) ;
assign n2197 =  ( n2193 ) | ( n2196 )  ;
assign n2198 = ~ ( n2197 ) ;
assign n2199 =  ( n2172 ) | ( n2198 )  ;
assign n2200 = ~ ( n118 ) ;
assign n2201 =  ( n2200 ) | ( n110 )  ;
assign n2202 = ~ ( n2201 ) ;
assign n2203 =  ( n2202 ) | ( n200 )  ;
assign n2204 = ~ ( n286 ) ;
assign n2205 =  ( n304 ) ^ ( n2204 )  ;
assign n2206 =  ( n2205 ) ^ ( n118 )  ;
assign n2207 = ~ ( n110 ) ;
assign n2208 =  ( n2206 ) ^ ( n2207 )  ;
assign n2209 = ~ ( n2208 ) ;
assign n2210 =  ( n2203 ) | ( n2209 )  ;
assign n2211 = ~ ( n434 ) ;
assign n2212 =  ( n2210 ) | ( n2211 )  ;
assign n2213 = ~ ( n546 ) ;
assign n2214 =  ( n2212 ) | ( n2213 )  ;
assign n2215 = ~ ( n676 ) ;
assign n2216 =  ( n2214 ) | ( n2215 )  ;
assign n2217 = ~ ( n786 ) ;
assign n2218 =  ( n2216 ) | ( n2217 )  ;
assign n2219 = ~ ( n894 ) ;
assign n2220 =  ( n2218 ) | ( n2219 )  ;
assign n2221 = ~ ( n913 ) ;
assign n2222 =  ( n2220 ) | ( n2221 )  ;
assign n2223 = ~ ( n1008 ) ;
assign n2224 =  ( n2222 ) | ( n2223 )  ;
assign n2225 = ~ ( n1092 ) ;
assign n2226 =  ( n2224 ) | ( n2225 )  ;
assign n2227 = ~ ( n1182 ) ;
assign n2228 =  ( n2226 ) | ( n2227 )  ;
assign n2229 = ~ ( n1198 ) ;
assign n2230 =  ( n2228 ) | ( n2229 )  ;
assign n2231 = ~ ( n1282 ) ;
assign n2232 =  ( n2230 ) | ( n2231 )  ;
assign n2233 = ~ ( n1351 ) ;
assign n2234 =  ( n2232 ) | ( n2233 )  ;
assign n2235 = ~ ( n1358 ) ;
assign n2236 =  ( n2234 ) | ( n2235 )  ;
assign n2237 =  ( n1401 ) | ( n1450 )  ;
assign n2238 =  ( n2237 ) | ( n1699 )  ;
assign n2239 = ~ ( n2238 ) ;
assign n2240 =  ( n2236 ) | ( n2239 )  ;
assign n2241 = ~ ( n2240 ) ;
assign n2242 =  ( n2199 ) | ( n2241 )  ;
assign n2243 = ~ ( n1531 ) ;
assign n2244 =  ( n2242 ) | ( n2243 )  ;
assign n2245 =  ( n2244 ) | ( n1546 )  ;
assign n2246 = ~ ( n2245 ) ;
assign n2247 = ~ ( n118 ) ;
assign n2248 =  ( n2247 ) | ( n110 )  ;
assign n2249 = ~ ( n2248 ) ;
assign n2250 = ~ ( n177 ) ;
assign n2251 =  ( n2249 ) | ( n2250 )  ;
assign n2252 = ~ ( n1563 ) ;
assign n2253 =  ( n2251 ) | ( n2252 )  ;
assign n2254 = ~ ( n1589 ) ;
assign n2255 =  ( n2253 ) | ( n2254 )  ;
assign n2256 = ~ ( n2197 ) ;
assign n2257 =  ( n2255 ) | ( n2256 )  ;
assign n2258 = ~ ( n2240 ) ;
assign n2259 =  ( n2257 ) | ( n2258 )  ;
assign n2260 = ~ ( n2259 ) ;
assign n2261 = ~ ( n1531 ) ;
assign n2262 =  ( n2261 ) | ( n1546 )  ;
assign n2263 = ~ ( n2262 ) ;
assign n2264 =  ( n2260 ) ^ ( n2263 )  ;
assign n2265 = ~ ( n2264 ) ;
assign n2266 = ~ ( n118 ) ;
assign n2267 =  ( n2266 ) | ( n110 )  ;
assign n2268 = ~ ( n2267 ) ;
assign n2269 =  ( n2265 ) | ( n2268 )  ;
assign n2270 = ~ ( n177 ) ;
assign n2271 =  ( n2269 ) | ( n2270 )  ;
assign n2272 = ~ ( n1563 ) ;
assign n2273 =  ( n2271 ) | ( n2272 )  ;
assign n2274 = ~ ( n1589 ) ;
assign n2275 =  ( n2273 ) | ( n2274 )  ;
assign n2276 = ~ ( n2197 ) ;
assign n2277 =  ( n2275 ) | ( n2276 )  ;
assign n2278 = ~ ( n2240 ) ;
assign n2279 =  ( n2277 ) | ( n2278 )  ;
assign n2280 = ~ ( n1531 ) ;
assign n2281 =  ( n2279 ) | ( n2280 )  ;
assign n2282 =  ( n2281 ) | ( n1546 )  ;
assign n2283 = ~ ( n2282 ) ;
assign n2284 =  ( n2246 ) | ( n2283 )  ;
assign n2285 = ~ ( n2264 ) ;
assign n2286 = ~ ( n118 ) ;
assign n2287 =  ( n2286 ) | ( n110 )  ;
assign n2288 = ~ ( n150 ) ;
assign n2289 = ~ ( n160 ) ;
assign n2290 =  ( n2288 ) | ( n2289 )  ;
assign n2291 = ~ ( n75 ) ;
assign n2292 =  ( n2291 ) ^ ( n100 )  ;
assign n2293 = ~ ( n2292 ) ;
assign n2294 =  ( n2290 ) | ( n2293 )  ;
assign n2295 = ~ ( n171 ) ;
assign n2296 =  ( n2294 ) | ( n2295 )  ;
assign n2297 = ~ ( n110 ) ;
assign n2298 =  ( n118 ) ^ ( n2297 )  ;
assign n2299 = ~ ( n2298 ) ;
assign n2300 =  ( n2296 ) | ( n2299 )  ;
assign n2301 = ~ ( n118 ) ;
assign n2302 =  ( n2301 ) | ( n110 )  ;
assign n2303 = ~ ( n2302 ) ;
assign n2304 =  ( n2300 ) | ( n2303 )  ;
assign n2305 = ~ ( n2304 ) ;
assign n2306 = ~ ( n292 ) ;
assign n2307 = ~ ( n416 ) ;
assign n2308 =  ( n2306 ) | ( n2307 )  ;
assign n2309 = ~ ( n635 ) ;
assign n2310 =  ( n2308 ) | ( n2309 )  ;
assign n2311 = ~ ( n1777 ) ;
assign n2312 =  ( n2310 ) | ( n2311 )  ;
assign n2313 = ~ ( n286 ) ;
assign n2314 =  ( n304 ) ^ ( n2313 )  ;
assign n2315 =  ( n2314 ) ^ ( n118 )  ;
assign n2316 = ~ ( n110 ) ;
assign n2317 =  ( n2315 ) ^ ( n2316 )  ;
assign n2318 = ~ ( n2317 ) ;
assign n2319 = ~ ( n434 ) ;
assign n2320 =  ( n2318 ) | ( n2319 )  ;
assign n2321 = ~ ( n546 ) ;
assign n2322 =  ( n2320 ) | ( n2321 )  ;
assign n2323 = ~ ( n676 ) ;
assign n2324 =  ( n2322 ) | ( n2323 )  ;
assign n2325 = ~ ( n786 ) ;
assign n2326 =  ( n2324 ) | ( n2325 )  ;
assign n2327 = ~ ( n894 ) ;
assign n2328 =  ( n2326 ) | ( n2327 )  ;
assign n2329 = ~ ( n913 ) ;
assign n2330 =  ( n2328 ) | ( n2329 )  ;
assign n2331 = ~ ( n1008 ) ;
assign n2332 =  ( n2330 ) | ( n2331 )  ;
assign n2333 =  ( n1075 ) | ( n1163 )  ;
assign n2334 =  ( n2333 ) | ( n1250 )  ;
assign n2335 =  ( n2334 ) | ( n1821 )  ;
assign n2336 = ~ ( n2335 ) ;
assign n2337 =  ( n2332 ) | ( n2336 )  ;
assign n2338 = ~ ( n2337 ) ;
assign n2339 =  ( n2312 ) | ( n2338 )  ;
assign n2340 = ~ ( n286 ) ;
assign n2341 =  ( n304 ) ^ ( n2340 )  ;
assign n2342 =  ( n2341 ) ^ ( n118 )  ;
assign n2343 = ~ ( n110 ) ;
assign n2344 =  ( n2342 ) ^ ( n2343 )  ;
assign n2345 = ~ ( n2344 ) ;
assign n2346 = ~ ( n434 ) ;
assign n2347 =  ( n2345 ) | ( n2346 )  ;
assign n2348 = ~ ( n546 ) ;
assign n2349 =  ( n2347 ) | ( n2348 )  ;
assign n2350 = ~ ( n676 ) ;
assign n2351 =  ( n2349 ) | ( n2350 )  ;
assign n2352 = ~ ( n786 ) ;
assign n2353 =  ( n2351 ) | ( n2352 )  ;
assign n2354 = ~ ( n894 ) ;
assign n2355 =  ( n2353 ) | ( n2354 )  ;
assign n2356 = ~ ( n913 ) ;
assign n2357 =  ( n2355 ) | ( n2356 )  ;
assign n2358 = ~ ( n1008 ) ;
assign n2359 =  ( n2357 ) | ( n2358 )  ;
assign n2360 = ~ ( n1092 ) ;
assign n2361 =  ( n2359 ) | ( n2360 )  ;
assign n2362 = ~ ( n1182 ) ;
assign n2363 =  ( n2361 ) | ( n2362 )  ;
assign n2364 = ~ ( n1198 ) ;
assign n2365 =  ( n2363 ) | ( n2364 )  ;
assign n2366 = ~ ( n1282 ) ;
assign n2367 =  ( n2365 ) | ( n2366 )  ;
assign n2368 = ~ ( n1351 ) ;
assign n2369 =  ( n2367 ) | ( n2368 )  ;
assign n2370 = ~ ( n1358 ) ;
assign n2371 =  ( n2369 ) | ( n2370 )  ;
assign n2372 = ~ ( n1407 ) ;
assign n2373 =  ( n2371 ) | ( n2372 )  ;
assign n2374 = ~ ( n1466 ) ;
assign n2375 =  ( n2373 ) | ( n2374 )  ;
assign n2376 =  ( n1434 ) ^ ( n1444 )  ;
assign n2377 = ~ ( n2376 ) ;
assign n2378 =  ( n2375 ) | ( n2377 )  ;
assign n2379 = ~ ( n1497 ) ;
assign n2380 =  ( n2378 ) | ( n2379 )  ;
assign n2381 = ~ ( n1506 ) ;
assign n2382 =  ( n2380 ) | ( n2381 )  ;
assign n2383 = ki[1:1] ;
assign n2384 = ~ ( n2383 ) ;
assign n2385 =  ( n2382 ) | ( n2384 )  ;
assign n2386 = ~ ( n2385 ) ;
assign n2387 =  ( n2339 ) | ( n2386 )  ;
assign n2388 = ~ ( n2387 ) ;
assign n2389 =  ( n200 ) | ( n2388 )  ;
assign n2390 = ~ ( n2389 ) ;
assign n2391 =  ( n2305 ) | ( n2390 )  ;
assign n2392 =  ( n2287 ) ^ ( n2391 )  ;
assign n2393 = ~ ( n2392 ) ;
assign n2394 = ~ ( n1531 ) ;
assign n2395 =  ( n2393 ) | ( n2394 )  ;
assign n2396 =  ( n2395 ) | ( n1546 )  ;
assign n2397 = ~ ( n2396 ) ;
assign n2398 = ~ ( n118 ) ;
assign n2399 =  ( n2398 ) | ( n110 )  ;
assign n2400 =  ( n2399 ) ^ ( n2391 )  ;
assign n2401 = ~ ( n1531 ) ;
assign n2402 =  ( n2401 ) | ( n1546 )  ;
assign n2403 = ~ ( n2402 ) ;
assign n2404 =  ( n2400 ) ^ ( n2403 )  ;
assign n2405 = ~ ( n2404 ) ;
assign n2406 = ~ ( n195 ) ;
assign n2407 = ~ ( n118 ) ;
assign n2408 =  ( n2407 ) | ( n110 )  ;
assign n2409 =  ( n2406 ) ^ ( n2408 )  ;
assign n2410 =  ( n2409 ) ^ ( n2387 )  ;
assign n2411 = ~ ( n2410 ) ;
assign n2412 =  ( n2405 ) | ( n2411 )  ;
assign n2413 = ~ ( n1531 ) ;
assign n2414 =  ( n2412 ) | ( n2413 )  ;
assign n2415 =  ( n2414 ) | ( n1546 )  ;
assign n2416 = ~ ( n2415 ) ;
assign n2417 =  ( n2397 ) | ( n2416 )  ;
assign n2418 = ~ ( n2417 ) ;
assign n2419 =  ( n2285 ) | ( n2418 )  ;
assign n2420 = ~ ( n2419 ) ;
assign n2421 =  ( n2284 ) | ( n2420 )  ;
assign n2422 = ~ ( n2264 ) ;
assign n2423 = ~ ( n2404 ) ;
assign n2424 =  ( n2422 ) | ( n2423 )  ;
assign n2425 = ~ ( n195 ) ;
assign n2426 = ~ ( n118 ) ;
assign n2427 =  ( n2426 ) | ( n110 )  ;
assign n2428 =  ( n2425 ) ^ ( n2427 )  ;
assign n2429 =  ( n2428 ) ^ ( n2387 )  ;
assign n2430 = ~ ( n1531 ) ;
assign n2431 =  ( n2430 ) | ( n1546 )  ;
assign n2432 = ~ ( n2431 ) ;
assign n2433 =  ( n2429 ) ^ ( n2432 )  ;
assign n2434 = ~ ( n2433 ) ;
assign n2435 =  ( n2424 ) | ( n2434 )  ;
assign n2436 = ~ ( n286 ) ;
assign n2437 =  ( n304 ) ^ ( n2436 )  ;
assign n2438 =  ( n2437 ) ^ ( n118 )  ;
assign n2439 = ~ ( n110 ) ;
assign n2440 =  ( n2438 ) ^ ( n2439 )  ;
assign n2441 =  ( n376 ) | ( n394 )  ;
assign n2442 = ~ ( n2441 ) ;
assign n2443 = ~ ( n414 ) ;
assign n2444 =  ( n2442 ) | ( n2443 )  ;
assign n2445 = ~ ( n2444 ) ;
assign n2446 = ~ ( n434 ) ;
assign n2447 =  ( n524 ) | ( n632 )  ;
assign n2448 =  ( n2447 ) | ( n1586 )  ;
assign n2449 =  ( n2448 ) | ( n1927 )  ;
assign n2450 = ~ ( n546 ) ;
assign n2451 = ~ ( n676 ) ;
assign n2452 =  ( n2450 ) | ( n2451 )  ;
assign n2453 = ~ ( n786 ) ;
assign n2454 =  ( n2452 ) | ( n2453 )  ;
assign n2455 = ~ ( n894 ) ;
assign n2456 =  ( n2454 ) | ( n2455 )  ;
assign n2457 = ~ ( n913 ) ;
assign n2458 =  ( n2456 ) | ( n2457 )  ;
assign n2459 = ~ ( n1008 ) ;
assign n2460 =  ( n2458 ) | ( n2459 )  ;
assign n2461 = ~ ( n1092 ) ;
assign n2462 =  ( n2460 ) | ( n2461 )  ;
assign n2463 = ~ ( n1182 ) ;
assign n2464 =  ( n2462 ) | ( n2463 )  ;
assign n2465 =  ( n1651 ) | ( n1664 )  ;
assign n2466 =  ( n2465 ) | ( n1973 )  ;
assign n2467 = ~ ( n2466 ) ;
assign n2468 =  ( n2464 ) | ( n2467 )  ;
assign n2469 = ~ ( n2468 ) ;
assign n2470 =  ( n2449 ) | ( n2469 )  ;
assign n2471 = ~ ( n546 ) ;
assign n2472 = ~ ( n676 ) ;
assign n2473 =  ( n2471 ) | ( n2472 )  ;
assign n2474 = ~ ( n786 ) ;
assign n2475 =  ( n2473 ) | ( n2474 )  ;
assign n2476 = ~ ( n894 ) ;
assign n2477 =  ( n2475 ) | ( n2476 )  ;
assign n2478 = ~ ( n913 ) ;
assign n2479 =  ( n2477 ) | ( n2478 )  ;
assign n2480 = ~ ( n1008 ) ;
assign n2481 =  ( n2479 ) | ( n2480 )  ;
assign n2482 = ~ ( n1092 ) ;
assign n2483 =  ( n2481 ) | ( n2482 )  ;
assign n2484 = ~ ( n1182 ) ;
assign n2485 =  ( n2483 ) | ( n2484 )  ;
assign n2486 = ~ ( n1198 ) ;
assign n2487 =  ( n2485 ) | ( n2486 )  ;
assign n2488 = ~ ( n1282 ) ;
assign n2489 =  ( n2487 ) | ( n2488 )  ;
assign n2490 = ~ ( n1351 ) ;
assign n2491 =  ( n2489 ) | ( n2490 )  ;
assign n2492 = ~ ( n1358 ) ;
assign n2493 =  ( n2491 ) | ( n2492 )  ;
assign n2494 = ~ ( n1407 ) ;
assign n2495 =  ( n2493 ) | ( n2494 )  ;
assign n2496 = ~ ( n1466 ) ;
assign n2497 =  ( n2495 ) | ( n2496 )  ;
assign n2498 =  ( n1434 ) ^ ( n1444 )  ;
assign n2499 = ~ ( n2498 ) ;
assign n2500 =  ( n2497 ) | ( n2499 )  ;
assign n2501 = ~ ( n1497 ) ;
assign n2502 =  ( n2500 ) | ( n2501 )  ;
assign n2503 = ~ ( n1506 ) ;
assign n2504 =  ( n2502 ) | ( n2503 )  ;
assign n2505 = ki[1:1] ;
assign n2506 = ~ ( n2505 ) ;
assign n2507 =  ( n2504 ) | ( n2506 )  ;
assign n2508 = ~ ( n2507 ) ;
assign n2509 =  ( n2470 ) | ( n2508 )  ;
assign n2510 = ~ ( n2509 ) ;
assign n2511 =  ( n2446 ) | ( n2510 )  ;
assign n2512 = ~ ( n2511 ) ;
assign n2513 =  ( n2445 ) | ( n2512 )  ;
assign n2514 =  ( n2440 ) ^ ( n2513 )  ;
assign n2515 = ~ ( n2514 ) ;
assign n2516 = ~ ( n1531 ) ;
assign n2517 =  ( n2515 ) | ( n2516 )  ;
assign n2518 =  ( n2517 ) | ( n1546 )  ;
assign n2519 = ~ ( n2518 ) ;
assign n2520 = ~ ( n286 ) ;
assign n2521 =  ( n304 ) ^ ( n2520 )  ;
assign n2522 =  ( n2521 ) ^ ( n118 )  ;
assign n2523 = ~ ( n110 ) ;
assign n2524 =  ( n2522 ) ^ ( n2523 )  ;
assign n2525 =  ( n2445 ) | ( n2512 )  ;
assign n2526 =  ( n2524 ) ^ ( n2525 )  ;
assign n2527 = ~ ( n1531 ) ;
assign n2528 =  ( n2527 ) | ( n1546 )  ;
assign n2529 = ~ ( n2528 ) ;
assign n2530 =  ( n2526 ) ^ ( n2529 )  ;
assign n2531 = ~ ( n2530 ) ;
assign n2532 =  ( n376 ) | ( n394 )  ;
assign n2533 =  ( bv_1_1_n2 ) ^ ( n2532 )  ;
assign n2534 =  ( n2533 ) ^ ( n406 )  ;
assign n2535 = ~ ( n268 ) ;
assign n2536 =  ( n2534 ) ^ ( n2535 )  ;
assign n2537 = ~ ( n100 ) ;
assign n2538 =  ( n75 ) | ( n2537 )  ;
assign n2539 = ~ ( n2538 ) ;
assign n2540 =  ( n2536 ) ^ ( n2539 )  ;
assign n2541 =  ( n2540 ) ^ ( n110 )  ;
assign n2542 =  ( n524 ) | ( n632 )  ;
assign n2543 =  ( n2542 ) | ( n1586 )  ;
assign n2544 =  ( n2543 ) | ( n1927 )  ;
assign n2545 =  ( n2544 ) | ( n2469 )  ;
assign n2546 =  ( n2545 ) | ( n2508 )  ;
assign n2547 =  ( n2541 ) ^ ( n2546 )  ;
assign n2548 = ~ ( n2547 ) ;
assign n2549 =  ( n2531 ) | ( n2548 )  ;
assign n2550 =  ( n1531 ) ^ ( n1546 )  ;
assign n2551 = ~ ( n2550 ) ;
assign n2552 =  ( n2549 ) | ( n2551 )  ;
assign n2553 = ~ ( n2552 ) ;
assign n2554 =  ( n2519 ) | ( n2553 )  ;
assign n2555 = ~ ( n2530 ) ;
assign n2556 =  ( n376 ) | ( n394 )  ;
assign n2557 =  ( bv_1_1_n2 ) ^ ( n2556 )  ;
assign n2558 =  ( n2557 ) ^ ( n406 )  ;
assign n2559 = ~ ( n268 ) ;
assign n2560 =  ( n2558 ) ^ ( n2559 )  ;
assign n2561 = ~ ( n100 ) ;
assign n2562 =  ( n75 ) | ( n2561 )  ;
assign n2563 = ~ ( n2562 ) ;
assign n2564 =  ( n2560 ) ^ ( n2563 )  ;
assign n2565 =  ( n2564 ) ^ ( n110 )  ;
assign n2566 =  ( n524 ) | ( n632 )  ;
assign n2567 =  ( n2566 ) | ( n1586 )  ;
assign n2568 =  ( n2567 ) | ( n1927 )  ;
assign n2569 =  ( n2568 ) | ( n2469 )  ;
assign n2570 =  ( n2569 ) | ( n2508 )  ;
assign n2571 =  ( n2565 ) ^ ( n2570 )  ;
assign n2572 =  ( n2571 ) ^ ( n1531 )  ;
assign n2573 =  ( n2572 ) ^ ( n1546 )  ;
assign n2574 = ~ ( n2573 ) ;
assign n2575 =  ( n2555 ) | ( n2574 )  ;
assign n2576 =  ( bv_1_1_n2 ) ^ ( n535 )  ;
assign n2577 =  ( n2576 ) ^ ( n385 )  ;
assign n2578 =  ( n2577 ) ^ ( n365 )  ;
assign n2579 = ~ ( n150 ) ;
assign n2580 = ~ ( n160 ) ;
assign n2581 =  ( n2579 ) | ( n2580 )  ;
assign n2582 = ~ ( n2581 ) ;
assign n2583 =  ( n2578 ) ^ ( n2582 )  ;
assign n2584 = ~ ( n75 ) ;
assign n2585 =  ( n2583 ) ^ ( n2584 )  ;
assign n2586 =  ( n2585 ) ^ ( n100 )  ;
assign n2587 = ~ ( n573 ) ;
assign n2588 = ~ ( n583 ) ;
assign n2589 =  ( n2587 ) | ( n2588 )  ;
assign n2590 =  ( n462 ) ^ ( n482 )  ;
assign n2591 = ~ ( n2590 ) ;
assign n2592 =  ( n2589 ) | ( n2591 )  ;
assign n2593 = ~ ( n594 ) ;
assign n2594 =  ( n2592 ) | ( n2593 )  ;
assign n2595 = ~ ( n610 ) ;
assign n2596 =  ( n2594 ) | ( n2595 )  ;
assign n2597 = ~ ( n629 ) ;
assign n2598 =  ( n2596 ) | ( n2597 )  ;
assign n2599 = ~ ( n2598 ) ;
assign n2600 = ~ ( n676 ) ;
assign n2601 =  ( n766 ) | ( n872 )  ;
assign n2602 =  ( n2601 ) | ( n985 )  ;
assign n2603 =  ( n2602 ) | ( n1254 )  ;
assign n2604 =  ( n2603 ) | ( n1516 )  ;
assign n2605 = ~ ( n2604 ) ;
assign n2606 =  ( n2600 ) | ( n2605 )  ;
assign n2607 = ~ ( n2606 ) ;
assign n2608 =  ( n2599 ) | ( n2607 )  ;
assign n2609 =  ( n2586 ) ^ ( n2608 )  ;
assign n2610 = ~ ( n2609 ) ;
assign n2611 =  ( n1531 ) ^ ( n1546 )  ;
assign n2612 = ~ ( n2611 ) ;
assign n2613 =  ( n2610 ) | ( n2612 )  ;
assign n2614 = ~ ( n2613 ) ;
assign n2615 =  ( bv_1_1_n2 ) ^ ( n535 )  ;
assign n2616 =  ( n2615 ) ^ ( n385 )  ;
assign n2617 =  ( n2616 ) ^ ( n365 )  ;
assign n2618 = ~ ( n150 ) ;
assign n2619 = ~ ( n160 ) ;
assign n2620 =  ( n2618 ) | ( n2619 )  ;
assign n2621 = ~ ( n2620 ) ;
assign n2622 =  ( n2617 ) ^ ( n2621 )  ;
assign n2623 = ~ ( n75 ) ;
assign n2624 =  ( n2622 ) ^ ( n2623 )  ;
assign n2625 =  ( n2624 ) ^ ( n100 )  ;
assign n2626 =  ( n2599 ) | ( n2607 )  ;
assign n2627 =  ( n2625 ) ^ ( n2626 )  ;
assign n2628 =  ( n2627 ) ^ ( n1531 )  ;
assign n2629 =  ( n2628 ) ^ ( n1546 )  ;
assign n2630 = ~ ( n2629 ) ;
assign n2631 =  ( n667 ) ^ ( n621 )  ;
assign n2632 =  ( n2631 ) ^ ( n502 )  ;
assign n2633 = ~ ( n227 ) ;
assign n2634 = ~ ( n247 ) ;
assign n2635 =  ( n2633 ) | ( n2634 )  ;
assign n2636 = ~ ( n2635 ) ;
assign n2637 =  ( n2632 ) ^ ( n2636 )  ;
assign n2638 =  ( n2637 ) ^ ( n150 )  ;
assign n2639 =  ( n2638 ) ^ ( n160 )  ;
assign n2640 =  ( n766 ) | ( n872 )  ;
assign n2641 =  ( n2640 ) | ( n985 )  ;
assign n2642 =  ( n2641 ) | ( n1254 )  ;
assign n2643 =  ( n2642 ) | ( n1516 )  ;
assign n2644 =  ( n2639 ) ^ ( n2643 )  ;
assign n2645 = ~ ( n2644 ) ;
assign n2646 =  ( n2630 ) | ( n2645 )  ;
assign n2647 =  ( n1531 ) ^ ( n1546 )  ;
assign n2648 = ~ ( n2647 ) ;
assign n2649 =  ( n2646 ) | ( n2648 )  ;
assign n2650 = ~ ( n2649 ) ;
assign n2651 =  ( n2614 ) | ( n2650 )  ;
assign n2652 = ~ ( n2651 ) ;
assign n2653 =  ( n2575 ) | ( n2652 )  ;
assign n2654 = ~ ( n2653 ) ;
assign n2655 =  ( n2554 ) | ( n2654 )  ;
assign n2656 = ~ ( n2655 ) ;
assign n2657 =  ( n2435 ) | ( n2656 )  ;
assign n2658 = ~ ( n2657 ) ;
assign n2659 =  ( n2421 ) | ( n2658 )  ;
assign n2660 = ~ ( n2659 ) ;
assign n2661 =  ( n2163 ) | ( n2660 )  ;
assign n2662 = ~ ( n2661 ) ;
assign n2663 =  ( n2156 ) | ( n2662 )  ;
assign n2664 = ~ ( n1728 ) ;
assign n2665 = ~ ( n1871 ) ;
assign n2666 =  ( n2664 ) | ( n2665 )  ;
assign n2667 = ~ ( n2021 ) ;
assign n2668 =  ( n2666 ) | ( n2667 )  ;
assign n2669 = ~ ( n2130 ) ;
assign n2670 =  ( n2668 ) | ( n2669 )  ;
assign n2671 = ~ ( n2264 ) ;
assign n2672 =  ( n2670 ) | ( n2671 )  ;
assign n2673 = ~ ( n2404 ) ;
assign n2674 =  ( n2672 ) | ( n2673 )  ;
assign n2675 = ~ ( n2433 ) ;
assign n2676 =  ( n2674 ) | ( n2675 )  ;
assign n2677 = ~ ( n2530 ) ;
assign n2678 =  ( n2676 ) | ( n2677 )  ;
assign n2679 = ~ ( n2573 ) ;
assign n2680 =  ( n2678 ) | ( n2679 )  ;
assign n2681 = ~ ( n2629 ) ;
assign n2682 =  ( n2680 ) | ( n2681 )  ;
assign n2683 =  ( n667 ) ^ ( n621 )  ;
assign n2684 =  ( n2683 ) ^ ( n502 )  ;
assign n2685 = ~ ( n227 ) ;
assign n2686 = ~ ( n247 ) ;
assign n2687 =  ( n2685 ) | ( n2686 )  ;
assign n2688 = ~ ( n2687 ) ;
assign n2689 =  ( n2684 ) ^ ( n2688 )  ;
assign n2690 =  ( n2689 ) ^ ( n150 )  ;
assign n2691 =  ( n2690 ) ^ ( n160 )  ;
assign n2692 =  ( n766 ) | ( n872 )  ;
assign n2693 =  ( n2692 ) | ( n985 )  ;
assign n2694 =  ( n2693 ) | ( n1254 )  ;
assign n2695 =  ( n2694 ) | ( n1516 )  ;
assign n2696 =  ( n2691 ) ^ ( n2695 )  ;
assign n2697 =  ( n2696 ) ^ ( n1531 )  ;
assign n2698 =  ( n2697 ) ^ ( n1546 )  ;
assign n2699 = ~ ( n2698 ) ;
assign n2700 =  ( n2682 ) | ( n2699 )  ;
assign n2701 =  ( n777 ) ^ ( n755 )  ;
assign n2702 =  ( n2701 ) ^ ( n603 )  ;
assign n2703 = ~ ( n336 ) ;
assign n2704 = ~ ( n345 ) ;
assign n2705 =  ( n2703 ) | ( n2704 )  ;
assign n2706 = ~ ( n2705 ) ;
assign n2707 =  ( n2702 ) ^ ( n2706 )  ;
assign n2708 =  ( n2707 ) ^ ( n227 )  ;
assign n2709 =  ( n2708 ) ^ ( n247 )  ;
assign n2710 = ~ ( n813 ) ;
assign n2711 = ~ ( n823 ) ;
assign n2712 =  ( n2710 ) | ( n2711 )  ;
assign n2713 =  ( n704 ) ^ ( n717 )  ;
assign n2714 = ~ ( n2713 ) ;
assign n2715 =  ( n2712 ) | ( n2714 )  ;
assign n2716 = ~ ( n834 ) ;
assign n2717 =  ( n2715 ) | ( n2716 )  ;
assign n2718 = ~ ( n850 ) ;
assign n2719 =  ( n2717 ) | ( n2718 )  ;
assign n2720 = ~ ( n869 ) ;
assign n2721 =  ( n2719 ) | ( n2720 )  ;
assign n2722 = ~ ( n2721 ) ;
assign n2723 = ~ ( n894 ) ;
assign n2724 =  ( n1625 ) | ( n1632 )  ;
assign n2725 =  ( n2724 ) | ( n1668 )  ;
assign n2726 =  ( n2725 ) | ( n1703 )  ;
assign n2727 = ~ ( n2726 ) ;
assign n2728 =  ( n2723 ) | ( n2727 )  ;
assign n2729 = ~ ( n2728 ) ;
assign n2730 =  ( n2722 ) | ( n2729 )  ;
assign n2731 =  ( n2709 ) ^ ( n2730 )  ;
assign n2732 = ~ ( n2731 ) ;
assign n2733 =  ( n1531 ) ^ ( n1546 )  ;
assign n2734 = ~ ( n2733 ) ;
assign n2735 =  ( n2732 ) | ( n2734 )  ;
assign n2736 = ~ ( n2735 ) ;
assign n2737 =  ( n777 ) ^ ( n755 )  ;
assign n2738 =  ( n2737 ) ^ ( n603 )  ;
assign n2739 = ~ ( n336 ) ;
assign n2740 = ~ ( n345 ) ;
assign n2741 =  ( n2739 ) | ( n2740 )  ;
assign n2742 = ~ ( n2741 ) ;
assign n2743 =  ( n2738 ) ^ ( n2742 )  ;
assign n2744 =  ( n2743 ) ^ ( n227 )  ;
assign n2745 =  ( n2744 ) ^ ( n247 )  ;
assign n2746 =  ( n2722 ) | ( n2729 )  ;
assign n2747 =  ( n2745 ) ^ ( n2746 )  ;
assign n2748 =  ( n2747 ) ^ ( n1531 )  ;
assign n2749 =  ( n2748 ) ^ ( n1546 )  ;
assign n2750 = ~ ( n2749 ) ;
assign n2751 =  ( n885 ) ^ ( n861 )  ;
assign n2752 =  ( n2751 ) ^ ( n737 )  ;
assign n2753 = ~ ( n462 ) ;
assign n2754 = ~ ( n482 ) ;
assign n2755 =  ( n2753 ) | ( n2754 )  ;
assign n2756 = ~ ( n2755 ) ;
assign n2757 =  ( n2752 ) ^ ( n2756 )  ;
assign n2758 =  ( n2757 ) ^ ( n336 )  ;
assign n2759 =  ( n2758 ) ^ ( n345 )  ;
assign n2760 =  ( n1625 ) | ( n1632 )  ;
assign n2761 =  ( n2760 ) | ( n1668 )  ;
assign n2762 =  ( n2761 ) | ( n1703 )  ;
assign n2763 =  ( n2759 ) ^ ( n2762 )  ;
assign n2764 = ~ ( n2763 ) ;
assign n2765 =  ( n2750 ) | ( n2764 )  ;
assign n2766 =  ( n1531 ) ^ ( n1546 )  ;
assign n2767 = ~ ( n2766 ) ;
assign n2768 =  ( n2765 ) | ( n2767 )  ;
assign n2769 = ~ ( n2768 ) ;
assign n2770 =  ( n2736 ) | ( n2769 )  ;
assign n2771 = ~ ( n2749 ) ;
assign n2772 =  ( n885 ) ^ ( n861 )  ;
assign n2773 =  ( n2772 ) ^ ( n737 )  ;
assign n2774 = ~ ( n462 ) ;
assign n2775 = ~ ( n482 ) ;
assign n2776 =  ( n2774 ) | ( n2775 )  ;
assign n2777 = ~ ( n2776 ) ;
assign n2778 =  ( n2773 ) ^ ( n2777 )  ;
assign n2779 =  ( n2778 ) ^ ( n336 )  ;
assign n2780 =  ( n2779 ) ^ ( n345 )  ;
assign n2781 =  ( n1625 ) | ( n1632 )  ;
assign n2782 =  ( n2781 ) | ( n1668 )  ;
assign n2783 =  ( n2782 ) | ( n1703 )  ;
assign n2784 =  ( n2780 ) ^ ( n2783 )  ;
assign n2785 =  ( n2784 ) ^ ( n1531 )  ;
assign n2786 =  ( n2785 ) ^ ( n1546 )  ;
assign n2787 = ~ ( n2786 ) ;
assign n2788 =  ( n2771 ) | ( n2787 )  ;
assign n2789 =  ( n905 ) ^ ( n843 )  ;
assign n2790 = ~ ( n573 ) ;
assign n2791 = ~ ( n583 ) ;
assign n2792 =  ( n2790 ) | ( n2791 )  ;
assign n2793 = ~ ( n2792 ) ;
assign n2794 =  ( n2789 ) ^ ( n2793 )  ;
assign n2795 =  ( n2794 ) ^ ( n462 )  ;
assign n2796 =  ( n2795 ) ^ ( n482 )  ;
assign n2797 = ~ ( n941 ) ;
assign n2798 = ~ ( n955 ) ;
assign n2799 =  ( n2797 ) | ( n2798 )  ;
assign n2800 =  ( n813 ) ^ ( n823 )  ;
assign n2801 = ~ ( n2800 ) ;
assign n2802 =  ( n2799 ) | ( n2801 )  ;
assign n2803 = ~ ( n966 ) ;
assign n2804 =  ( n2802 ) | ( n2803 )  ;
assign n2805 = ~ ( n982 ) ;
assign n2806 =  ( n2804 ) | ( n2805 )  ;
assign n2807 = ~ ( n2806 ) ;
assign n2808 = ~ ( n1008 ) ;
assign n2809 =  ( n1075 ) | ( n1163 )  ;
assign n2810 =  ( n2809 ) | ( n1250 )  ;
assign n2811 =  ( n2810 ) | ( n1821 )  ;
assign n2812 =  ( n2811 ) | ( n1848 )  ;
assign n2813 = ~ ( n2812 ) ;
assign n2814 =  ( n2808 ) | ( n2813 )  ;
assign n2815 = ~ ( n2814 ) ;
assign n2816 =  ( n2807 ) | ( n2815 )  ;
assign n2817 =  ( n2796 ) ^ ( n2816 )  ;
assign n2818 = ~ ( n2817 ) ;
assign n2819 =  ( n1531 ) ^ ( n1546 )  ;
assign n2820 = ~ ( n2819 ) ;
assign n2821 =  ( n2818 ) | ( n2820 )  ;
assign n2822 = ~ ( n2821 ) ;
assign n2823 =  ( n905 ) ^ ( n843 )  ;
assign n2824 = ~ ( n573 ) ;
assign n2825 = ~ ( n583 ) ;
assign n2826 =  ( n2824 ) | ( n2825 )  ;
assign n2827 = ~ ( n2826 ) ;
assign n2828 =  ( n2823 ) ^ ( n2827 )  ;
assign n2829 =  ( n2828 ) ^ ( n462 )  ;
assign n2830 =  ( n2829 ) ^ ( n482 )  ;
assign n2831 =  ( n2807 ) | ( n2815 )  ;
assign n2832 =  ( n2830 ) ^ ( n2831 )  ;
assign n2833 =  ( n2832 ) ^ ( n1531 )  ;
assign n2834 =  ( n2833 ) ^ ( n1546 )  ;
assign n2835 = ~ ( n2834 ) ;
assign n2836 =  ( n1000 ) ^ ( n975 )  ;
assign n2837 = ~ ( n704 ) ;
assign n2838 = ~ ( n717 ) ;
assign n2839 =  ( n2837 ) | ( n2838 )  ;
assign n2840 = ~ ( n2839 ) ;
assign n2841 =  ( n2836 ) ^ ( n2840 )  ;
assign n2842 =  ( n2841 ) ^ ( n573 )  ;
assign n2843 =  ( n2842 ) ^ ( n583 )  ;
assign n2844 =  ( n1075 ) | ( n1163 )  ;
assign n2845 =  ( n2844 ) | ( n1250 )  ;
assign n2846 =  ( n2845 ) | ( n1821 )  ;
assign n2847 =  ( n2846 ) | ( n1848 )  ;
assign n2848 =  ( n2843 ) ^ ( n2847 )  ;
assign n2849 = ~ ( n2848 ) ;
assign n2850 =  ( n2835 ) | ( n2849 )  ;
assign n2851 =  ( n1531 ) ^ ( n1546 )  ;
assign n2852 = ~ ( n2851 ) ;
assign n2853 =  ( n2850 ) | ( n2852 )  ;
assign n2854 = ~ ( n2853 ) ;
assign n2855 =  ( n2822 ) | ( n2854 )  ;
assign n2856 = ~ ( n2855 ) ;
assign n2857 =  ( n2788 ) | ( n2856 )  ;
assign n2858 = ~ ( n2857 ) ;
assign n2859 =  ( n2770 ) | ( n2858 )  ;
assign n2860 = ~ ( n2749 ) ;
assign n2861 = ~ ( n2786 ) ;
assign n2862 =  ( n2860 ) | ( n2861 )  ;
assign n2863 = ~ ( n2834 ) ;
assign n2864 =  ( n2862 ) | ( n2863 )  ;
assign n2865 =  ( n1000 ) ^ ( n975 )  ;
assign n2866 = ~ ( n704 ) ;
assign n2867 = ~ ( n717 ) ;
assign n2868 =  ( n2866 ) | ( n2867 )  ;
assign n2869 = ~ ( n2868 ) ;
assign n2870 =  ( n2865 ) ^ ( n2869 )  ;
assign n2871 =  ( n2870 ) ^ ( n573 )  ;
assign n2872 =  ( n2871 ) ^ ( n583 )  ;
assign n2873 =  ( n1075 ) | ( n1163 )  ;
assign n2874 =  ( n2873 ) | ( n1250 )  ;
assign n2875 =  ( n2874 ) | ( n1821 )  ;
assign n2876 =  ( n2875 ) | ( n1848 )  ;
assign n2877 =  ( n2872 ) ^ ( n2876 )  ;
assign n2878 =  ( n2877 ) ^ ( n1531 )  ;
assign n2879 =  ( n2878 ) ^ ( n1546 )  ;
assign n2880 = ~ ( n2879 ) ;
assign n2881 =  ( n2864 ) | ( n2880 )  ;
assign n2882 =  ( n1084 ) ^ ( n1065 )  ;
assign n2883 = ~ ( n813 ) ;
assign n2884 = ~ ( n823 ) ;
assign n2885 =  ( n2883 ) | ( n2884 )  ;
assign n2886 = ~ ( n2885 ) ;
assign n2887 =  ( n2882 ) ^ ( n2886 )  ;
assign n2888 =  ( n2887 ) ^ ( n704 )  ;
assign n2889 =  ( n2888 ) ^ ( n717 )  ;
assign n2890 = ~ ( n1119 ) ;
assign n2891 = ~ ( n1133 ) ;
assign n2892 =  ( n2890 ) | ( n2891 )  ;
assign n2893 =  ( n1036 ) ^ ( n1045 )  ;
assign n2894 = ~ ( n2893 ) ;
assign n2895 =  ( n2892 ) | ( n2894 )  ;
assign n2896 = ~ ( n1144 ) ;
assign n2897 =  ( n2895 ) | ( n2896 )  ;
assign n2898 = ~ ( n1160 ) ;
assign n2899 =  ( n2897 ) | ( n2898 )  ;
assign n2900 = ~ ( n2899 ) ;
assign n2901 = ~ ( n1182 ) ;
assign n2902 =  ( n1651 ) | ( n1664 )  ;
assign n2903 =  ( n2902 ) | ( n1973 )  ;
assign n2904 =  ( n2903 ) | ( n1996 )  ;
assign n2905 = ~ ( n2904 ) ;
assign n2906 =  ( n2901 ) | ( n2905 )  ;
assign n2907 = ~ ( n2906 ) ;
assign n2908 =  ( n2900 ) | ( n2907 )  ;
assign n2909 =  ( n2889 ) ^ ( n2908 )  ;
assign n2910 = ~ ( n2909 ) ;
assign n2911 =  ( n1531 ) ^ ( n1546 )  ;
assign n2912 = ~ ( n2911 ) ;
assign n2913 =  ( n2910 ) | ( n2912 )  ;
assign n2914 = ~ ( n2913 ) ;
assign n2915 =  ( n1084 ) ^ ( n1065 )  ;
assign n2916 = ~ ( n813 ) ;
assign n2917 = ~ ( n823 ) ;
assign n2918 =  ( n2916 ) | ( n2917 )  ;
assign n2919 = ~ ( n2918 ) ;
assign n2920 =  ( n2915 ) ^ ( n2919 )  ;
assign n2921 =  ( n2920 ) ^ ( n704 )  ;
assign n2922 =  ( n2921 ) ^ ( n717 )  ;
assign n2923 =  ( n2900 ) | ( n2907 )  ;
assign n2924 =  ( n2922 ) ^ ( n2923 )  ;
assign n2925 =  ( n2924 ) ^ ( n1531 )  ;
assign n2926 =  ( n2925 ) ^ ( n1546 )  ;
assign n2927 = ~ ( n2926 ) ;
assign n2928 =  ( n1174 ) ^ ( n1153 )  ;
assign n2929 = ~ ( n941 ) ;
assign n2930 = ~ ( n955 ) ;
assign n2931 =  ( n2929 ) | ( n2930 )  ;
assign n2932 = ~ ( n2931 ) ;
assign n2933 =  ( n2928 ) ^ ( n2932 )  ;
assign n2934 =  ( n2933 ) ^ ( n813 )  ;
assign n2935 =  ( n2934 ) ^ ( n823 )  ;
assign n2936 =  ( n1651 ) | ( n1664 )  ;
assign n2937 =  ( n2936 ) | ( n1973 )  ;
assign n2938 =  ( n2937 ) | ( n1996 )  ;
assign n2939 =  ( n2935 ) ^ ( n2938 )  ;
assign n2940 = ~ ( n2939 ) ;
assign n2941 =  ( n2927 ) | ( n2940 )  ;
assign n2942 =  ( n1531 ) ^ ( n1546 )  ;
assign n2943 = ~ ( n2942 ) ;
assign n2944 =  ( n2941 ) | ( n2943 )  ;
assign n2945 = ~ ( n2944 ) ;
assign n2946 =  ( n2914 ) | ( n2945 )  ;
assign n2947 = ~ ( n2926 ) ;
assign n2948 =  ( n1174 ) ^ ( n1153 )  ;
assign n2949 = ~ ( n941 ) ;
assign n2950 = ~ ( n955 ) ;
assign n2951 =  ( n2949 ) | ( n2950 )  ;
assign n2952 = ~ ( n2951 ) ;
assign n2953 =  ( n2948 ) ^ ( n2952 )  ;
assign n2954 =  ( n2953 ) ^ ( n813 )  ;
assign n2955 =  ( n2954 ) ^ ( n823 )  ;
assign n2956 =  ( n1651 ) | ( n1664 )  ;
assign n2957 =  ( n2956 ) | ( n1973 )  ;
assign n2958 =  ( n2957 ) | ( n1996 )  ;
assign n2959 =  ( n2955 ) ^ ( n2958 )  ;
assign n2960 =  ( n2959 ) ^ ( n1531 )  ;
assign n2961 =  ( n2960 ) ^ ( n1546 )  ;
assign n2962 = ~ ( n2961 ) ;
assign n2963 =  ( n2947 ) | ( n2962 )  ;
assign n2964 = ~ ( n1036 ) ;
assign n2965 = ~ ( n1045 ) ;
assign n2966 =  ( n2964 ) | ( n2965 )  ;
assign n2967 = ~ ( n2966 ) ;
assign n2968 =  ( n1191 ) ^ ( n2967 )  ;
assign n2969 =  ( n2968 ) ^ ( n941 )  ;
assign n2970 =  ( n2969 ) ^ ( n955 )  ;
assign n2971 = ~ ( n1226 ) ;
assign n2972 = ~ ( n1236 ) ;
assign n2973 =  ( n2971 ) | ( n2972 )  ;
assign n2974 =  ( n1119 ) ^ ( n1133 )  ;
assign n2975 = ~ ( n2974 ) ;
assign n2976 =  ( n2973 ) | ( n2975 )  ;
assign n2977 = ~ ( n1247 ) ;
assign n2978 =  ( n2976 ) | ( n2977 )  ;
assign n2979 = ~ ( n2978 ) ;
assign n2980 = ~ ( n1282 ) ;
assign n2981 =  ( n1337 ) | ( n1454 )  ;
assign n2982 =  ( n2981 ) | ( n1512 )  ;
assign n2983 = ~ ( n2982 ) ;
assign n2984 =  ( n2980 ) | ( n2983 )  ;
assign n2985 = ~ ( n2984 ) ;
assign n2986 =  ( n2979 ) | ( n2985 )  ;
assign n2987 =  ( n2970 ) ^ ( n2986 )  ;
assign n2988 = ~ ( n2987 ) ;
assign n2989 =  ( n1531 ) ^ ( n1546 )  ;
assign n2990 = ~ ( n2989 ) ;
assign n2991 =  ( n2988 ) | ( n2990 )  ;
assign n2992 = ~ ( n2991 ) ;
assign n2993 = ~ ( n1036 ) ;
assign n2994 = ~ ( n1045 ) ;
assign n2995 =  ( n2993 ) | ( n2994 )  ;
assign n2996 = ~ ( n2995 ) ;
assign n2997 =  ( n1191 ) ^ ( n2996 )  ;
assign n2998 =  ( n2997 ) ^ ( n941 )  ;
assign n2999 =  ( n2998 ) ^ ( n955 )  ;
assign n3000 =  ( n2979 ) | ( n2985 )  ;
assign n3001 =  ( n2999 ) ^ ( n3000 )  ;
assign n3002 =  ( n3001 ) ^ ( n1531 )  ;
assign n3003 =  ( n3002 ) ^ ( n1546 )  ;
assign n3004 = ~ ( n3003 ) ;
assign n3005 = ~ ( n1119 ) ;
assign n3006 = ~ ( n1133 ) ;
assign n3007 =  ( n3005 ) | ( n3006 )  ;
assign n3008 = ~ ( n3007 ) ;
assign n3009 =  ( n1275 ) ^ ( n3008 )  ;
assign n3010 =  ( n3009 ) ^ ( n1036 )  ;
assign n3011 =  ( n3010 ) ^ ( n1045 )  ;
assign n3012 =  ( n1337 ) | ( n1454 )  ;
assign n3013 =  ( n3012 ) | ( n1512 )  ;
assign n3014 =  ( n3011 ) ^ ( n3013 )  ;
assign n3015 = ~ ( n3014 ) ;
assign n3016 =  ( n3004 ) | ( n3015 )  ;
assign n3017 =  ( n1531 ) ^ ( n1546 )  ;
assign n3018 = ~ ( n3017 ) ;
assign n3019 =  ( n3016 ) | ( n3018 )  ;
assign n3020 = ~ ( n3019 ) ;
assign n3021 =  ( n2992 ) | ( n3020 )  ;
assign n3022 = ~ ( n3021 ) ;
assign n3023 =  ( n2963 ) | ( n3022 )  ;
assign n3024 = ~ ( n3023 ) ;
assign n3025 =  ( n2946 ) | ( n3024 )  ;
assign n3026 = ~ ( n3025 ) ;
assign n3027 =  ( n2881 ) | ( n3026 )  ;
assign n3028 = ~ ( n3027 ) ;
assign n3029 =  ( n2859 ) | ( n3028 )  ;
assign n3030 = ~ ( n2749 ) ;
assign n3031 = ~ ( n2786 ) ;
assign n3032 =  ( n3030 ) | ( n3031 )  ;
assign n3033 = ~ ( n2834 ) ;
assign n3034 =  ( n3032 ) | ( n3033 )  ;
assign n3035 = ~ ( n2879 ) ;
assign n3036 =  ( n3034 ) | ( n3035 )  ;
assign n3037 = ~ ( n2926 ) ;
assign n3038 =  ( n3036 ) | ( n3037 )  ;
assign n3039 = ~ ( n2961 ) ;
assign n3040 =  ( n3038 ) | ( n3039 )  ;
assign n3041 = ~ ( n3003 ) ;
assign n3042 =  ( n3040 ) | ( n3041 )  ;
assign n3043 = ~ ( n1119 ) ;
assign n3044 = ~ ( n1133 ) ;
assign n3045 =  ( n3043 ) | ( n3044 )  ;
assign n3046 = ~ ( n3045 ) ;
assign n3047 =  ( n1275 ) ^ ( n3046 )  ;
assign n3048 =  ( n3047 ) ^ ( n1036 )  ;
assign n3049 =  ( n3048 ) ^ ( n1045 )  ;
assign n3050 =  ( n1337 ) | ( n1454 )  ;
assign n3051 =  ( n3050 ) | ( n1512 )  ;
assign n3052 =  ( n3049 ) ^ ( n3051 )  ;
assign n3053 =  ( n3052 ) ^ ( n1531 )  ;
assign n3054 =  ( n3053 ) ^ ( n1546 )  ;
assign n3055 = ~ ( n3054 ) ;
assign n3056 =  ( n3042 ) | ( n3055 )  ;
assign n3057 = ~ ( n1226 ) ;
assign n3058 = ~ ( n1236 ) ;
assign n3059 =  ( n3057 ) | ( n3058 )  ;
assign n3060 = ~ ( n3059 ) ;
assign n3061 =  ( n1344 ) ^ ( n3060 )  ;
assign n3062 =  ( n3061 ) ^ ( n1119 )  ;
assign n3063 =  ( n3062 ) ^ ( n1133 )  ;
assign n3064 = ~ ( n1358 ) ;
assign n3065 =  ( n1401 ) | ( n1450 )  ;
assign n3066 =  ( n3065 ) | ( n1699 )  ;
assign n3067 = ~ ( n3066 ) ;
assign n3068 =  ( n3064 ) | ( n3067 )  ;
assign n3069 = ~ ( n3068 ) ;
assign n3070 =  ( n3063 ) ^ ( n3069 )  ;
assign n3071 = ~ ( n3070 ) ;
assign n3072 =  ( n1531 ) ^ ( n1546 )  ;
assign n3073 = ~ ( n3072 ) ;
assign n3074 =  ( n3071 ) | ( n3073 )  ;
assign n3075 = ~ ( n3074 ) ;
assign n3076 = ~ ( n1226 ) ;
assign n3077 = ~ ( n1236 ) ;
assign n3078 =  ( n3076 ) | ( n3077 )  ;
assign n3079 = ~ ( n3078 ) ;
assign n3080 =  ( n1344 ) ^ ( n3079 )  ;
assign n3081 =  ( n3080 ) ^ ( n1119 )  ;
assign n3082 =  ( n3081 ) ^ ( n1133 )  ;
assign n3083 =  ( n3082 ) ^ ( n3069 )  ;
assign n3084 =  ( n3083 ) ^ ( n1531 )  ;
assign n3085 =  ( n3084 ) ^ ( n1546 )  ;
assign n3086 = ~ ( n3085 ) ;
assign n3087 = ~ ( n1310 ) ;
assign n3088 = ~ ( n1323 ) ;
assign n3089 =  ( n3087 ) | ( n3088 )  ;
assign n3090 = ~ ( n3089 ) ;
assign n3091 =  ( n3090 ) ^ ( n1226 )  ;
assign n3092 =  ( n3091 ) ^ ( n1236 )  ;
assign n3093 =  ( n1401 ) | ( n1450 )  ;
assign n3094 =  ( n3093 ) | ( n1699 )  ;
assign n3095 =  ( n3092 ) ^ ( n3094 )  ;
assign n3096 = ~ ( n3095 ) ;
assign n3097 =  ( n3086 ) | ( n3096 )  ;
assign n3098 =  ( n1531 ) ^ ( n1546 )  ;
assign n3099 = ~ ( n3098 ) ;
assign n3100 =  ( n3097 ) | ( n3099 )  ;
assign n3101 = ~ ( n3100 ) ;
assign n3102 =  ( n3075 ) | ( n3101 )  ;
assign n3103 = ~ ( n3085 ) ;
assign n3104 = ~ ( n1310 ) ;
assign n3105 = ~ ( n1323 ) ;
assign n3106 =  ( n3104 ) | ( n3105 )  ;
assign n3107 = ~ ( n3106 ) ;
assign n3108 =  ( n3107 ) ^ ( n1226 )  ;
assign n3109 =  ( n3108 ) ^ ( n1236 )  ;
assign n3110 =  ( n1401 ) | ( n1450 )  ;
assign n3111 =  ( n3110 ) | ( n1699 )  ;
assign n3112 =  ( n3109 ) ^ ( n3111 )  ;
assign n3113 =  ( n3112 ) ^ ( n1531 )  ;
assign n3114 =  ( n3113 ) ^ ( n1546 )  ;
assign n3115 = ~ ( n3114 ) ;
assign n3116 =  ( n3103 ) | ( n3115 )  ;
assign n3117 = ~ ( n1386 ) ;
assign n3118 = ~ ( n1395 ) ;
assign n3119 =  ( n3117 ) | ( n3118 )  ;
assign n3120 = ~ ( n3119 ) ;
assign n3121 =  ( n3120 ) ^ ( n1310 )  ;
assign n3122 =  ( n3121 ) ^ ( n1323 )  ;
assign n3123 = ~ ( n1434 ) ;
assign n3124 = ~ ( n1444 ) ;
assign n3125 =  ( n3123 ) | ( n3124 )  ;
assign n3126 =  ( n1386 ) ^ ( n1395 )  ;
assign n3127 = ~ ( n3126 ) ;
assign n3128 =  ( n3125 ) | ( n3127 )  ;
assign n3129 = ~ ( n3128 ) ;
assign n3130 = ~ ( n1466 ) ;
assign n3131 =  ( n1434 ) ^ ( n1444 )  ;
assign n3132 = ~ ( n3131 ) ;
assign n3133 =  ( n3130 ) | ( n3132 )  ;
assign n3134 = ~ ( n1497 ) ;
assign n3135 =  ( n3133 ) | ( n3134 )  ;
assign n3136 = ~ ( n1506 ) ;
assign n3137 =  ( n3135 ) | ( n3136 )  ;
assign n3138 = ki[1:1] ;
assign n3139 = ~ ( n3138 ) ;
assign n3140 =  ( n3137 ) | ( n3139 )  ;
assign n3141 = ~ ( n3140 ) ;
assign n3142 =  ( n3129 ) | ( n3141 )  ;
assign n3143 =  ( n3122 ) ^ ( n3142 )  ;
assign n3144 = ~ ( n3143 ) ;
assign n3145 =  ( n1531 ) ^ ( n1546 )  ;
assign n3146 = ~ ( n3145 ) ;
assign n3147 =  ( n3144 ) | ( n3146 )  ;
assign n3148 = ~ ( n3147 ) ;
assign n3149 = ~ ( n1386 ) ;
assign n3150 = ~ ( n1395 ) ;
assign n3151 =  ( n3149 ) | ( n3150 )  ;
assign n3152 = ~ ( n3151 ) ;
assign n3153 =  ( n3152 ) ^ ( n1310 )  ;
assign n3154 =  ( n3153 ) ^ ( n1323 )  ;
assign n3155 =  ( n3129 ) | ( n3141 )  ;
assign n3156 =  ( n3154 ) ^ ( n3155 )  ;
assign n3157 =  ( n3156 ) ^ ( n1531 )  ;
assign n3158 =  ( n3157 ) ^ ( n1546 )  ;
assign n3159 = ~ ( n3158 ) ;
assign n3160 = ~ ( n1434 ) ;
assign n3161 = ~ ( n1444 ) ;
assign n3162 =  ( n3160 ) | ( n3161 )  ;
assign n3163 = ~ ( n3162 ) ;
assign n3164 =  ( n3163 ) ^ ( n1386 )  ;
assign n3165 =  ( n3164 ) ^ ( n1395 )  ;
assign n3166 =  ( n1434 ) ^ ( n1444 )  ;
assign n3167 = ~ ( n3166 ) ;
assign n3168 = ~ ( n1497 ) ;
assign n3169 =  ( n3167 ) | ( n3168 )  ;
assign n3170 = ~ ( n1506 ) ;
assign n3171 =  ( n3169 ) | ( n3170 )  ;
assign n3172 = ki[1:1] ;
assign n3173 = ~ ( n3172 ) ;
assign n3174 =  ( n3171 ) | ( n3173 )  ;
assign n3175 = ~ ( n3174 ) ;
assign n3176 =  ( n3165 ) ^ ( n3175 )  ;
assign n3177 = ~ ( n3176 ) ;
assign n3178 =  ( n3159 ) | ( n3177 )  ;
assign n3179 =  ( n1531 ) ^ ( n1546 )  ;
assign n3180 = ~ ( n3179 ) ;
assign n3181 =  ( n3178 ) | ( n3180 )  ;
assign n3182 = ~ ( n3181 ) ;
assign n3183 =  ( n3148 ) | ( n3182 )  ;
assign n3184 = ~ ( n3183 ) ;
assign n3185 =  ( n3116 ) | ( n3184 )  ;
assign n3186 = ~ ( n3185 ) ;
assign n3187 =  ( n3102 ) | ( n3186 )  ;
assign n3188 = ~ ( n3085 ) ;
assign n3189 = ~ ( n3114 ) ;
assign n3190 =  ( n3188 ) | ( n3189 )  ;
assign n3191 = ~ ( n3158 ) ;
assign n3192 =  ( n3190 ) | ( n3191 )  ;
assign n3193 = ~ ( n1434 ) ;
assign n3194 = ~ ( n1444 ) ;
assign n3195 =  ( n3193 ) | ( n3194 )  ;
assign n3196 = ~ ( n3195 ) ;
assign n3197 =  ( n3196 ) ^ ( n1386 )  ;
assign n3198 =  ( n3197 ) ^ ( n1395 )  ;
assign n3199 =  ( n3198 ) ^ ( n3175 )  ;
assign n3200 =  ( n3199 ) ^ ( n1531 )  ;
assign n3201 =  ( n3200 ) ^ ( n1546 )  ;
assign n3202 = ~ ( n3201 ) ;
assign n3203 =  ( n3192 ) | ( n3202 )  ;
assign n3204 =  ( n1434 ) ^ ( n1444 )  ;
assign n3205 = ~ ( n1497 ) ;
assign n3206 = ~ ( n1506 ) ;
assign n3207 =  ( n3205 ) | ( n3206 )  ;
assign n3208 = ki[1:1] ;
assign n3209 = ~ ( n3208 ) ;
assign n3210 =  ( n3207 ) | ( n3209 )  ;
assign n3211 = ~ ( n3210 ) ;
assign n3212 =  ( n3204 ) ^ ( n3211 )  ;
assign n3213 = ~ ( n3212 ) ;
assign n3214 =  ( n1531 ) ^ ( n1546 )  ;
assign n3215 = ~ ( n3214 ) ;
assign n3216 =  ( n3213 ) | ( n3215 )  ;
assign n3217 = ~ ( n3216 ) ;
assign n3218 =  ( n1434 ) ^ ( n1444 )  ;
assign n3219 =  ( n3218 ) ^ ( n3211 )  ;
assign n3220 =  ( n3219 ) ^ ( n1531 )  ;
assign n3221 =  ( n3220 ) ^ ( n1546 )  ;
assign n3222 = ~ ( n3221 ) ;
assign n3223 = ~ ( n1506 ) ;
assign n3224 = ki[1:1] ;
assign n3225 = ~ ( n3224 ) ;
assign n3226 =  ( n3223 ) | ( n3225 )  ;
assign n3227 = ~ ( n3226 ) ;
assign n3228 =  ( n1497 ) ^ ( n3227 )  ;
assign n3229 = ~ ( n3228 ) ;
assign n3230 =  ( n3222 ) | ( n3229 )  ;
assign n3231 = ~ ( n1540 ) ;
assign n3232 = kd[1:1] ;
assign n3233 = ~ ( n3232 ) ;
assign n3234 =  ( n3231 ) | ( n3233 )  ;
assign n3235 = ~ ( n3234 ) ;
assign n3236 =  ( n1531 ) ^ ( n3235 )  ;
assign n3237 = ~ ( n3236 ) ;
assign n3238 =  ( n3230 ) | ( n3237 )  ;
assign n3239 = ~ ( n3238 ) ;
assign n3240 =  ( n3217 ) | ( n3239 )  ;
assign n3241 =  ( n1434 ) ^ ( n1444 )  ;
assign n3242 =  ( n3241 ) ^ ( n3211 )  ;
assign n3243 =  ( n3242 ) ^ ( n1531 )  ;
assign n3244 =  ( n3243 ) ^ ( n1546 )  ;
assign n3245 = ~ ( n3244 ) ;
assign n3246 =  ( n1497 ) ^ ( n3227 )  ;
assign n3247 =  ( n3246 ) ^ ( n1531 )  ;
assign n3248 =  ( n3247 ) ^ ( n3235 )  ;
assign n3249 = ~ ( n3248 ) ;
assign n3250 =  ( n3245 ) | ( n3249 )  ;
assign n3251 = ki[1:1] ;
assign n3252 =  ( n1506 ) ^ ( n3251 )  ;
assign n3253 = ~ ( n3252 ) ;
assign n3254 =  ( n3250 ) | ( n3253 )  ;
assign n3255 = kd[1:1] ;
assign n3256 =  ( n1540 ) ^ ( n3255 )  ;
assign n3257 = ~ ( n3256 ) ;
assign n3258 =  ( n3254 ) | ( n3257 )  ;
assign n3259 = ~ ( n3258 ) ;
assign n3260 =  ( n3240 ) | ( n3259 )  ;
assign n3261 = ~ ( n3260 ) ;
assign n3262 =  ( n3203 ) | ( n3261 )  ;
assign n3263 = ~ ( n3262 ) ;
assign n3264 =  ( n3187 ) | ( n3263 )  ;
assign n3265 = ~ ( n3264 ) ;
assign n3266 =  ( n3056 ) | ( n3265 )  ;
assign n3267 = ~ ( n3266 ) ;
assign n3268 =  ( n3029 ) | ( n3267 )  ;
assign n3269 = ~ ( n3268 ) ;
assign n3270 =  ( n2700 ) | ( n3269 )  ;
assign n3271 = ~ ( n3270 ) ;
assign n3272 =  ( n2663 ) | ( n3271 )  ;
assign n3273 =  ( n1549 ) ^ ( n3272 )  ;
assign n3274 = ~ ( n1723 ) ;
assign n3275 = ~ ( n1531 ) ;
assign n3276 =  ( n3275 ) | ( n1546 )  ;
assign n3277 = ~ ( n3276 ) ;
assign n3278 =  ( n3274 ) ^ ( n3277 )  ;
assign n3279 = ~ ( n1711 ) ;
assign n3280 = ~ ( n1728 ) ;
assign n3281 = ~ ( n1856 ) ;
assign n3282 = ~ ( n1885 ) ;
assign n3283 =  ( n3281 ) | ( n3282 )  ;
assign n3284 = ~ ( n1871 ) ;
assign n3285 = ~ ( n2004 ) ;
assign n3286 = ~ ( n2037 ) ;
assign n3287 =  ( n3285 ) | ( n3286 )  ;
assign n3288 = ~ ( n3287 ) ;
assign n3289 =  ( n3284 ) | ( n3288 )  ;
assign n3290 = ~ ( n3289 ) ;
assign n3291 =  ( n3283 ) | ( n3290 )  ;
assign n3292 = ~ ( n1871 ) ;
assign n3293 = ~ ( n2021 ) ;
assign n3294 =  ( n3292 ) | ( n3293 )  ;
assign n3295 = ~ ( n2113 ) ;
assign n3296 = ~ ( n2146 ) ;
assign n3297 =  ( n3295 ) | ( n3296 )  ;
assign n3298 = ~ ( n2130 ) ;
assign n3299 = ~ ( n2245 ) ;
assign n3300 = ~ ( n2282 ) ;
assign n3301 =  ( n3299 ) | ( n3300 )  ;
assign n3302 = ~ ( n3301 ) ;
assign n3303 =  ( n3298 ) | ( n3302 )  ;
assign n3304 = ~ ( n3303 ) ;
assign n3305 =  ( n3297 ) | ( n3304 )  ;
assign n3306 = ~ ( n3305 ) ;
assign n3307 =  ( n3294 ) | ( n3306 )  ;
assign n3308 = ~ ( n3307 ) ;
assign n3309 =  ( n3291 ) | ( n3308 )  ;
assign n3310 = ~ ( n1871 ) ;
assign n3311 = ~ ( n2021 ) ;
assign n3312 =  ( n3310 ) | ( n3311 )  ;
assign n3313 = ~ ( n2130 ) ;
assign n3314 =  ( n3312 ) | ( n3313 )  ;
assign n3315 = ~ ( n2264 ) ;
assign n3316 =  ( n3314 ) | ( n3315 )  ;
assign n3317 = ~ ( n1531 ) ;
assign n3318 =  ( n2393 ) | ( n3317 )  ;
assign n3319 =  ( n3318 ) | ( n1546 )  ;
assign n3320 = ~ ( n3319 ) ;
assign n3321 = ~ ( n2404 ) ;
assign n3322 =  ( n3321 ) | ( n2411 )  ;
assign n3323 = ~ ( n1531 ) ;
assign n3324 =  ( n3322 ) | ( n3323 )  ;
assign n3325 =  ( n3324 ) | ( n1546 )  ;
assign n3326 = ~ ( n3325 ) ;
assign n3327 =  ( n3320 ) | ( n3326 )  ;
assign n3328 = ~ ( n2404 ) ;
assign n3329 = ~ ( n2433 ) ;
assign n3330 =  ( n3328 ) | ( n3329 )  ;
assign n3331 = ~ ( n2518 ) ;
assign n3332 =  ( n3331 ) | ( n2553 )  ;
assign n3333 = ~ ( n3332 ) ;
assign n3334 =  ( n3330 ) | ( n3333 )  ;
assign n3335 = ~ ( n3334 ) ;
assign n3336 =  ( n3327 ) | ( n3335 )  ;
assign n3337 = ~ ( n2404 ) ;
assign n3338 = ~ ( n2433 ) ;
assign n3339 =  ( n3337 ) | ( n3338 )  ;
assign n3340 = ~ ( n2530 ) ;
assign n3341 =  ( n3339 ) | ( n3340 )  ;
assign n3342 = ~ ( n2573 ) ;
assign n3343 =  ( n3341 ) | ( n3342 )  ;
assign n3344 =  ( n2614 ) | ( n2650 )  ;
assign n3345 = ~ ( n2629 ) ;
assign n3346 = ~ ( n2698 ) ;
assign n3347 =  ( n3345 ) | ( n3346 )  ;
assign n3348 =  ( n2736 ) | ( n2769 )  ;
assign n3349 = ~ ( n3348 ) ;
assign n3350 =  ( n3347 ) | ( n3349 )  ;
assign n3351 = ~ ( n3350 ) ;
assign n3352 =  ( n3344 ) | ( n3351 )  ;
assign n3353 = ~ ( n3352 ) ;
assign n3354 =  ( n3343 ) | ( n3353 )  ;
assign n3355 = ~ ( n3354 ) ;
assign n3356 =  ( n3336 ) | ( n3355 )  ;
assign n3357 = ~ ( n3356 ) ;
assign n3358 =  ( n3316 ) | ( n3357 )  ;
assign n3359 = ~ ( n3358 ) ;
assign n3360 =  ( n3309 ) | ( n3359 )  ;
assign n3361 = ~ ( n1871 ) ;
assign n3362 = ~ ( n2021 ) ;
assign n3363 =  ( n3361 ) | ( n3362 )  ;
assign n3364 = ~ ( n2130 ) ;
assign n3365 =  ( n3363 ) | ( n3364 )  ;
assign n3366 = ~ ( n2264 ) ;
assign n3367 =  ( n3365 ) | ( n3366 )  ;
assign n3368 = ~ ( n2404 ) ;
assign n3369 =  ( n3367 ) | ( n3368 )  ;
assign n3370 = ~ ( n2433 ) ;
assign n3371 =  ( n3369 ) | ( n3370 )  ;
assign n3372 = ~ ( n2530 ) ;
assign n3373 =  ( n3371 ) | ( n3372 )  ;
assign n3374 = ~ ( n2573 ) ;
assign n3375 =  ( n3373 ) | ( n3374 )  ;
assign n3376 = ~ ( n2629 ) ;
assign n3377 =  ( n3375 ) | ( n3376 )  ;
assign n3378 = ~ ( n2698 ) ;
assign n3379 =  ( n3377 ) | ( n3378 )  ;
assign n3380 = ~ ( n2749 ) ;
assign n3381 =  ( n3379 ) | ( n3380 )  ;
assign n3382 = ~ ( n2786 ) ;
assign n3383 =  ( n3381 ) | ( n3382 )  ;
assign n3384 =  ( n2822 ) | ( n2854 )  ;
assign n3385 = ~ ( n2834 ) ;
assign n3386 = ~ ( n2879 ) ;
assign n3387 =  ( n3385 ) | ( n3386 )  ;
assign n3388 =  ( n2914 ) | ( n2945 )  ;
assign n3389 = ~ ( n3388 ) ;
assign n3390 =  ( n3387 ) | ( n3389 )  ;
assign n3391 = ~ ( n3390 ) ;
assign n3392 =  ( n3384 ) | ( n3391 )  ;
assign n3393 = ~ ( n2834 ) ;
assign n3394 = ~ ( n2879 ) ;
assign n3395 =  ( n3393 ) | ( n3394 )  ;
assign n3396 = ~ ( n2926 ) ;
assign n3397 =  ( n3395 ) | ( n3396 )  ;
assign n3398 = ~ ( n2961 ) ;
assign n3399 =  ( n3397 ) | ( n3398 )  ;
assign n3400 =  ( n2992 ) | ( n3020 )  ;
assign n3401 = ~ ( n3003 ) ;
assign n3402 = ~ ( n3054 ) ;
assign n3403 =  ( n3401 ) | ( n3402 )  ;
assign n3404 =  ( n3075 ) | ( n3101 )  ;
assign n3405 = ~ ( n3404 ) ;
assign n3406 =  ( n3403 ) | ( n3405 )  ;
assign n3407 = ~ ( n3406 ) ;
assign n3408 =  ( n3400 ) | ( n3407 )  ;
assign n3409 = ~ ( n3408 ) ;
assign n3410 =  ( n3399 ) | ( n3409 )  ;
assign n3411 = ~ ( n3410 ) ;
assign n3412 =  ( n3392 ) | ( n3411 )  ;
assign n3413 = ~ ( n2834 ) ;
assign n3414 = ~ ( n2879 ) ;
assign n3415 =  ( n3413 ) | ( n3414 )  ;
assign n3416 = ~ ( n2926 ) ;
assign n3417 =  ( n3415 ) | ( n3416 )  ;
assign n3418 = ~ ( n2961 ) ;
assign n3419 =  ( n3417 ) | ( n3418 )  ;
assign n3420 = ~ ( n3003 ) ;
assign n3421 =  ( n3419 ) | ( n3420 )  ;
assign n3422 = ~ ( n3054 ) ;
assign n3423 =  ( n3421 ) | ( n3422 )  ;
assign n3424 = ~ ( n3085 ) ;
assign n3425 =  ( n3423 ) | ( n3424 )  ;
assign n3426 = ~ ( n3114 ) ;
assign n3427 =  ( n3425 ) | ( n3426 )  ;
assign n3428 =  ( n3148 ) | ( n3182 )  ;
assign n3429 = ~ ( n3158 ) ;
assign n3430 = ~ ( n3201 ) ;
assign n3431 =  ( n3429 ) | ( n3430 )  ;
assign n3432 =  ( n3217 ) | ( n3239 )  ;
assign n3433 = ~ ( n3432 ) ;
assign n3434 =  ( n3431 ) | ( n3433 )  ;
assign n3435 = ~ ( n3434 ) ;
assign n3436 =  ( n3428 ) | ( n3435 )  ;
assign n3437 = ~ ( n3158 ) ;
assign n3438 = ~ ( n3201 ) ;
assign n3439 =  ( n3437 ) | ( n3438 )  ;
assign n3440 =  ( n1434 ) ^ ( n1444 )  ;
assign n3441 =  ( n3440 ) ^ ( n3211 )  ;
assign n3442 =  ( n3441 ) ^ ( n1531 )  ;
assign n3443 =  ( n3442 ) ^ ( n1546 )  ;
assign n3444 = ~ ( n3443 ) ;
assign n3445 =  ( n3439 ) | ( n3444 )  ;
assign n3446 =  ( n1497 ) ^ ( n3227 )  ;
assign n3447 =  ( n3446 ) ^ ( n1531 )  ;
assign n3448 =  ( n3447 ) ^ ( n3235 )  ;
assign n3449 = ~ ( n3448 ) ;
assign n3450 =  ( n3445 ) | ( n3449 )  ;
assign n3451 = ki[1:1] ;
assign n3452 =  ( n1506 ) ^ ( n3451 )  ;
assign n3453 = ~ ( n3452 ) ;
assign n3454 =  ( n3450 ) | ( n3453 )  ;
assign n3455 = kd[1:1] ;
assign n3456 =  ( n1540 ) ^ ( n3455 )  ;
assign n3457 = ~ ( n3456 ) ;
assign n3458 =  ( n3454 ) | ( n3457 )  ;
assign n3459 = ~ ( n3458 ) ;
assign n3460 =  ( n3436 ) | ( n3459 )  ;
assign n3461 = ~ ( n3460 ) ;
assign n3462 =  ( n3427 ) | ( n3461 )  ;
assign n3463 = ~ ( n3462 ) ;
assign n3464 =  ( n3412 ) | ( n3463 )  ;
assign n3465 = ~ ( n3464 ) ;
assign n3466 =  ( n3383 ) | ( n3465 )  ;
assign n3467 = ~ ( n3466 ) ;
assign n3468 =  ( n3360 ) | ( n3467 )  ;
assign n3469 = ~ ( n3468 ) ;
assign n3470 =  ( n3280 ) | ( n3469 )  ;
assign n3471 = ~ ( n3470 ) ;
assign n3472 =  ( n3279 ) | ( n3471 )  ;
assign n3473 =  ( n3278 ) ^ ( n3472 )  ;
assign n3474 =  { ( n3273 ) , ( n3473 ) }  ;
assign n3475 = ~ ( n1723 ) ;
assign n3476 = ~ ( n1531 ) ;
assign n3477 =  ( n3476 ) | ( n1546 )  ;
assign n3478 = ~ ( n3477 ) ;
assign n3479 =  ( n3475 ) ^ ( n3478 )  ;
assign n3480 =  ( n3479 ) ^ ( n3468 )  ;
assign n3481 =  { ( n3474 ) , ( n3480 ) }  ;
assign n3482 = ~ ( n1866 ) ;
assign n3483 = ~ ( n1531 ) ;
assign n3484 =  ( n3483 ) | ( n1546 )  ;
assign n3485 = ~ ( n3484 ) ;
assign n3486 =  ( n3482 ) ^ ( n3485 )  ;
assign n3487 = ~ ( n1856 ) ;
assign n3488 = ~ ( n1871 ) ;
assign n3489 = ~ ( n2004 ) ;
assign n3490 = ~ ( n2037 ) ;
assign n3491 =  ( n3489 ) | ( n3490 )  ;
assign n3492 = ~ ( n2150 ) ;
assign n3493 =  ( n3491 ) | ( n3492 )  ;
assign n3494 = ~ ( n2021 ) ;
assign n3495 = ~ ( n2130 ) ;
assign n3496 =  ( n3494 ) | ( n3495 )  ;
assign n3497 = ~ ( n2245 ) ;
assign n3498 = ~ ( n2282 ) ;
assign n3499 =  ( n3497 ) | ( n3498 )  ;
assign n3500 = ~ ( n2264 ) ;
assign n3501 = ~ ( n2417 ) ;
assign n3502 =  ( n3500 ) | ( n3501 )  ;
assign n3503 = ~ ( n3502 ) ;
assign n3504 =  ( n3499 ) | ( n3503 )  ;
assign n3505 = ~ ( n3504 ) ;
assign n3506 =  ( n3496 ) | ( n3505 )  ;
assign n3507 = ~ ( n3506 ) ;
assign n3508 =  ( n3493 ) | ( n3507 )  ;
assign n3509 = ~ ( n2021 ) ;
assign n3510 = ~ ( n2130 ) ;
assign n3511 =  ( n3509 ) | ( n3510 )  ;
assign n3512 = ~ ( n2264 ) ;
assign n3513 =  ( n3511 ) | ( n3512 )  ;
assign n3514 = ~ ( n2404 ) ;
assign n3515 =  ( n3513 ) | ( n3514 )  ;
assign n3516 = ~ ( n2433 ) ;
assign n3517 =  ( n3515 ) | ( n3516 )  ;
assign n3518 = ~ ( n2518 ) ;
assign n3519 =  ( n3518 ) | ( n2553 )  ;
assign n3520 =  ( n3519 ) | ( n2654 )  ;
assign n3521 = ~ ( n2530 ) ;
assign n3522 = ~ ( n2573 ) ;
assign n3523 =  ( n3521 ) | ( n3522 )  ;
assign n3524 = ~ ( n2629 ) ;
assign n3525 =  ( n3523 ) | ( n3524 )  ;
assign n3526 = ~ ( n2698 ) ;
assign n3527 =  ( n3525 ) | ( n3526 )  ;
assign n3528 =  ( n2736 ) | ( n2769 )  ;
assign n3529 =  ( n3528 ) | ( n2858 )  ;
assign n3530 = ~ ( n3529 ) ;
assign n3531 =  ( n3527 ) | ( n3530 )  ;
assign n3532 = ~ ( n3531 ) ;
assign n3533 =  ( n3520 ) | ( n3532 )  ;
assign n3534 = ~ ( n3533 ) ;
assign n3535 =  ( n3517 ) | ( n3534 )  ;
assign n3536 = ~ ( n3535 ) ;
assign n3537 =  ( n3508 ) | ( n3536 )  ;
assign n3538 = ~ ( n2021 ) ;
assign n3539 = ~ ( n2130 ) ;
assign n3540 =  ( n3538 ) | ( n3539 )  ;
assign n3541 = ~ ( n2264 ) ;
assign n3542 =  ( n3540 ) | ( n3541 )  ;
assign n3543 = ~ ( n2404 ) ;
assign n3544 =  ( n3542 ) | ( n3543 )  ;
assign n3545 = ~ ( n2433 ) ;
assign n3546 =  ( n3544 ) | ( n3545 )  ;
assign n3547 = ~ ( n2530 ) ;
assign n3548 =  ( n3546 ) | ( n3547 )  ;
assign n3549 = ~ ( n2573 ) ;
assign n3550 =  ( n3548 ) | ( n3549 )  ;
assign n3551 = ~ ( n2629 ) ;
assign n3552 =  ( n3550 ) | ( n3551 )  ;
assign n3553 = ~ ( n2698 ) ;
assign n3554 =  ( n3552 ) | ( n3553 )  ;
assign n3555 = ~ ( n2749 ) ;
assign n3556 =  ( n3554 ) | ( n3555 )  ;
assign n3557 = ~ ( n2786 ) ;
assign n3558 =  ( n3556 ) | ( n3557 )  ;
assign n3559 = ~ ( n2834 ) ;
assign n3560 =  ( n3558 ) | ( n3559 )  ;
assign n3561 = ~ ( n2879 ) ;
assign n3562 =  ( n3560 ) | ( n3561 )  ;
assign n3563 =  ( n2914 ) | ( n2945 )  ;
assign n3564 =  ( n3563 ) | ( n3024 )  ;
assign n3565 = ~ ( n2926 ) ;
assign n3566 = ~ ( n2961 ) ;
assign n3567 =  ( n3565 ) | ( n3566 )  ;
assign n3568 = ~ ( n3003 ) ;
assign n3569 =  ( n3567 ) | ( n3568 )  ;
assign n3570 = ~ ( n3054 ) ;
assign n3571 =  ( n3569 ) | ( n3570 )  ;
assign n3572 =  ( n3075 ) | ( n3101 )  ;
assign n3573 =  ( n3572 ) | ( n3186 )  ;
assign n3574 = ~ ( n3573 ) ;
assign n3575 =  ( n3571 ) | ( n3574 )  ;
assign n3576 = ~ ( n3575 ) ;
assign n3577 =  ( n3564 ) | ( n3576 )  ;
assign n3578 = ~ ( n2926 ) ;
assign n3579 = ~ ( n2961 ) ;
assign n3580 =  ( n3578 ) | ( n3579 )  ;
assign n3581 = ~ ( n3003 ) ;
assign n3582 =  ( n3580 ) | ( n3581 )  ;
assign n3583 = ~ ( n3054 ) ;
assign n3584 =  ( n3582 ) | ( n3583 )  ;
assign n3585 = ~ ( n3085 ) ;
assign n3586 =  ( n3584 ) | ( n3585 )  ;
assign n3587 = ~ ( n3114 ) ;
assign n3588 =  ( n3586 ) | ( n3587 )  ;
assign n3589 = ~ ( n3158 ) ;
assign n3590 =  ( n3588 ) | ( n3589 )  ;
assign n3591 = ~ ( n3201 ) ;
assign n3592 =  ( n3590 ) | ( n3591 )  ;
assign n3593 =  ( n3217 ) | ( n3239 )  ;
assign n3594 = ~ ( n3258 ) ;
assign n3595 =  ( n3593 ) | ( n3594 )  ;
assign n3596 = ~ ( n3595 ) ;
assign n3597 =  ( n3592 ) | ( n3596 )  ;
assign n3598 = ~ ( n3597 ) ;
assign n3599 =  ( n3577 ) | ( n3598 )  ;
assign n3600 = ~ ( n3599 ) ;
assign n3601 =  ( n3562 ) | ( n3600 )  ;
assign n3602 = ~ ( n3601 ) ;
assign n3603 =  ( n3537 ) | ( n3602 )  ;
assign n3604 = ~ ( n3603 ) ;
assign n3605 =  ( n3488 ) | ( n3604 )  ;
assign n3606 = ~ ( n3605 ) ;
assign n3607 =  ( n3487 ) | ( n3606 )  ;
assign n3608 =  ( n3486 ) ^ ( n3607 )  ;
assign n3609 =  { ( n3481 ) , ( n3608 ) }  ;
assign n3610 = ~ ( n1866 ) ;
assign n3611 = ~ ( n1531 ) ;
assign n3612 =  ( n3611 ) | ( n1546 )  ;
assign n3613 = ~ ( n3612 ) ;
assign n3614 =  ( n3610 ) ^ ( n3613 )  ;
assign n3615 =  ( n3614 ) ^ ( n3603 )  ;
assign n3616 =  { ( n3609 ) , ( n3615 ) }  ;
assign n3617 = ~ ( n2016 ) ;
assign n3618 = ~ ( n1531 ) ;
assign n3619 =  ( n3618 ) | ( n1546 )  ;
assign n3620 = ~ ( n3619 ) ;
assign n3621 =  ( n3617 ) ^ ( n3620 )  ;
assign n3622 = ~ ( n2004 ) ;
assign n3623 = ~ ( n2021 ) ;
assign n3624 = ~ ( n2113 ) ;
assign n3625 = ~ ( n2146 ) ;
assign n3626 =  ( n3624 ) | ( n3625 )  ;
assign n3627 = ~ ( n3303 ) ;
assign n3628 =  ( n3626 ) | ( n3627 )  ;
assign n3629 = ~ ( n2130 ) ;
assign n3630 = ~ ( n2264 ) ;
assign n3631 =  ( n3629 ) | ( n3630 )  ;
assign n3632 = ~ ( n1531 ) ;
assign n3633 =  ( n2393 ) | ( n3632 )  ;
assign n3634 =  ( n3633 ) | ( n1546 )  ;
assign n3635 = ~ ( n3634 ) ;
assign n3636 = ~ ( n2404 ) ;
assign n3637 =  ( n3636 ) | ( n2411 )  ;
assign n3638 = ~ ( n1531 ) ;
assign n3639 =  ( n3637 ) | ( n3638 )  ;
assign n3640 =  ( n3639 ) | ( n1546 )  ;
assign n3641 = ~ ( n3640 ) ;
assign n3642 =  ( n3635 ) | ( n3641 )  ;
assign n3643 = ~ ( n3334 ) ;
assign n3644 =  ( n3642 ) | ( n3643 )  ;
assign n3645 = ~ ( n3644 ) ;
assign n3646 =  ( n3631 ) | ( n3645 )  ;
assign n3647 = ~ ( n3646 ) ;
assign n3648 =  ( n3628 ) | ( n3647 )  ;
assign n3649 = ~ ( n2130 ) ;
assign n3650 = ~ ( n2264 ) ;
assign n3651 =  ( n3649 ) | ( n3650 )  ;
assign n3652 = ~ ( n2404 ) ;
assign n3653 =  ( n3651 ) | ( n3652 )  ;
assign n3654 = ~ ( n2433 ) ;
assign n3655 =  ( n3653 ) | ( n3654 )  ;
assign n3656 = ~ ( n2530 ) ;
assign n3657 =  ( n3655 ) | ( n3656 )  ;
assign n3658 = ~ ( n2573 ) ;
assign n3659 =  ( n3657 ) | ( n3658 )  ;
assign n3660 =  ( n2614 ) | ( n2650 )  ;
assign n3661 =  ( n3660 ) | ( n3351 )  ;
assign n3662 = ~ ( n2629 ) ;
assign n3663 = ~ ( n2698 ) ;
assign n3664 =  ( n3662 ) | ( n3663 )  ;
assign n3665 = ~ ( n2749 ) ;
assign n3666 =  ( n3664 ) | ( n3665 )  ;
assign n3667 = ~ ( n2786 ) ;
assign n3668 =  ( n3666 ) | ( n3667 )  ;
assign n3669 =  ( n2822 ) | ( n2854 )  ;
assign n3670 =  ( n3669 ) | ( n3391 )  ;
assign n3671 = ~ ( n3670 ) ;
assign n3672 =  ( n3668 ) | ( n3671 )  ;
assign n3673 = ~ ( n3672 ) ;
assign n3674 =  ( n3661 ) | ( n3673 )  ;
assign n3675 = ~ ( n3674 ) ;
assign n3676 =  ( n3659 ) | ( n3675 )  ;
assign n3677 = ~ ( n3676 ) ;
assign n3678 =  ( n3648 ) | ( n3677 )  ;
assign n3679 = ~ ( n2130 ) ;
assign n3680 = ~ ( n2264 ) ;
assign n3681 =  ( n3679 ) | ( n3680 )  ;
assign n3682 = ~ ( n2404 ) ;
assign n3683 =  ( n3681 ) | ( n3682 )  ;
assign n3684 = ~ ( n2433 ) ;
assign n3685 =  ( n3683 ) | ( n3684 )  ;
assign n3686 = ~ ( n2530 ) ;
assign n3687 =  ( n3685 ) | ( n3686 )  ;
assign n3688 = ~ ( n2573 ) ;
assign n3689 =  ( n3687 ) | ( n3688 )  ;
assign n3690 = ~ ( n2629 ) ;
assign n3691 =  ( n3689 ) | ( n3690 )  ;
assign n3692 = ~ ( n2698 ) ;
assign n3693 =  ( n3691 ) | ( n3692 )  ;
assign n3694 = ~ ( n2749 ) ;
assign n3695 =  ( n3693 ) | ( n3694 )  ;
assign n3696 = ~ ( n2786 ) ;
assign n3697 =  ( n3695 ) | ( n3696 )  ;
assign n3698 = ~ ( n2834 ) ;
assign n3699 =  ( n3697 ) | ( n3698 )  ;
assign n3700 = ~ ( n2879 ) ;
assign n3701 =  ( n3699 ) | ( n3700 )  ;
assign n3702 = ~ ( n2926 ) ;
assign n3703 =  ( n3701 ) | ( n3702 )  ;
assign n3704 = ~ ( n2961 ) ;
assign n3705 =  ( n3703 ) | ( n3704 )  ;
assign n3706 =  ( n2992 ) | ( n3020 )  ;
assign n3707 =  ( n3706 ) | ( n3407 )  ;
assign n3708 = ~ ( n3003 ) ;
assign n3709 = ~ ( n3054 ) ;
assign n3710 =  ( n3708 ) | ( n3709 )  ;
assign n3711 = ~ ( n3085 ) ;
assign n3712 =  ( n3710 ) | ( n3711 )  ;
assign n3713 = ~ ( n3114 ) ;
assign n3714 =  ( n3712 ) | ( n3713 )  ;
assign n3715 =  ( n3148 ) | ( n3182 )  ;
assign n3716 =  ( n3715 ) | ( n3435 )  ;
assign n3717 = ~ ( n3716 ) ;
assign n3718 =  ( n3714 ) | ( n3717 )  ;
assign n3719 = ~ ( n3718 ) ;
assign n3720 =  ( n3707 ) | ( n3719 )  ;
assign n3721 = ~ ( n3003 ) ;
assign n3722 = ~ ( n3054 ) ;
assign n3723 =  ( n3721 ) | ( n3722 )  ;
assign n3724 = ~ ( n3085 ) ;
assign n3725 =  ( n3723 ) | ( n3724 )  ;
assign n3726 = ~ ( n3114 ) ;
assign n3727 =  ( n3725 ) | ( n3726 )  ;
assign n3728 = ~ ( n3158 ) ;
assign n3729 =  ( n3727 ) | ( n3728 )  ;
assign n3730 = ~ ( n3201 ) ;
assign n3731 =  ( n3729 ) | ( n3730 )  ;
assign n3732 =  ( n1434 ) ^ ( n1444 )  ;
assign n3733 =  ( n3732 ) ^ ( n3211 )  ;
assign n3734 =  ( n3733 ) ^ ( n1531 )  ;
assign n3735 =  ( n3734 ) ^ ( n1546 )  ;
assign n3736 = ~ ( n3735 ) ;
assign n3737 =  ( n3731 ) | ( n3736 )  ;
assign n3738 =  ( n1497 ) ^ ( n3227 )  ;
assign n3739 =  ( n3738 ) ^ ( n1531 )  ;
assign n3740 =  ( n3739 ) ^ ( n3235 )  ;
assign n3741 = ~ ( n3740 ) ;
assign n3742 =  ( n3737 ) | ( n3741 )  ;
assign n3743 = ki[1:1] ;
assign n3744 =  ( n1506 ) ^ ( n3743 )  ;
assign n3745 = ~ ( n3744 ) ;
assign n3746 =  ( n3742 ) | ( n3745 )  ;
assign n3747 = kd[1:1] ;
assign n3748 =  ( n1540 ) ^ ( n3747 )  ;
assign n3749 = ~ ( n3748 ) ;
assign n3750 =  ( n3746 ) | ( n3749 )  ;
assign n3751 = ~ ( n3750 ) ;
assign n3752 =  ( n3720 ) | ( n3751 )  ;
assign n3753 = ~ ( n3752 ) ;
assign n3754 =  ( n3705 ) | ( n3753 )  ;
assign n3755 = ~ ( n3754 ) ;
assign n3756 =  ( n3678 ) | ( n3755 )  ;
assign n3757 = ~ ( n3756 ) ;
assign n3758 =  ( n3623 ) | ( n3757 )  ;
assign n3759 = ~ ( n3758 ) ;
assign n3760 =  ( n3622 ) | ( n3759 )  ;
assign n3761 =  ( n3621 ) ^ ( n3760 )  ;
assign n3762 =  { ( n3616 ) , ( n3761 ) }  ;
assign n3763 = ~ ( n2016 ) ;
assign n3764 = ~ ( n1531 ) ;
assign n3765 =  ( n3764 ) | ( n1546 )  ;
assign n3766 = ~ ( n3765 ) ;
assign n3767 =  ( n3763 ) ^ ( n3766 )  ;
assign n3768 =  ( n3767 ) ^ ( n3756 )  ;
assign n3769 =  { ( n3762 ) , ( n3768 ) }  ;
assign n3770 = ~ ( n2125 ) ;
assign n3771 = ~ ( n1531 ) ;
assign n3772 =  ( n3771 ) | ( n1546 )  ;
assign n3773 = ~ ( n3772 ) ;
assign n3774 =  ( n3770 ) ^ ( n3773 )  ;
assign n3775 = ~ ( n2113 ) ;
assign n3776 = ~ ( n2130 ) ;
assign n3777 = ~ ( n2245 ) ;
assign n3778 = ~ ( n2282 ) ;
assign n3779 =  ( n3777 ) | ( n3778 )  ;
assign n3780 = ~ ( n2264 ) ;
assign n3781 = ~ ( n2417 ) ;
assign n3782 =  ( n3780 ) | ( n3781 )  ;
assign n3783 = ~ ( n3782 ) ;
assign n3784 =  ( n3779 ) | ( n3783 )  ;
assign n3785 = ~ ( n2657 ) ;
assign n3786 =  ( n3784 ) | ( n3785 )  ;
assign n3787 = ~ ( n2264 ) ;
assign n3788 = ~ ( n2404 ) ;
assign n3789 =  ( n3787 ) | ( n3788 )  ;
assign n3790 = ~ ( n2433 ) ;
assign n3791 =  ( n3789 ) | ( n3790 )  ;
assign n3792 = ~ ( n2530 ) ;
assign n3793 =  ( n3791 ) | ( n3792 )  ;
assign n3794 = ~ ( n2573 ) ;
assign n3795 =  ( n3793 ) | ( n3794 )  ;
assign n3796 = ~ ( n2629 ) ;
assign n3797 =  ( n3795 ) | ( n3796 )  ;
assign n3798 = ~ ( n2698 ) ;
assign n3799 =  ( n3797 ) | ( n3798 )  ;
assign n3800 =  ( n2736 ) | ( n2769 )  ;
assign n3801 =  ( n3800 ) | ( n2858 )  ;
assign n3802 =  ( n3801 ) | ( n3028 )  ;
assign n3803 = ~ ( n3802 ) ;
assign n3804 =  ( n3799 ) | ( n3803 )  ;
assign n3805 = ~ ( n3804 ) ;
assign n3806 =  ( n3786 ) | ( n3805 )  ;
assign n3807 = ~ ( n2264 ) ;
assign n3808 = ~ ( n2404 ) ;
assign n3809 =  ( n3807 ) | ( n3808 )  ;
assign n3810 = ~ ( n2433 ) ;
assign n3811 =  ( n3809 ) | ( n3810 )  ;
assign n3812 = ~ ( n2530 ) ;
assign n3813 =  ( n3811 ) | ( n3812 )  ;
assign n3814 = ~ ( n2573 ) ;
assign n3815 =  ( n3813 ) | ( n3814 )  ;
assign n3816 = ~ ( n2629 ) ;
assign n3817 =  ( n3815 ) | ( n3816 )  ;
assign n3818 = ~ ( n2698 ) ;
assign n3819 =  ( n3817 ) | ( n3818 )  ;
assign n3820 = ~ ( n2749 ) ;
assign n3821 =  ( n3819 ) | ( n3820 )  ;
assign n3822 = ~ ( n2786 ) ;
assign n3823 =  ( n3821 ) | ( n3822 )  ;
assign n3824 = ~ ( n2834 ) ;
assign n3825 =  ( n3823 ) | ( n3824 )  ;
assign n3826 = ~ ( n2879 ) ;
assign n3827 =  ( n3825 ) | ( n3826 )  ;
assign n3828 = ~ ( n2926 ) ;
assign n3829 =  ( n3827 ) | ( n3828 )  ;
assign n3830 = ~ ( n2961 ) ;
assign n3831 =  ( n3829 ) | ( n3830 )  ;
assign n3832 = ~ ( n3003 ) ;
assign n3833 =  ( n3831 ) | ( n3832 )  ;
assign n3834 = ~ ( n3054 ) ;
assign n3835 =  ( n3833 ) | ( n3834 )  ;
assign n3836 =  ( n3075 ) | ( n3101 )  ;
assign n3837 =  ( n3836 ) | ( n3186 )  ;
assign n3838 = ~ ( n3262 ) ;
assign n3839 =  ( n3837 ) | ( n3838 )  ;
assign n3840 = ~ ( n3839 ) ;
assign n3841 =  ( n3835 ) | ( n3840 )  ;
assign n3842 = ~ ( n3841 ) ;
assign n3843 =  ( n3806 ) | ( n3842 )  ;
assign n3844 = ~ ( n3843 ) ;
assign n3845 =  ( n3776 ) | ( n3844 )  ;
assign n3846 = ~ ( n3845 ) ;
assign n3847 =  ( n3775 ) | ( n3846 )  ;
assign n3848 =  ( n3774 ) ^ ( n3847 )  ;
assign n3849 =  { ( n3769 ) , ( n3848 ) }  ;
assign n3850 = ~ ( n2125 ) ;
assign n3851 = ~ ( n1531 ) ;
assign n3852 =  ( n3851 ) | ( n1546 )  ;
assign n3853 = ~ ( n3852 ) ;
assign n3854 =  ( n3850 ) ^ ( n3853 )  ;
assign n3855 =  ( n3854 ) ^ ( n3843 )  ;
assign n3856 =  { ( n3849 ) , ( n3855 ) }  ;
assign n3857 = ~ ( n2259 ) ;
assign n3858 = ~ ( n1531 ) ;
assign n3859 =  ( n3858 ) | ( n1546 )  ;
assign n3860 = ~ ( n3859 ) ;
assign n3861 =  ( n3857 ) ^ ( n3860 )  ;
assign n3862 = ~ ( n2245 ) ;
assign n3863 = ~ ( n2264 ) ;
assign n3864 = ~ ( n1531 ) ;
assign n3865 =  ( n2393 ) | ( n3864 )  ;
assign n3866 =  ( n3865 ) | ( n1546 )  ;
assign n3867 = ~ ( n3866 ) ;
assign n3868 = ~ ( n2404 ) ;
assign n3869 =  ( n3868 ) | ( n2411 )  ;
assign n3870 = ~ ( n1531 ) ;
assign n3871 =  ( n3869 ) | ( n3870 )  ;
assign n3872 =  ( n3871 ) | ( n1546 )  ;
assign n3873 = ~ ( n3872 ) ;
assign n3874 =  ( n3867 ) | ( n3873 )  ;
assign n3875 = ~ ( n3334 ) ;
assign n3876 =  ( n3874 ) | ( n3875 )  ;
assign n3877 =  ( n3876 ) | ( n3355 )  ;
assign n3878 = ~ ( n2404 ) ;
assign n3879 = ~ ( n2433 ) ;
assign n3880 =  ( n3878 ) | ( n3879 )  ;
assign n3881 = ~ ( n2530 ) ;
assign n3882 =  ( n3880 ) | ( n3881 )  ;
assign n3883 = ~ ( n2573 ) ;
assign n3884 =  ( n3882 ) | ( n3883 )  ;
assign n3885 = ~ ( n2629 ) ;
assign n3886 =  ( n3884 ) | ( n3885 )  ;
assign n3887 = ~ ( n2698 ) ;
assign n3888 =  ( n3886 ) | ( n3887 )  ;
assign n3889 = ~ ( n2749 ) ;
assign n3890 =  ( n3888 ) | ( n3889 )  ;
assign n3891 = ~ ( n2786 ) ;
assign n3892 =  ( n3890 ) | ( n3891 )  ;
assign n3893 =  ( n2822 ) | ( n2854 )  ;
assign n3894 =  ( n3893 ) | ( n3391 )  ;
assign n3895 =  ( n3894 ) | ( n3411 )  ;
assign n3896 = ~ ( n3895 ) ;
assign n3897 =  ( n3892 ) | ( n3896 )  ;
assign n3898 = ~ ( n3897 ) ;
assign n3899 =  ( n3877 ) | ( n3898 )  ;
assign n3900 = ~ ( n2404 ) ;
assign n3901 = ~ ( n2433 ) ;
assign n3902 =  ( n3900 ) | ( n3901 )  ;
assign n3903 = ~ ( n2530 ) ;
assign n3904 =  ( n3902 ) | ( n3903 )  ;
assign n3905 = ~ ( n2573 ) ;
assign n3906 =  ( n3904 ) | ( n3905 )  ;
assign n3907 = ~ ( n2629 ) ;
assign n3908 =  ( n3906 ) | ( n3907 )  ;
assign n3909 = ~ ( n2698 ) ;
assign n3910 =  ( n3908 ) | ( n3909 )  ;
assign n3911 = ~ ( n2749 ) ;
assign n3912 =  ( n3910 ) | ( n3911 )  ;
assign n3913 = ~ ( n2786 ) ;
assign n3914 =  ( n3912 ) | ( n3913 )  ;
assign n3915 = ~ ( n2834 ) ;
assign n3916 =  ( n3914 ) | ( n3915 )  ;
assign n3917 = ~ ( n2879 ) ;
assign n3918 =  ( n3916 ) | ( n3917 )  ;
assign n3919 = ~ ( n2926 ) ;
assign n3920 =  ( n3918 ) | ( n3919 )  ;
assign n3921 = ~ ( n2961 ) ;
assign n3922 =  ( n3920 ) | ( n3921 )  ;
assign n3923 = ~ ( n3003 ) ;
assign n3924 =  ( n3922 ) | ( n3923 )  ;
assign n3925 = ~ ( n3054 ) ;
assign n3926 =  ( n3924 ) | ( n3925 )  ;
assign n3927 = ~ ( n3085 ) ;
assign n3928 =  ( n3926 ) | ( n3927 )  ;
assign n3929 = ~ ( n3114 ) ;
assign n3930 =  ( n3928 ) | ( n3929 )  ;
assign n3931 =  ( n3148 ) | ( n3182 )  ;
assign n3932 =  ( n3931 ) | ( n3435 )  ;
assign n3933 = ~ ( n3458 ) ;
assign n3934 =  ( n3932 ) | ( n3933 )  ;
assign n3935 = ~ ( n3934 ) ;
assign n3936 =  ( n3930 ) | ( n3935 )  ;
assign n3937 = ~ ( n3936 ) ;
assign n3938 =  ( n3899 ) | ( n3937 )  ;
assign n3939 = ~ ( n3938 ) ;
assign n3940 =  ( n3863 ) | ( n3939 )  ;
assign n3941 = ~ ( n3940 ) ;
assign n3942 =  ( n3862 ) | ( n3941 )  ;
assign n3943 =  ( n3861 ) ^ ( n3942 )  ;
assign n3944 =  { ( n3856 ) , ( n3943 ) }  ;
assign n3945 = ~ ( n2259 ) ;
assign n3946 = ~ ( n1531 ) ;
assign n3947 =  ( n3946 ) | ( n1546 )  ;
assign n3948 = ~ ( n3947 ) ;
assign n3949 =  ( n3945 ) ^ ( n3948 )  ;
assign n3950 =  ( n3949 ) ^ ( n3938 )  ;
assign n3951 =  { ( n3944 ) , ( n3950 ) }  ;
assign n3952 = ~ ( n118 ) ;
assign n3953 =  ( n3952 ) | ( n110 )  ;
assign n3954 =  ( n3953 ) ^ ( n2391 )  ;
assign n3955 = ~ ( n1531 ) ;
assign n3956 =  ( n3955 ) | ( n1546 )  ;
assign n3957 = ~ ( n3956 ) ;
assign n3958 =  ( n3954 ) ^ ( n3957 )  ;
assign n3959 = ~ ( n1531 ) ;
assign n3960 =  ( n2411 ) | ( n3959 )  ;
assign n3961 =  ( n3960 ) | ( n1546 )  ;
assign n3962 = ~ ( n3961 ) ;
assign n3963 = ~ ( n2433 ) ;
assign n3964 = ~ ( n2518 ) ;
assign n3965 =  ( n3964 ) | ( n2553 )  ;
assign n3966 =  ( n3965 ) | ( n2654 )  ;
assign n3967 =  ( n3966 ) | ( n3532 )  ;
assign n3968 = ~ ( n2530 ) ;
assign n3969 = ~ ( n2573 ) ;
assign n3970 =  ( n3968 ) | ( n3969 )  ;
assign n3971 = ~ ( n2629 ) ;
assign n3972 =  ( n3970 ) | ( n3971 )  ;
assign n3973 = ~ ( n2698 ) ;
assign n3974 =  ( n3972 ) | ( n3973 )  ;
assign n3975 = ~ ( n2749 ) ;
assign n3976 =  ( n3974 ) | ( n3975 )  ;
assign n3977 = ~ ( n2786 ) ;
assign n3978 =  ( n3976 ) | ( n3977 )  ;
assign n3979 = ~ ( n2834 ) ;
assign n3980 =  ( n3978 ) | ( n3979 )  ;
assign n3981 = ~ ( n2879 ) ;
assign n3982 =  ( n3980 ) | ( n3981 )  ;
assign n3983 =  ( n2914 ) | ( n2945 )  ;
assign n3984 =  ( n3983 ) | ( n3024 )  ;
assign n3985 =  ( n3984 ) | ( n3576 )  ;
assign n3986 = ~ ( n3985 ) ;
assign n3987 =  ( n3982 ) | ( n3986 )  ;
assign n3988 = ~ ( n3987 ) ;
assign n3989 =  ( n3967 ) | ( n3988 )  ;
assign n3990 = ~ ( n2530 ) ;
assign n3991 = ~ ( n2573 ) ;
assign n3992 =  ( n3990 ) | ( n3991 )  ;
assign n3993 = ~ ( n2629 ) ;
assign n3994 =  ( n3992 ) | ( n3993 )  ;
assign n3995 = ~ ( n2698 ) ;
assign n3996 =  ( n3994 ) | ( n3995 )  ;
assign n3997 = ~ ( n2749 ) ;
assign n3998 =  ( n3996 ) | ( n3997 )  ;
assign n3999 = ~ ( n2786 ) ;
assign n4000 =  ( n3998 ) | ( n3999 )  ;
assign n4001 = ~ ( n2834 ) ;
assign n4002 =  ( n4000 ) | ( n4001 )  ;
assign n4003 = ~ ( n2879 ) ;
assign n4004 =  ( n4002 ) | ( n4003 )  ;
assign n4005 = ~ ( n2926 ) ;
assign n4006 =  ( n4004 ) | ( n4005 )  ;
assign n4007 = ~ ( n2961 ) ;
assign n4008 =  ( n4006 ) | ( n4007 )  ;
assign n4009 = ~ ( n3003 ) ;
assign n4010 =  ( n4008 ) | ( n4009 )  ;
assign n4011 = ~ ( n3054 ) ;
assign n4012 =  ( n4010 ) | ( n4011 )  ;
assign n4013 = ~ ( n3085 ) ;
assign n4014 =  ( n4012 ) | ( n4013 )  ;
assign n4015 = ~ ( n3114 ) ;
assign n4016 =  ( n4014 ) | ( n4015 )  ;
assign n4017 = ~ ( n3158 ) ;
assign n4018 =  ( n4016 ) | ( n4017 )  ;
assign n4019 = ~ ( n3201 ) ;
assign n4020 =  ( n4018 ) | ( n4019 )  ;
assign n4021 =  ( n3217 ) | ( n3239 )  ;
assign n4022 = ~ ( n3258 ) ;
assign n4023 =  ( n4021 ) | ( n4022 )  ;
assign n4024 = ~ ( n4023 ) ;
assign n4025 =  ( n4020 ) | ( n4024 )  ;
assign n4026 = ~ ( n4025 ) ;
assign n4027 =  ( n3989 ) | ( n4026 )  ;
assign n4028 = ~ ( n4027 ) ;
assign n4029 =  ( n3963 ) | ( n4028 )  ;
assign n4030 = ~ ( n4029 ) ;
assign n4031 =  ( n3962 ) | ( n4030 )  ;
assign n4032 =  ( n3958 ) ^ ( n4031 )  ;
assign n4033 =  { ( n3951 ) , ( n4032 ) }  ;
assign n4034 = ~ ( n195 ) ;
assign n4035 = ~ ( n118 ) ;
assign n4036 =  ( n4035 ) | ( n110 )  ;
assign n4037 =  ( n4034 ) ^ ( n4036 )  ;
assign n4038 =  ( n4037 ) ^ ( n2387 )  ;
assign n4039 = ~ ( n1531 ) ;
assign n4040 =  ( n4039 ) | ( n1546 )  ;
assign n4041 = ~ ( n4040 ) ;
assign n4042 =  ( n4038 ) ^ ( n4041 )  ;
assign n4043 = ~ ( n2518 ) ;
assign n4044 =  ( n4043 ) | ( n2553 )  ;
assign n4045 =  ( n4044 ) | ( n2654 )  ;
assign n4046 =  ( n4045 ) | ( n3532 )  ;
assign n4047 =  ( n4046 ) | ( n3988 )  ;
assign n4048 = ~ ( n4025 ) ;
assign n4049 =  ( n4047 ) | ( n4048 )  ;
assign n4050 =  ( n4042 ) ^ ( n4049 )  ;
assign n4051 =  { ( n4033 ) , ( n4050 ) }  ;
assign n4052 = ~ ( n286 ) ;
assign n4053 =  ( n304 ) ^ ( n4052 )  ;
assign n4054 =  ( n4053 ) ^ ( n118 )  ;
assign n4055 = ~ ( n110 ) ;
assign n4056 =  ( n4054 ) ^ ( n4055 )  ;
assign n4057 =  ( n2445 ) | ( n2512 )  ;
assign n4058 =  ( n4056 ) ^ ( n4057 )  ;
assign n4059 = ~ ( n1531 ) ;
assign n4060 =  ( n4059 ) | ( n1546 )  ;
assign n4061 = ~ ( n4060 ) ;
assign n4062 =  ( n4058 ) ^ ( n4061 )  ;
assign n4063 = ~ ( n2547 ) ;
assign n4064 =  ( n1531 ) ^ ( n1546 )  ;
assign n4065 = ~ ( n4064 ) ;
assign n4066 =  ( n4063 ) | ( n4065 )  ;
assign n4067 = ~ ( n4066 ) ;
assign n4068 = ~ ( n2573 ) ;
assign n4069 =  ( n2614 ) | ( n2650 )  ;
assign n4070 =  ( n4069 ) | ( n3351 )  ;
assign n4071 =  ( n4070 ) | ( n3673 )  ;
assign n4072 = ~ ( n2629 ) ;
assign n4073 = ~ ( n2698 ) ;
assign n4074 =  ( n4072 ) | ( n4073 )  ;
assign n4075 = ~ ( n2749 ) ;
assign n4076 =  ( n4074 ) | ( n4075 )  ;
assign n4077 = ~ ( n2786 ) ;
assign n4078 =  ( n4076 ) | ( n4077 )  ;
assign n4079 = ~ ( n2834 ) ;
assign n4080 =  ( n4078 ) | ( n4079 )  ;
assign n4081 = ~ ( n2879 ) ;
assign n4082 =  ( n4080 ) | ( n4081 )  ;
assign n4083 = ~ ( n2926 ) ;
assign n4084 =  ( n4082 ) | ( n4083 )  ;
assign n4085 = ~ ( n2961 ) ;
assign n4086 =  ( n4084 ) | ( n4085 )  ;
assign n4087 =  ( n2992 ) | ( n3020 )  ;
assign n4088 =  ( n4087 ) | ( n3407 )  ;
assign n4089 =  ( n4088 ) | ( n3719 )  ;
assign n4090 = ~ ( n4089 ) ;
assign n4091 =  ( n4086 ) | ( n4090 )  ;
assign n4092 = ~ ( n4091 ) ;
assign n4093 =  ( n4071 ) | ( n4092 )  ;
assign n4094 = ~ ( n2629 ) ;
assign n4095 = ~ ( n2698 ) ;
assign n4096 =  ( n4094 ) | ( n4095 )  ;
assign n4097 = ~ ( n2749 ) ;
assign n4098 =  ( n4096 ) | ( n4097 )  ;
assign n4099 = ~ ( n2786 ) ;
assign n4100 =  ( n4098 ) | ( n4099 )  ;
assign n4101 = ~ ( n2834 ) ;
assign n4102 =  ( n4100 ) | ( n4101 )  ;
assign n4103 = ~ ( n2879 ) ;
assign n4104 =  ( n4102 ) | ( n4103 )  ;
assign n4105 = ~ ( n2926 ) ;
assign n4106 =  ( n4104 ) | ( n4105 )  ;
assign n4107 = ~ ( n2961 ) ;
assign n4108 =  ( n4106 ) | ( n4107 )  ;
assign n4109 = ~ ( n3003 ) ;
assign n4110 =  ( n4108 ) | ( n4109 )  ;
assign n4111 = ~ ( n3054 ) ;
assign n4112 =  ( n4110 ) | ( n4111 )  ;
assign n4113 = ~ ( n3085 ) ;
assign n4114 =  ( n4112 ) | ( n4113 )  ;
assign n4115 = ~ ( n3114 ) ;
assign n4116 =  ( n4114 ) | ( n4115 )  ;
assign n4117 = ~ ( n3158 ) ;
assign n4118 =  ( n4116 ) | ( n4117 )  ;
assign n4119 = ~ ( n3201 ) ;
assign n4120 =  ( n4118 ) | ( n4119 )  ;
assign n4121 =  ( n1434 ) ^ ( n1444 )  ;
assign n4122 =  ( n4121 ) ^ ( n3211 )  ;
assign n4123 =  ( n4122 ) ^ ( n1531 )  ;
assign n4124 =  ( n4123 ) ^ ( n1546 )  ;
assign n4125 = ~ ( n4124 ) ;
assign n4126 =  ( n4120 ) | ( n4125 )  ;
assign n4127 =  ( n1497 ) ^ ( n3227 )  ;
assign n4128 =  ( n4127 ) ^ ( n1531 )  ;
assign n4129 =  ( n4128 ) ^ ( n3235 )  ;
assign n4130 = ~ ( n4129 ) ;
assign n4131 =  ( n4126 ) | ( n4130 )  ;
assign n4132 = ki[1:1] ;
assign n4133 =  ( n1506 ) ^ ( n4132 )  ;
assign n4134 = ~ ( n4133 ) ;
assign n4135 =  ( n4131 ) | ( n4134 )  ;
assign n4136 = kd[1:1] ;
assign n4137 =  ( n1540 ) ^ ( n4136 )  ;
assign n4138 = ~ ( n4137 ) ;
assign n4139 =  ( n4135 ) | ( n4138 )  ;
assign n4140 = ~ ( n4139 ) ;
assign n4141 =  ( n4093 ) | ( n4140 )  ;
assign n4142 = ~ ( n4141 ) ;
assign n4143 =  ( n4068 ) | ( n4142 )  ;
assign n4144 = ~ ( n4143 ) ;
assign n4145 =  ( n4067 ) | ( n4144 )  ;
assign n4146 =  ( n4062 ) ^ ( n4145 )  ;
assign n4147 =  { ( n4051 ) , ( n4146 ) }  ;
assign n4148 =  ( n376 ) | ( n394 )  ;
assign n4149 =  ( bv_1_1_n2 ) ^ ( n4148 )  ;
assign n4150 =  ( n4149 ) ^ ( n406 )  ;
assign n4151 = ~ ( n268 ) ;
assign n4152 =  ( n4150 ) ^ ( n4151 )  ;
assign n4153 = ~ ( n100 ) ;
assign n4154 =  ( n75 ) | ( n4153 )  ;
assign n4155 = ~ ( n4154 ) ;
assign n4156 =  ( n4152 ) ^ ( n4155 )  ;
assign n4157 =  ( n4156 ) ^ ( n110 )  ;
assign n4158 =  ( n524 ) | ( n632 )  ;
assign n4159 =  ( n4158 ) | ( n1586 )  ;
assign n4160 =  ( n4159 ) | ( n1927 )  ;
assign n4161 =  ( n4160 ) | ( n2469 )  ;
assign n4162 =  ( n4161 ) | ( n2508 )  ;
assign n4163 =  ( n4157 ) ^ ( n4162 )  ;
assign n4164 =  ( n4163 ) ^ ( n1531 )  ;
assign n4165 =  ( n4164 ) ^ ( n1546 )  ;
assign n4166 =  ( n2614 ) | ( n2650 )  ;
assign n4167 =  ( n4166 ) | ( n3351 )  ;
assign n4168 =  ( n4167 ) | ( n3673 )  ;
assign n4169 =  ( n4168 ) | ( n4092 )  ;
assign n4170 = ~ ( n4139 ) ;
assign n4171 =  ( n4169 ) | ( n4170 )  ;
assign n4172 =  ( n4165 ) ^ ( n4171 )  ;
assign n4173 =  { ( n4147 ) , ( n4172 ) }  ;
assign n4174 =  ( bv_1_1_n2 ) ^ ( n535 )  ;
assign n4175 =  ( n4174 ) ^ ( n385 )  ;
assign n4176 =  ( n4175 ) ^ ( n365 )  ;
assign n4177 = ~ ( n150 ) ;
assign n4178 = ~ ( n160 ) ;
assign n4179 =  ( n4177 ) | ( n4178 )  ;
assign n4180 = ~ ( n4179 ) ;
assign n4181 =  ( n4176 ) ^ ( n4180 )  ;
assign n4182 = ~ ( n75 ) ;
assign n4183 =  ( n4181 ) ^ ( n4182 )  ;
assign n4184 =  ( n4183 ) ^ ( n100 )  ;
assign n4185 =  ( n2599 ) | ( n2607 )  ;
assign n4186 =  ( n4184 ) ^ ( n4185 )  ;
assign n4187 =  ( n4186 ) ^ ( n1531 )  ;
assign n4188 =  ( n4187 ) ^ ( n1546 )  ;
assign n4189 = ~ ( n2644 ) ;
assign n4190 =  ( n1531 ) ^ ( n1546 )  ;
assign n4191 = ~ ( n4190 ) ;
assign n4192 =  ( n4189 ) | ( n4191 )  ;
assign n4193 = ~ ( n4192 ) ;
assign n4194 = ~ ( n2698 ) ;
assign n4195 =  ( n2736 ) | ( n2769 )  ;
assign n4196 =  ( n4195 ) | ( n2858 )  ;
assign n4197 =  ( n4196 ) | ( n3028 )  ;
assign n4198 = ~ ( n3266 ) ;
assign n4199 =  ( n4197 ) | ( n4198 )  ;
assign n4200 = ~ ( n4199 ) ;
assign n4201 =  ( n4194 ) | ( n4200 )  ;
assign n4202 = ~ ( n4201 ) ;
assign n4203 =  ( n4193 ) | ( n4202 )  ;
assign n4204 =  ( n4188 ) ^ ( n4203 )  ;
assign n4205 =  { ( n4173 ) , ( n4204 ) }  ;
assign n4206 =  ( n667 ) ^ ( n621 )  ;
assign n4207 =  ( n4206 ) ^ ( n502 )  ;
assign n4208 = ~ ( n227 ) ;
assign n4209 = ~ ( n247 ) ;
assign n4210 =  ( n4208 ) | ( n4209 )  ;
assign n4211 = ~ ( n4210 ) ;
assign n4212 =  ( n4207 ) ^ ( n4211 )  ;
assign n4213 =  ( n4212 ) ^ ( n150 )  ;
assign n4214 =  ( n4213 ) ^ ( n160 )  ;
assign n4215 =  ( n766 ) | ( n872 )  ;
assign n4216 =  ( n4215 ) | ( n985 )  ;
assign n4217 =  ( n4216 ) | ( n1254 )  ;
assign n4218 =  ( n4217 ) | ( n1516 )  ;
assign n4219 =  ( n4214 ) ^ ( n4218 )  ;
assign n4220 =  ( n4219 ) ^ ( n1531 )  ;
assign n4221 =  ( n4220 ) ^ ( n1546 )  ;
assign n4222 =  ( n2736 ) | ( n2769 )  ;
assign n4223 =  ( n4222 ) | ( n2858 )  ;
assign n4224 =  ( n4223 ) | ( n3028 )  ;
assign n4225 = ~ ( n3266 ) ;
assign n4226 =  ( n4224 ) | ( n4225 )  ;
assign n4227 =  ( n4221 ) ^ ( n4226 )  ;
assign n4228 =  { ( n4205 ) , ( n4227 ) }  ;
assign n4229 =  ( n777 ) ^ ( n755 )  ;
assign n4230 =  ( n4229 ) ^ ( n603 )  ;
assign n4231 = ~ ( n336 ) ;
assign n4232 = ~ ( n345 ) ;
assign n4233 =  ( n4231 ) | ( n4232 )  ;
assign n4234 = ~ ( n4233 ) ;
assign n4235 =  ( n4230 ) ^ ( n4234 )  ;
assign n4236 =  ( n4235 ) ^ ( n227 )  ;
assign n4237 =  ( n4236 ) ^ ( n247 )  ;
assign n4238 =  ( n2722 ) | ( n2729 )  ;
assign n4239 =  ( n4237 ) ^ ( n4238 )  ;
assign n4240 =  ( n4239 ) ^ ( n1531 )  ;
assign n4241 =  ( n4240 ) ^ ( n1546 )  ;
assign n4242 = ~ ( n2763 ) ;
assign n4243 =  ( n1531 ) ^ ( n1546 )  ;
assign n4244 = ~ ( n4243 ) ;
assign n4245 =  ( n4242 ) | ( n4244 )  ;
assign n4246 = ~ ( n4245 ) ;
assign n4247 = ~ ( n2786 ) ;
assign n4248 =  ( n2822 ) | ( n2854 )  ;
assign n4249 =  ( n4248 ) | ( n3391 )  ;
assign n4250 =  ( n4249 ) | ( n3411 )  ;
assign n4251 = ~ ( n3462 ) ;
assign n4252 =  ( n4250 ) | ( n4251 )  ;
assign n4253 = ~ ( n4252 ) ;
assign n4254 =  ( n4247 ) | ( n4253 )  ;
assign n4255 = ~ ( n4254 ) ;
assign n4256 =  ( n4246 ) | ( n4255 )  ;
assign n4257 =  ( n4241 ) ^ ( n4256 )  ;
assign n4258 =  { ( n4228 ) , ( n4257 ) }  ;
assign n4259 =  ( n885 ) ^ ( n861 )  ;
assign n4260 =  ( n4259 ) ^ ( n737 )  ;
assign n4261 = ~ ( n462 ) ;
assign n4262 = ~ ( n482 ) ;
assign n4263 =  ( n4261 ) | ( n4262 )  ;
assign n4264 = ~ ( n4263 ) ;
assign n4265 =  ( n4260 ) ^ ( n4264 )  ;
assign n4266 =  ( n4265 ) ^ ( n336 )  ;
assign n4267 =  ( n4266 ) ^ ( n345 )  ;
assign n4268 =  ( n1625 ) | ( n1632 )  ;
assign n4269 =  ( n4268 ) | ( n1668 )  ;
assign n4270 =  ( n4269 ) | ( n1703 )  ;
assign n4271 =  ( n4267 ) ^ ( n4270 )  ;
assign n4272 =  ( n4271 ) ^ ( n1531 )  ;
assign n4273 =  ( n4272 ) ^ ( n1546 )  ;
assign n4274 =  ( n2822 ) | ( n2854 )  ;
assign n4275 =  ( n4274 ) | ( n3391 )  ;
assign n4276 =  ( n4275 ) | ( n3411 )  ;
assign n4277 = ~ ( n3462 ) ;
assign n4278 =  ( n4276 ) | ( n4277 )  ;
assign n4279 =  ( n4273 ) ^ ( n4278 )  ;
assign n4280 =  { ( n4258 ) , ( n4279 ) }  ;
assign n4281 =  ( n905 ) ^ ( n843 )  ;
assign n4282 = ~ ( n573 ) ;
assign n4283 = ~ ( n583 ) ;
assign n4284 =  ( n4282 ) | ( n4283 )  ;
assign n4285 = ~ ( n4284 ) ;
assign n4286 =  ( n4281 ) ^ ( n4285 )  ;
assign n4287 =  ( n4286 ) ^ ( n462 )  ;
assign n4288 =  ( n4287 ) ^ ( n482 )  ;
assign n4289 =  ( n2807 ) | ( n2815 )  ;
assign n4290 =  ( n4288 ) ^ ( n4289 )  ;
assign n4291 =  ( n4290 ) ^ ( n1531 )  ;
assign n4292 =  ( n4291 ) ^ ( n1546 )  ;
assign n4293 = ~ ( n2848 ) ;
assign n4294 =  ( n1531 ) ^ ( n1546 )  ;
assign n4295 = ~ ( n4294 ) ;
assign n4296 =  ( n4293 ) | ( n4295 )  ;
assign n4297 = ~ ( n4296 ) ;
assign n4298 = ~ ( n2879 ) ;
assign n4299 =  ( n2914 ) | ( n2945 )  ;
assign n4300 =  ( n4299 ) | ( n3024 )  ;
assign n4301 =  ( n4300 ) | ( n3576 )  ;
assign n4302 = ~ ( n3597 ) ;
assign n4303 =  ( n4301 ) | ( n4302 )  ;
assign n4304 = ~ ( n4303 ) ;
assign n4305 =  ( n4298 ) | ( n4304 )  ;
assign n4306 = ~ ( n4305 ) ;
assign n4307 =  ( n4297 ) | ( n4306 )  ;
assign n4308 =  ( n4292 ) ^ ( n4307 )  ;
assign n4309 =  { ( n4280 ) , ( n4308 ) }  ;
assign n4310 =  ( n1000 ) ^ ( n975 )  ;
assign n4311 = ~ ( n704 ) ;
assign n4312 = ~ ( n717 ) ;
assign n4313 =  ( n4311 ) | ( n4312 )  ;
assign n4314 = ~ ( n4313 ) ;
assign n4315 =  ( n4310 ) ^ ( n4314 )  ;
assign n4316 =  ( n4315 ) ^ ( n573 )  ;
assign n4317 =  ( n4316 ) ^ ( n583 )  ;
assign n4318 =  ( n1075 ) | ( n1163 )  ;
assign n4319 =  ( n4318 ) | ( n1250 )  ;
assign n4320 =  ( n4319 ) | ( n1821 )  ;
assign n4321 =  ( n4320 ) | ( n1848 )  ;
assign n4322 =  ( n4317 ) ^ ( n4321 )  ;
assign n4323 =  ( n4322 ) ^ ( n1531 )  ;
assign n4324 =  ( n4323 ) ^ ( n1546 )  ;
assign n4325 =  ( n2914 ) | ( n2945 )  ;
assign n4326 =  ( n4325 ) | ( n3024 )  ;
assign n4327 =  ( n4326 ) | ( n3576 )  ;
assign n4328 = ~ ( n3597 ) ;
assign n4329 =  ( n4327 ) | ( n4328 )  ;
assign n4330 =  ( n4324 ) ^ ( n4329 )  ;
assign n4331 =  { ( n4309 ) , ( n4330 ) }  ;
assign n4332 =  ( n1084 ) ^ ( n1065 )  ;
assign n4333 = ~ ( n813 ) ;
assign n4334 = ~ ( n823 ) ;
assign n4335 =  ( n4333 ) | ( n4334 )  ;
assign n4336 = ~ ( n4335 ) ;
assign n4337 =  ( n4332 ) ^ ( n4336 )  ;
assign n4338 =  ( n4337 ) ^ ( n704 )  ;
assign n4339 =  ( n4338 ) ^ ( n717 )  ;
assign n4340 =  ( n2900 ) | ( n2907 )  ;
assign n4341 =  ( n4339 ) ^ ( n4340 )  ;
assign n4342 =  ( n4341 ) ^ ( n1531 )  ;
assign n4343 =  ( n4342 ) ^ ( n1546 )  ;
assign n4344 = ~ ( n2939 ) ;
assign n4345 =  ( n1531 ) ^ ( n1546 )  ;
assign n4346 = ~ ( n4345 ) ;
assign n4347 =  ( n4344 ) | ( n4346 )  ;
assign n4348 = ~ ( n4347 ) ;
assign n4349 = ~ ( n2961 ) ;
assign n4350 =  ( n2992 ) | ( n3020 )  ;
assign n4351 =  ( n4350 ) | ( n3407 )  ;
assign n4352 =  ( n4351 ) | ( n3719 )  ;
assign n4353 = ~ ( n3750 ) ;
assign n4354 =  ( n4352 ) | ( n4353 )  ;
assign n4355 = ~ ( n4354 ) ;
assign n4356 =  ( n4349 ) | ( n4355 )  ;
assign n4357 = ~ ( n4356 ) ;
assign n4358 =  ( n4348 ) | ( n4357 )  ;
assign n4359 =  ( n4343 ) ^ ( n4358 )  ;
assign n4360 =  { ( n4331 ) , ( n4359 ) }  ;
assign n4361 =  ( n1174 ) ^ ( n1153 )  ;
assign n4362 = ~ ( n941 ) ;
assign n4363 = ~ ( n955 ) ;
assign n4364 =  ( n4362 ) | ( n4363 )  ;
assign n4365 = ~ ( n4364 ) ;
assign n4366 =  ( n4361 ) ^ ( n4365 )  ;
assign n4367 =  ( n4366 ) ^ ( n813 )  ;
assign n4368 =  ( n4367 ) ^ ( n823 )  ;
assign n4369 =  ( n1651 ) | ( n1664 )  ;
assign n4370 =  ( n4369 ) | ( n1973 )  ;
assign n4371 =  ( n4370 ) | ( n1996 )  ;
assign n4372 =  ( n4368 ) ^ ( n4371 )  ;
assign n4373 =  ( n4372 ) ^ ( n1531 )  ;
assign n4374 =  ( n4373 ) ^ ( n1546 )  ;
assign n4375 =  ( n2992 ) | ( n3020 )  ;
assign n4376 =  ( n4375 ) | ( n3407 )  ;
assign n4377 =  ( n4376 ) | ( n3719 )  ;
assign n4378 = ~ ( n3750 ) ;
assign n4379 =  ( n4377 ) | ( n4378 )  ;
assign n4380 =  ( n4374 ) ^ ( n4379 )  ;
assign n4381 =  { ( n4360 ) , ( n4380 ) }  ;
assign n4382 = ~ ( n1036 ) ;
assign n4383 = ~ ( n1045 ) ;
assign n4384 =  ( n4382 ) | ( n4383 )  ;
assign n4385 = ~ ( n4384 ) ;
assign n4386 =  ( n1191 ) ^ ( n4385 )  ;
assign n4387 =  ( n4386 ) ^ ( n941 )  ;
assign n4388 =  ( n4387 ) ^ ( n955 )  ;
assign n4389 =  ( n2979 ) | ( n2985 )  ;
assign n4390 =  ( n4388 ) ^ ( n4389 )  ;
assign n4391 =  ( n4390 ) ^ ( n1531 )  ;
assign n4392 =  ( n4391 ) ^ ( n1546 )  ;
assign n4393 = ~ ( n3014 ) ;
assign n4394 =  ( n1531 ) ^ ( n1546 )  ;
assign n4395 = ~ ( n4394 ) ;
assign n4396 =  ( n4393 ) | ( n4395 )  ;
assign n4397 = ~ ( n4396 ) ;
assign n4398 = ~ ( n3054 ) ;
assign n4399 =  ( n3075 ) | ( n3101 )  ;
assign n4400 =  ( n4399 ) | ( n3186 )  ;
assign n4401 = ~ ( n3262 ) ;
assign n4402 =  ( n4400 ) | ( n4401 )  ;
assign n4403 = ~ ( n4402 ) ;
assign n4404 =  ( n4398 ) | ( n4403 )  ;
assign n4405 = ~ ( n4404 ) ;
assign n4406 =  ( n4397 ) | ( n4405 )  ;
assign n4407 =  ( n4392 ) ^ ( n4406 )  ;
assign n4408 =  { ( n4381 ) , ( n4407 ) }  ;
assign n4409 = ~ ( n1119 ) ;
assign n4410 = ~ ( n1133 ) ;
assign n4411 =  ( n4409 ) | ( n4410 )  ;
assign n4412 = ~ ( n4411 ) ;
assign n4413 =  ( n1275 ) ^ ( n4412 )  ;
assign n4414 =  ( n4413 ) ^ ( n1036 )  ;
assign n4415 =  ( n4414 ) ^ ( n1045 )  ;
assign n4416 =  ( n1337 ) | ( n1454 )  ;
assign n4417 =  ( n4416 ) | ( n1512 )  ;
assign n4418 =  ( n4415 ) ^ ( n4417 )  ;
assign n4419 =  ( n4418 ) ^ ( n1531 )  ;
assign n4420 =  ( n4419 ) ^ ( n1546 )  ;
assign n4421 =  ( n3075 ) | ( n3101 )  ;
assign n4422 =  ( n4421 ) | ( n3186 )  ;
assign n4423 = ~ ( n3262 ) ;
assign n4424 =  ( n4422 ) | ( n4423 )  ;
assign n4425 =  ( n4420 ) ^ ( n4424 )  ;
assign n4426 =  { ( n4408 ) , ( n4425 ) }  ;
assign n4427 = ~ ( n1226 ) ;
assign n4428 = ~ ( n1236 ) ;
assign n4429 =  ( n4427 ) | ( n4428 )  ;
assign n4430 = ~ ( n4429 ) ;
assign n4431 =  ( n1344 ) ^ ( n4430 )  ;
assign n4432 =  ( n4431 ) ^ ( n1119 )  ;
assign n4433 =  ( n4432 ) ^ ( n1133 )  ;
assign n4434 =  ( n4433 ) ^ ( n3069 )  ;
assign n4435 =  ( n4434 ) ^ ( n1531 )  ;
assign n4436 =  ( n4435 ) ^ ( n1546 )  ;
assign n4437 = ~ ( n3095 ) ;
assign n4438 =  ( n1531 ) ^ ( n1546 )  ;
assign n4439 = ~ ( n4438 ) ;
assign n4440 =  ( n4437 ) | ( n4439 )  ;
assign n4441 = ~ ( n4440 ) ;
assign n4442 = ~ ( n3114 ) ;
assign n4443 =  ( n3148 ) | ( n3182 )  ;
assign n4444 =  ( n4443 ) | ( n3435 )  ;
assign n4445 = ~ ( n3458 ) ;
assign n4446 =  ( n4444 ) | ( n4445 )  ;
assign n4447 = ~ ( n4446 ) ;
assign n4448 =  ( n4442 ) | ( n4447 )  ;
assign n4449 = ~ ( n4448 ) ;
assign n4450 =  ( n4441 ) | ( n4449 )  ;
assign n4451 =  ( n4436 ) ^ ( n4450 )  ;
assign n4452 =  { ( n4426 ) , ( n4451 ) }  ;
assign n4453 = ~ ( n1310 ) ;
assign n4454 = ~ ( n1323 ) ;
assign n4455 =  ( n4453 ) | ( n4454 )  ;
assign n4456 = ~ ( n4455 ) ;
assign n4457 =  ( n4456 ) ^ ( n1226 )  ;
assign n4458 =  ( n4457 ) ^ ( n1236 )  ;
assign n4459 =  ( n1401 ) | ( n1450 )  ;
assign n4460 =  ( n4459 ) | ( n1699 )  ;
assign n4461 =  ( n4458 ) ^ ( n4460 )  ;
assign n4462 =  ( n4461 ) ^ ( n1531 )  ;
assign n4463 =  ( n4462 ) ^ ( n1546 )  ;
assign n4464 =  ( n3148 ) | ( n3182 )  ;
assign n4465 =  ( n4464 ) | ( n3435 )  ;
assign n4466 = ~ ( n3458 ) ;
assign n4467 =  ( n4465 ) | ( n4466 )  ;
assign n4468 =  ( n4463 ) ^ ( n4467 )  ;
assign n4469 =  { ( n4452 ) , ( n4468 ) }  ;
assign n4470 = ~ ( n1386 ) ;
assign n4471 = ~ ( n1395 ) ;
assign n4472 =  ( n4470 ) | ( n4471 )  ;
assign n4473 = ~ ( n4472 ) ;
assign n4474 =  ( n4473 ) ^ ( n1310 )  ;
assign n4475 =  ( n4474 ) ^ ( n1323 )  ;
assign n4476 =  ( n3129 ) | ( n3141 )  ;
assign n4477 =  ( n4475 ) ^ ( n4476 )  ;
assign n4478 =  ( n4477 ) ^ ( n1531 )  ;
assign n4479 =  ( n4478 ) ^ ( n1546 )  ;
assign n4480 = ~ ( n3176 ) ;
assign n4481 =  ( n1531 ) ^ ( n1546 )  ;
assign n4482 = ~ ( n4481 ) ;
assign n4483 =  ( n4480 ) | ( n4482 )  ;
assign n4484 = ~ ( n4483 ) ;
assign n4485 = ~ ( n3201 ) ;
assign n4486 =  ( n3217 ) | ( n3239 )  ;
assign n4487 = ~ ( n3258 ) ;
assign n4488 =  ( n4486 ) | ( n4487 )  ;
assign n4489 = ~ ( n4488 ) ;
assign n4490 =  ( n4485 ) | ( n4489 )  ;
assign n4491 = ~ ( n4490 ) ;
assign n4492 =  ( n4484 ) | ( n4491 )  ;
assign n4493 =  ( n4479 ) ^ ( n4492 )  ;
assign n4494 =  { ( n4469 ) , ( n4493 ) }  ;
assign n4495 = ~ ( n1434 ) ;
assign n4496 = ~ ( n1444 ) ;
assign n4497 =  ( n4495 ) | ( n4496 )  ;
assign n4498 = ~ ( n4497 ) ;
assign n4499 =  ( n4498 ) ^ ( n1386 )  ;
assign n4500 =  ( n4499 ) ^ ( n1395 )  ;
assign n4501 =  ( n4500 ) ^ ( n3175 )  ;
assign n4502 =  ( n4501 ) ^ ( n1531 )  ;
assign n4503 =  ( n4502 ) ^ ( n1546 )  ;
assign n4504 =  ( n3217 ) | ( n3239 )  ;
assign n4505 = ~ ( n3258 ) ;
assign n4506 =  ( n4504 ) | ( n4505 )  ;
assign n4507 =  ( n4503 ) ^ ( n4506 )  ;
assign n4508 =  { ( n4494 ) , ( n4507 ) }  ;
assign n4509 =  ( n1434 ) ^ ( n1444 )  ;
assign n4510 =  ( n4509 ) ^ ( n3211 )  ;
assign n4511 =  ( n4510 ) ^ ( n1531 )  ;
assign n4512 =  ( n4511 ) ^ ( n1546 )  ;
assign n4513 =  ( n1497 ) ^ ( n3227 )  ;
assign n4514 = ~ ( n4513 ) ;
assign n4515 =  ( n1531 ) ^ ( n3235 )  ;
assign n4516 = ~ ( n4515 ) ;
assign n4517 =  ( n4514 ) | ( n4516 )  ;
assign n4518 = ~ ( n4517 ) ;
assign n4519 =  ( n1497 ) ^ ( n3227 )  ;
assign n4520 =  ( n4519 ) ^ ( n1531 )  ;
assign n4521 =  ( n4520 ) ^ ( n3235 )  ;
assign n4522 = ~ ( n4521 ) ;
assign n4523 = ki[1:1] ;
assign n4524 =  ( n1506 ) ^ ( n4523 )  ;
assign n4525 = ~ ( n4524 ) ;
assign n4526 =  ( n4522 ) | ( n4525 )  ;
assign n4527 = kd[1:1] ;
assign n4528 =  ( n1540 ) ^ ( n4527 )  ;
assign n4529 = ~ ( n4528 ) ;
assign n4530 =  ( n4526 ) | ( n4529 )  ;
assign n4531 = ~ ( n4530 ) ;
assign n4532 =  ( n4518 ) | ( n4531 )  ;
assign n4533 =  ( n4512 ) ^ ( n4532 )  ;
assign n4534 =  { ( n4508 ) , ( n4533 ) }  ;
assign n4535 =  ( n1497 ) ^ ( n3227 )  ;
assign n4536 =  ( n4535 ) ^ ( n1531 )  ;
assign n4537 =  ( n4536 ) ^ ( n3235 )  ;
assign n4538 = ki[1:1] ;
assign n4539 =  ( n1506 ) ^ ( n4538 )  ;
assign n4540 = ~ ( n4539 ) ;
assign n4541 = kd[1:1] ;
assign n4542 =  ( n1540 ) ^ ( n4541 )  ;
assign n4543 = ~ ( n4542 ) ;
assign n4544 =  ( n4540 ) | ( n4543 )  ;
assign n4545 = ~ ( n4544 ) ;
assign n4546 =  ( n4537 ) ^ ( n4545 )  ;
assign n4547 =  { ( n4534 ) , ( n4546 ) }  ;
assign n4548 = ki[1:1] ;
assign n4549 =  ( n1506 ) ^ ( n4548 )  ;
assign n4550 =  ( n4549 ) ^ ( n1540 )  ;
assign n4551 = kd[1:1] ;
assign n4552 =  ( n4550 ) ^ ( n4551 )  ;
assign n4553 =  { ( n4547 ) , ( n4552 ) }  ;
always @(posedge clk) begin
   if(rst) begin
       __COUNTER_start__n0 <= 0;
   end
   else if(__ILA_bar_valid__) begin
       if ( __ILA_bar_decode_of_i1__ ) begin 
           __COUNTER_start__n0 <= 1; end
       else if( (__COUNTER_start__n0 >= 1 ) && ( __COUNTER_start__n0 < 255 )) begin
           __COUNTER_start__n0 <= __COUNTER_start__n0 + 1; end
       if (__ILA_bar_decode_of_i1__) begin
           i_wb_data <= i_wb_data ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           kp <= kp ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           ki <= ki ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           kd <= kd ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           sp <= sp ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           pv <= pv ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           RS <= RS ;
       end
       if (__ILA_bar_decode_of_i1__) begin
           un <= n4553 ;
       end
   end
end
endmodule
