module FP16_TO_FP17_chn_o_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp16_to_fp17.v:168" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp16_to_fp17.v:169" *)
  output outsig;
  assign outsig = in_0;
endmodule
