module gfx_wbm_read_arbiter(master_busy_o, read_request_o, addr_o, sel_o, dat_i, ack_i, m0_read_request_i, m0_addr_i, m0_sel_i, m0_dat_o, m0_ack_o, m1_read_request_i, m1_addr_i, m1_sel_i, m1_dat_o, m1_ack_o, m2_read_request_i, m2_addr_i, m2_sel_i, m2_dat_o, m2_ack_o);
  wire _00_;
  wire _01_;
  wire _02_;
  wire _03_;
  wire _04_;
  wire [29:0] _05_;
  wire [3:0] _06_;
  input ack_i;
  output [31:2] addr_o;
  input [31:0] dat_i;
  output m0_ack_o;
  input [31:2] m0_addr_i;
  output [31:0] m0_dat_o;
  input m0_read_request_i;
  input [3:0] m0_sel_i;
  output m1_ack_o;
  input [31:2] m1_addr_i;
  output [31:0] m1_dat_o;
  input m1_read_request_i;
  input [3:0] m1_sel_i;
  output m2_ack_o;
  input [31:2] m2_addr_i;
  output [31:0] m2_dat_o;
  input m2_read_request_i;
  input [3:0] m2_sel_i;
  output master_busy_o;
  wire [2:0] master_sel;
  output read_request_o;
  output [3:0] sel_o;
  assign m0_ack_o = ack_i & master_sel[0];
  assign m1_ack_o = ack_i & master_sel[1];
  assign m2_ack_o = ack_i & m2_read_request_i;
  assign _00_ = m0_read_request_i & _01_;
  assign master_sel[0] = _00_ & _02_;
  assign master_sel[1] = m1_read_request_i & _02_;
  assign _01_ = ! m1_read_request_i;
  assign _02_ = ! m2_read_request_i;
  assign _03_ = m2_read_request_i | master_sel[1];
  assign read_request_o = _03_ | master_sel[0];
  assign _04_ = m0_read_request_i | m1_read_request_i;
  assign master_busy_o = _04_ | m2_read_request_i;
  assign _05_ = master_sel[1] ? m1_addr_i : m0_addr_i;
  assign addr_o = m2_read_request_i ? m2_addr_i : _05_;
  assign _06_ = master_sel[1] ? m1_sel_i : m0_sel_i;
  assign sel_o = m2_read_request_i ? m2_sel_i : _06_;
  assign m0_dat_o = dat_i;
  assign m1_dat_o = dat_i;
  assign m2_dat_o = dat_i;
  assign master_sel[2] = m2_read_request_i;
endmodule
