module S(clk, in, out);
  (* src = "S.v:11" *)
  wire [7:0] _000_;
  wire _001_;
  wire _002_;
  wire _003_;
  wire _004_;
  wire _005_;
  wire _006_;
  wire _007_;
  wire _008_;
  wire _009_;
  wire _010_;
  wire _011_;
  wire _012_;
  wire _013_;
  wire _014_;
  wire _015_;
  wire _016_;
  wire _017_;
  wire _018_;
  wire _019_;
  wire _020_;
  wire _021_;
  wire _022_;
  wire _023_;
  wire _024_;
  wire _025_;
  wire _026_;
  wire _027_;
  wire _028_;
  wire _029_;
  wire _030_;
  wire _031_;
  wire _032_;
  wire _033_;
  wire _034_;
  wire _035_;
  wire _036_;
  wire _037_;
  wire _038_;
  wire _039_;
  wire _040_;
  wire _041_;
  wire _042_;
  wire _043_;
  wire _044_;
  wire _045_;
  wire _046_;
  wire _047_;
  wire _048_;
  wire _049_;
  wire _050_;
  wire _051_;
  wire _052_;
  wire _053_;
  wire _054_;
  wire _055_;
  wire _056_;
  wire _057_;
  wire _058_;
  wire _059_;
  wire _060_;
  wire _061_;
  wire _062_;
  wire _063_;
  wire _064_;
  wire _065_;
  wire _066_;
  wire _067_;
  wire _068_;
  wire _069_;
  wire _070_;
  wire _071_;
  wire _072_;
  wire _073_;
  wire _074_;
  wire _075_;
  wire _076_;
  wire _077_;
  wire _078_;
  wire _079_;
  wire _080_;
  wire _081_;
  wire _082_;
  wire _083_;
  wire _084_;
  wire _085_;
  wire _086_;
  wire _087_;
  wire _088_;
  wire _089_;
  wire _090_;
  wire _091_;
  wire _092_;
  wire _093_;
  wire _094_;
  wire _095_;
  wire _096_;
  wire _097_;
  wire _098_;
  wire _099_;
  wire _100_;
  wire _101_;
  wire _102_;
  wire _103_;
  wire _104_;
  wire _105_;
  wire _106_;
  wire _107_;
  wire _108_;
  wire _109_;
  wire _110_;
  wire _111_;
  wire _112_;
  wire _113_;
  wire _114_;
  wire _115_;
  wire _116_;
  wire _117_;
  wire _118_;
  wire _119_;
  wire _120_;
  wire _121_;
  wire _122_;
  wire _123_;
  wire _124_;
  wire _125_;
  wire _126_;
  wire _127_;
  wire _128_;
  wire _129_;
  wire _130_;
  wire _131_;
  wire _132_;
  wire _133_;
  wire _134_;
  wire _135_;
  wire _136_;
  wire _137_;
  wire _138_;
  wire _139_;
  wire _140_;
  wire _141_;
  wire _142_;
  wire _143_;
  wire _144_;
  wire _145_;
  wire _146_;
  wire _147_;
  wire _148_;
  wire _149_;
  wire _150_;
  wire _151_;
  wire _152_;
  wire _153_;
  wire _154_;
  wire _155_;
  wire _156_;
  wire _157_;
  wire _158_;
  wire _159_;
  wire _160_;
  wire _161_;
  wire _162_;
  wire _163_;
  wire _164_;
  wire _165_;
  wire _166_;
  wire _167_;
  wire _168_;
  wire _169_;
  wire _170_;
  wire _171_;
  wire _172_;
  wire _173_;
  wire _174_;
  wire _175_;
  wire _176_;
  wire _177_;
  wire _178_;
  wire _179_;
  wire _180_;
  wire _181_;
  wire _182_;
  wire _183_;
  wire _184_;
  wire _185_;
  wire _186_;
  wire _187_;
  wire _188_;
  wire _189_;
  wire _190_;
  wire _191_;
  wire _192_;
  wire _193_;
  wire _194_;
  wire _195_;
  wire _196_;
  wire _197_;
  wire _198_;
  wire _199_;
  wire _200_;
  wire _201_;
  wire _202_;
  wire _203_;
  wire _204_;
  wire _205_;
  wire _206_;
  wire _207_;
  wire _208_;
  wire _209_;
  wire _210_;
  wire _211_;
  wire _212_;
  wire _213_;
  wire _214_;
  wire _215_;
  wire _216_;
  wire _217_;
  wire _218_;
  wire _219_;
  wire _220_;
  wire _221_;
  wire _222_;
  wire _223_;
  wire _224_;
  wire _225_;
  wire _226_;
  wire _227_;
  wire _228_;
  wire _229_;
  wire _230_;
  wire _231_;
  wire _232_;
  wire _233_;
  wire _234_;
  wire _235_;
  wire _236_;
  wire _237_;
  wire _238_;
  wire _239_;
  wire _240_;
  wire _241_;
  wire _242_;
  wire _243_;
  wire _244_;
  wire _245_;
  wire _246_;
  wire _247_;
  wire _248_;
  wire _249_;
  wire _250_;
  wire _251_;
  wire _252_;
  wire _253_;
  wire _254_;
  wire _255_;
  wire _256_;
  (* src = "S.v:5" *)
  input clk;
  (* src = "S.v:6" *)
  input [7:0] in;
  (* src = "S.v:7" *)
  output [7:0] out;
  reg [7:0] out;
  always @(posedge clk)
      out <= _000_;
  assign _001_ = in == (* src = "S.v:12" *) 8'h9e;
  assign _002_ = in == (* src = "S.v:12" *) 8'h9d;
  assign _003_ = in == (* src = "S.v:12" *) 8'h9c;
  assign _004_ = in == (* src = "S.v:12" *) 8'h9b;
  assign _005_ = in == (* src = "S.v:12" *) 8'h9a;
  assign _006_ = in == (* src = "S.v:12" *) 8'h99;
  assign _007_ = in == (* src = "S.v:12" *) 8'h98;
  assign _008_ = in == (* src = "S.v:12" *) 8'h97;
  assign _009_ = in == (* src = "S.v:12" *) 8'h96;
  assign _010_ = in == (* src = "S.v:12" *) 8'h95;
  assign _011_ = in == (* src = "S.v:12" *) 8'hf8;
  assign _012_ = in == (* src = "S.v:12" *) 8'h94;
  assign _013_ = in == (* src = "S.v:12" *) 8'h93;
  assign _014_ = in == (* src = "S.v:12" *) 8'h92;
  assign _015_ = in == (* src = "S.v:12" *) 8'h91;
  assign _016_ = in == (* src = "S.v:12" *) 8'h90;
  assign _017_ = in == (* src = "S.v:12" *) 8'h8f;
  assign _018_ = in == (* src = "S.v:12" *) 8'h8e;
  assign _019_ = in == (* src = "S.v:12" *) 8'h8d;
  assign _020_ = in == (* src = "S.v:12" *) 8'h8c;
  assign _021_ = in == (* src = "S.v:12" *) 8'h8b;
  assign _022_ = in == (* src = "S.v:12" *) 8'hf7;
  assign _023_ = in == (* src = "S.v:12" *) 8'h8a;
  assign _024_ = in == (* src = "S.v:12" *) 8'h89;
  assign _025_ = in == (* src = "S.v:12" *) 8'h88;
  assign _026_ = in == (* src = "S.v:12" *) 8'h87;
  assign _027_ = in == (* src = "S.v:12" *) 8'h86;
  assign _028_ = in == (* src = "S.v:12" *) 8'h85;
  assign _029_ = in == (* src = "S.v:12" *) 8'h84;
  assign _030_ = in == (* src = "S.v:12" *) 8'h83;
  assign _031_ = in == (* src = "S.v:12" *) 8'h82;
  assign _032_ = in == (* src = "S.v:12" *) 8'h81;
  assign _033_ = in == (* src = "S.v:12" *) 8'hf6;
  assign _034_ = in == (* src = "S.v:12" *) 8'h80;
  assign _035_ = in == (* src = "S.v:12" *) 7'h7f;
  assign _036_ = in == (* src = "S.v:12" *) 7'h7e;
  assign _037_ = in == (* src = "S.v:12" *) 7'h7d;
  assign _038_ = in == (* src = "S.v:12" *) 7'h7c;
  assign _039_ = in == (* src = "S.v:12" *) 7'h7b;
  assign _040_ = in == (* src = "S.v:12" *) 7'h7a;
  assign _041_ = in == (* src = "S.v:12" *) 7'h79;
  assign _042_ = in == (* src = "S.v:12" *) 7'h78;
  assign _043_ = in == (* src = "S.v:12" *) 7'h77;
  assign _044_ = in == (* src = "S.v:12" *) 8'hf5;
  assign _045_ = in == (* src = "S.v:12" *) 7'h76;
  assign _046_ = in == (* src = "S.v:12" *) 7'h75;
  assign _047_ = in == (* src = "S.v:12" *) 7'h74;
  assign _048_ = in == (* src = "S.v:12" *) 7'h73;
  assign _049_ = in == (* src = "S.v:12" *) 7'h72;
  assign _050_ = in == (* src = "S.v:12" *) 7'h71;
  assign _051_ = in == (* src = "S.v:12" *) 7'h70;
  assign _052_ = in == (* src = "S.v:12" *) 7'h6f;
  assign _053_ = in == (* src = "S.v:12" *) 7'h6e;
  assign _054_ = in == (* src = "S.v:12" *) 7'h6d;
  assign _055_ = in == (* src = "S.v:12" *) 8'hf4;
  assign _056_ = in == (* src = "S.v:12" *) 7'h6c;
  assign _057_ = in == (* src = "S.v:12" *) 7'h6b;
  assign _058_ = in == (* src = "S.v:12" *) 7'h6a;
  assign _059_ = in == (* src = "S.v:12" *) 7'h69;
  assign _060_ = in == (* src = "S.v:12" *) 7'h68;
  assign _061_ = in == (* src = "S.v:12" *) 7'h67;
  assign _062_ = in == (* src = "S.v:12" *) 7'h66;
  assign _063_ = in == (* src = "S.v:12" *) 7'h65;
  assign _064_ = in == (* src = "S.v:12" *) 7'h64;
  assign _065_ = in == (* src = "S.v:12" *) 7'h63;
  assign _066_ = in == (* src = "S.v:12" *) 8'hf3;
  assign _067_ = in == (* src = "S.v:12" *) 7'h62;
  assign _068_ = in == (* src = "S.v:12" *) 7'h61;
  assign _069_ = in == (* src = "S.v:12" *) 7'h60;
  assign _070_ = in == (* src = "S.v:12" *) 7'h5f;
  assign _071_ = in == (* src = "S.v:12" *) 7'h5e;
  assign _072_ = in == (* src = "S.v:12" *) 7'h5d;
  assign _073_ = in == (* src = "S.v:12" *) 7'h5c;
  assign _074_ = in == (* src = "S.v:12" *) 7'h5b;
  assign _075_ = in == (* src = "S.v:12" *) 7'h5a;
  assign _076_ = in == (* src = "S.v:12" *) 7'h59;
  assign _077_ = in == (* src = "S.v:12" *) 8'hf2;
  assign _078_ = in == (* src = "S.v:12" *) 7'h58;
  assign _079_ = in == (* src = "S.v:12" *) 7'h57;
  assign _080_ = in == (* src = "S.v:12" *) 7'h56;
  assign _081_ = in == (* src = "S.v:12" *) 7'h55;
  assign _082_ = in == (* src = "S.v:12" *) 7'h54;
  assign _083_ = in == (* src = "S.v:12" *) 7'h53;
  assign _084_ = in == (* src = "S.v:12" *) 7'h52;
  assign _085_ = in == (* src = "S.v:12" *) 7'h51;
  assign _086_ = in == (* src = "S.v:12" *) 7'h50;
  assign _087_ = in == (* src = "S.v:12" *) 7'h4f;
  assign _088_ = in == (* src = "S.v:12" *) 8'hf1;
  assign _089_ = in == (* src = "S.v:12" *) 7'h4e;
  assign _090_ = in == (* src = "S.v:12" *) 7'h4d;
  assign _091_ = in == (* src = "S.v:12" *) 7'h4c;
  assign _092_ = in == (* src = "S.v:12" *) 7'h4b;
  assign _093_ = in == (* src = "S.v:12" *) 7'h4a;
  assign _094_ = in == (* src = "S.v:12" *) 7'h49;
  assign _095_ = in == (* src = "S.v:12" *) 7'h48;
  assign _096_ = in == (* src = "S.v:12" *) 7'h47;
  assign _097_ = in == (* src = "S.v:12" *) 7'h46;
  assign _098_ = in == (* src = "S.v:12" *) 7'h45;
  assign _099_ = in == (* src = "S.v:12" *) 8'hf0;
  assign _100_ = in == (* src = "S.v:12" *) 7'h44;
  assign _101_ = in == (* src = "S.v:12" *) 7'h43;
  assign _102_ = in == (* src = "S.v:12" *) 7'h42;
  assign _103_ = in == (* src = "S.v:12" *) 7'h41;
  assign _104_ = in == (* src = "S.v:12" *) 7'h40;
  assign _105_ = in == (* src = "S.v:12" *) 6'h3f;
  assign _106_ = in == (* src = "S.v:12" *) 6'h3e;
  assign _107_ = in == (* src = "S.v:12" *) 6'h3d;
  assign _108_ = in == (* src = "S.v:12" *) 6'h3c;
  assign _109_ = in == (* src = "S.v:12" *) 6'h3b;
  assign _110_ = in == (* src = "S.v:12" *) 8'hef;
  function [7:0] _368_;
    input [7:0] a;
    input [2047:0] b;
    input [255:0] s;
    (* src = "S.v:12" *)
    (* parallel_case *)
    casez (s)
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1:
        _368_ = b[7:0];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?:
        _368_ = b[15:8];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??:
        _368_ = b[23:16];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???:
        _368_ = b[31:24];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????:
        _368_ = b[39:32];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????:
        _368_ = b[47:40];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????:
        _368_ = b[55:48];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????:
        _368_ = b[63:56];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????:
        _368_ = b[71:64];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????:
        _368_ = b[79:72];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????:
        _368_ = b[87:80];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????:
        _368_ = b[95:88];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????:
        _368_ = b[103:96];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????:
        _368_ = b[111:104];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????:
        _368_ = b[119:112];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????:
        _368_ = b[127:120];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????:
        _368_ = b[135:128];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????:
        _368_ = b[143:136];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????:
        _368_ = b[151:144];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????:
        _368_ = b[159:152];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????:
        _368_ = b[167:160];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????:
        _368_ = b[175:168];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????:
        _368_ = b[183:176];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????:
        _368_ = b[191:184];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????:
        _368_ = b[199:192];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????:
        _368_ = b[207:200];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????:
        _368_ = b[215:208];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????:
        _368_ = b[223:216];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????:
        _368_ = b[231:224];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????:
        _368_ = b[239:232];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????:
        _368_ = b[247:240];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????:
        _368_ = b[255:248];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????:
        _368_ = b[263:256];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????:
        _368_ = b[271:264];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????:
        _368_ = b[279:272];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????:
        _368_ = b[287:280];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????:
        _368_ = b[295:288];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????:
        _368_ = b[303:296];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????:
        _368_ = b[311:304];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????:
        _368_ = b[319:312];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????:
        _368_ = b[327:320];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????:
        _368_ = b[335:328];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????:
        _368_ = b[343:336];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????:
        _368_ = b[351:344];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????:
        _368_ = b[359:352];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????:
        _368_ = b[367:360];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????:
        _368_ = b[375:368];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????:
        _368_ = b[383:376];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????:
        _368_ = b[391:384];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????:
        _368_ = b[399:392];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????:
        _368_ = b[407:400];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????:
        _368_ = b[415:408];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????:
        _368_ = b[423:416];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????:
        _368_ = b[431:424];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????:
        _368_ = b[439:432];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????:
        _368_ = b[447:440];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????:
        _368_ = b[455:448];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????:
        _368_ = b[463:456];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????:
        _368_ = b[471:464];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????:
        _368_ = b[479:472];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????:
        _368_ = b[487:480];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????:
        _368_ = b[495:488];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????:
        _368_ = b[503:496];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????:
        _368_ = b[511:504];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????:
        _368_ = b[519:512];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????:
        _368_ = b[527:520];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????:
        _368_ = b[535:528];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????:
        _368_ = b[543:536];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????:
        _368_ = b[551:544];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????:
        _368_ = b[559:552];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????:
        _368_ = b[567:560];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????:
        _368_ = b[575:568];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????:
        _368_ = b[583:576];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????:
        _368_ = b[591:584];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????:
        _368_ = b[599:592];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????:
        _368_ = b[607:600];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????:
        _368_ = b[615:608];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????:
        _368_ = b[623:616];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????:
        _368_ = b[631:624];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????:
        _368_ = b[639:632];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[647:640];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[655:648];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[663:656];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[671:664];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[679:672];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[687:680];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[695:688];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[703:696];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[711:704];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[719:712];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[727:720];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[735:728];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[743:736];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[751:744];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[759:752];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[767:760];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[775:768];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[783:776];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[791:784];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[799:792];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[807:800];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[815:808];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[823:816];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[831:824];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[839:832];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[847:840];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[855:848];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[863:856];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[871:864];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[879:872];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[887:880];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[895:888];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[903:896];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[911:904];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[919:912];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[927:920];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[935:928];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[943:936];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[951:944];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[959:952];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[967:960];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[975:968];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[983:976];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[991:984];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[999:992];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1007:1000];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1015:1008];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1023:1016];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1031:1024];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1039:1032];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1047:1040];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1055:1048];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1063:1056];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1071:1064];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1079:1072];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1087:1080];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1095:1088];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1103:1096];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1111:1104];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1119:1112];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1127:1120];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1135:1128];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1143:1136];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1151:1144];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1159:1152];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1167:1160];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1175:1168];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1183:1176];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1191:1184];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1199:1192];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1207:1200];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1215:1208];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1223:1216];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1231:1224];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1239:1232];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1247:1240];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1255:1248];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1263:1256];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1271:1264];
      256'b????????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1279:1272];
      256'b???????????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1287:1280];
      256'b??????????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1295:1288];
      256'b?????????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1303:1296];
      256'b????????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1311:1304];
      256'b???????????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1319:1312];
      256'b??????????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1327:1320];
      256'b?????????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1335:1328];
      256'b????????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1343:1336];
      256'b???????????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1351:1344];
      256'b??????????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1359:1352];
      256'b?????????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1367:1360];
      256'b????????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1375:1368];
      256'b???????????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1383:1376];
      256'b??????????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1391:1384];
      256'b?????????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1399:1392];
      256'b????????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1407:1400];
      256'b???????????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1415:1408];
      256'b??????????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1423:1416];
      256'b?????????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1431:1424];
      256'b????????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1439:1432];
      256'b???????????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1447:1440];
      256'b??????????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1455:1448];
      256'b?????????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1463:1456];
      256'b????????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1471:1464];
      256'b???????????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1479:1472];
      256'b??????????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1487:1480];
      256'b?????????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1495:1488];
      256'b????????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1503:1496];
      256'b???????????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1511:1504];
      256'b??????????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1519:1512];
      256'b?????????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1527:1520];
      256'b????????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1535:1528];
      256'b???????????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1543:1536];
      256'b??????????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1551:1544];
      256'b?????????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1559:1552];
      256'b????????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1567:1560];
      256'b???????????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1575:1568];
      256'b??????????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1583:1576];
      256'b?????????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1591:1584];
      256'b????????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1599:1592];
      256'b???????????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1607:1600];
      256'b??????????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1615:1608];
      256'b?????????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1623:1616];
      256'b????????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1631:1624];
      256'b???????????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1639:1632];
      256'b??????????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1647:1640];
      256'b?????????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1655:1648];
      256'b????????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1663:1656];
      256'b???????????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1671:1664];
      256'b??????????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1679:1672];
      256'b?????????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1687:1680];
      256'b????????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1695:1688];
      256'b???????????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1703:1696];
      256'b??????????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1711:1704];
      256'b?????????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1719:1712];
      256'b????????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1727:1720];
      256'b???????????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1735:1728];
      256'b??????????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1743:1736];
      256'b?????????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1751:1744];
      256'b????????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1759:1752];
      256'b???????????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1767:1760];
      256'b??????????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1775:1768];
      256'b?????????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1783:1776];
      256'b????????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1791:1784];
      256'b???????????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1799:1792];
      256'b??????????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1807:1800];
      256'b?????????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1815:1808];
      256'b????????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1823:1816];
      256'b???????????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1831:1824];
      256'b??????????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1839:1832];
      256'b?????????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1847:1840];
      256'b????????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1855:1848];
      256'b???????????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1863:1856];
      256'b??????????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1871:1864];
      256'b?????????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1879:1872];
      256'b????????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1887:1880];
      256'b???????????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1895:1888];
      256'b??????????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1903:1896];
      256'b?????????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1911:1904];
      256'b????????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1919:1912];
      256'b???????????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1927:1920];
      256'b??????????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1935:1928];
      256'b?????????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1943:1936];
      256'b????????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1951:1944];
      256'b???????????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1959:1952];
      256'b??????????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1967:1960];
      256'b?????????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1975:1968];
      256'b????????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1983:1976];
      256'b???????1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1991:1984];
      256'b??????1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[1999:1992];
      256'b?????1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[2007:2000];
      256'b????1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[2015:2008];
      256'b???1????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[2023:2016];
      256'b??1?????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[2031:2024];
      256'b?1??????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[2039:2032];
      256'b1???????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????????:
        _368_ = b[2047:2040];
      default:
        _368_ = a;
    endcase
  endfunction
  assign _000_ = _368_(out, 2048'h637c777bf26b6fc53001672bfed7ab76ca82c97dfa5947f0add4a2af9ca472c0b7fd9326363ff7cc34a5e5f171d8311504c723c31896059a071280e2eb27b27509832c1a1b6e5aa0523bd6b329e32f8453d100ed20fcb15b6acbbe394a4c58cfd0efaafb434d338545f9027f503c9fa851a3408f929d38f5bcb6da2110fff3d2cd0c13ec5f974417c4a77e3d645d197360814fdc222a908846eeb814de5e0bdbe0323a0a4906245cc2d3ac629195e479e7c8376d8dd54ea96c56f4ea657aae08ba78252e1ca6b4c6e8dd741f4bbd8b8a703eb5664803f60e613557b986c11d9ee1f8981169d98e949b1e87e9ce5528df8ca1890dbfe6426841992d0fb054bb16, { _174_, _173_, _172_, _171_, _170_, _169_, _168_, _167_, _166_, _164_, _163_, _162_, _161_, _160_, _159_, _158_, _157_, _156_, _155_, _153_, _152_, _151_, _150_, _149_, _148_, _147_, _146_, _145_, _144_, _142_, _141_, _140_, _139_, _138_, _137_, _136_, _135_, _134_, _133_, _131_, _130_, _129_, _128_, _127_, _126_, _125_, _124_, _123_, _122_, _120_, _119_, _118_, _117_, _116_, _115_, _114_, _113_, _112_, _111_, _109_, _108_, _107_, _106_, _105_, _104_, _103_, _102_, _101_, _100_, _098_, _097_, _096_, _095_, _094_, _093_, _092_, _091_, _090_, _089_, _087_, _086_, _085_, _084_, _083_, _082_, _081_, _080_, _079_, _078_, _076_, _075_, _074_, _073_, _072_, _071_, _070_, _069_, _068_, _067_, _065_, _064_, _063_, _062_, _061_, _060_, _059_, _058_, _057_, _056_, _054_, _053_, _052_, _051_, _050_, _049_, _048_, _047_, _046_, _045_, _043_, _042_, _041_, _040_, _039_, _038_, _037_, _036_, _035_, _034_, _032_, _031_, _030_, _029_, _028_, _027_, _026_, _025_, _024_, _023_, _021_, _020_, _019_, _018_, _017_, _016_, _015_, _014_, _013_, _012_, _010_, _009_, _008_, _007_, _006_, _005_, _004_, _003_, _002_, _001_, _255_, _254_, _253_, _252_, _251_, _250_, _249_, _248_, _247_, _246_, _244_, _243_, _242_, _241_, _240_, _239_, _238_, _237_, _236_, _235_, _233_, _232_, _231_, _230_, _229_, _228_, _227_, _226_, _225_, _224_, _222_, _221_, _220_, _219_, _218_, _217_, _216_, _215_, _214_, _213_, _211_, _210_, _209_, _208_, _207_, _206_, _205_, _204_, _203_, _202_, _200_, _199_, _198_, _197_, _196_, _195_, _194_, _193_, _192_, _191_, _189_, _188_, _187_, _186_, _185_, _184_, _183_, _182_, _181_, _180_, _179_, _178_, _177_, _176_, _175_, _165_, _154_, _143_, _132_, _121_, _110_, _099_, _088_, _077_, _066_, _055_, _044_, _033_, _022_, _011_, _256_, _245_, _234_, _223_, _212_, _201_, _190_ });
  assign _111_ = in == (* src = "S.v:12" *) 6'h3a;
  assign _112_ = in == (* src = "S.v:12" *) 6'h39;
  assign _113_ = in == (* src = "S.v:12" *) 6'h38;
  assign _114_ = in == (* src = "S.v:12" *) 6'h37;
  assign _115_ = in == (* src = "S.v:12" *) 6'h36;
  assign _116_ = in == (* src = "S.v:12" *) 6'h35;
  assign _117_ = in == (* src = "S.v:12" *) 6'h34;
  assign _118_ = in == (* src = "S.v:12" *) 6'h33;
  assign _119_ = in == (* src = "S.v:12" *) 6'h32;
  assign _120_ = in == (* src = "S.v:12" *) 6'h31;
  assign _121_ = in == (* src = "S.v:12" *) 8'hee;
  assign _122_ = in == (* src = "S.v:12" *) 6'h30;
  assign _123_ = in == (* src = "S.v:12" *) 6'h2f;
  assign _124_ = in == (* src = "S.v:12" *) 6'h2e;
  assign _125_ = in == (* src = "S.v:12" *) 6'h2d;
  assign _126_ = in == (* src = "S.v:12" *) 6'h2c;
  assign _127_ = in == (* src = "S.v:12" *) 6'h2b;
  assign _128_ = in == (* src = "S.v:12" *) 6'h2a;
  assign _129_ = in == (* src = "S.v:12" *) 6'h29;
  assign _130_ = in == (* src = "S.v:12" *) 6'h28;
  assign _131_ = in == (* src = "S.v:12" *) 6'h27;
  assign _132_ = in == (* src = "S.v:12" *) 8'hed;
  assign _133_ = in == (* src = "S.v:12" *) 6'h26;
  assign _134_ = in == (* src = "S.v:12" *) 6'h25;
  assign _135_ = in == (* src = "S.v:12" *) 6'h24;
  assign _136_ = in == (* src = "S.v:12" *) 6'h23;
  assign _137_ = in == (* src = "S.v:12" *) 6'h22;
  assign _138_ = in == (* src = "S.v:12" *) 6'h21;
  assign _139_ = in == (* src = "S.v:12" *) 6'h20;
  assign _140_ = in == (* src = "S.v:12" *) 5'h1f;
  assign _141_ = in == (* src = "S.v:12" *) 5'h1e;
  assign _142_ = in == (* src = "S.v:12" *) 5'h1d;
  assign _143_ = in == (* src = "S.v:12" *) 8'hec;
  assign _144_ = in == (* src = "S.v:12" *) 5'h1c;
  assign _145_ = in == (* src = "S.v:12" *) 5'h1b;
  assign _146_ = in == (* src = "S.v:12" *) 5'h1a;
  assign _147_ = in == (* src = "S.v:12" *) 5'h19;
  assign _148_ = in == (* src = "S.v:12" *) 5'h18;
  assign _149_ = in == (* src = "S.v:12" *) 5'h17;
  assign _150_ = in == (* src = "S.v:12" *) 5'h16;
  assign _151_ = in == (* src = "S.v:12" *) 5'h15;
  assign _152_ = in == (* src = "S.v:12" *) 5'h14;
  assign _153_ = in == (* src = "S.v:12" *) 5'h13;
  assign _154_ = in == (* src = "S.v:12" *) 8'heb;
  assign _155_ = in == (* src = "S.v:12" *) 5'h12;
  assign _156_ = in == (* src = "S.v:12" *) 5'h11;
  assign _157_ = in == (* src = "S.v:12" *) 5'h10;
  assign _158_ = in == (* src = "S.v:12" *) 4'hf;
  assign _159_ = in == (* src = "S.v:12" *) 4'he;
  assign _160_ = in == (* src = "S.v:12" *) 4'hd;
  assign _161_ = in == (* src = "S.v:12" *) 4'hc;
  assign _162_ = in == (* src = "S.v:12" *) 4'hb;
  assign _163_ = in == (* src = "S.v:12" *) 4'ha;
  assign _164_ = in == (* src = "S.v:12" *) 4'h9;
  assign _165_ = in == (* src = "S.v:12" *) 8'hea;
  assign _166_ = in == (* src = "S.v:12" *) 4'h8;
  assign _167_ = in == (* src = "S.v:12" *) 3'h7;
  assign _168_ = in == (* src = "S.v:12" *) 3'h6;
  assign _169_ = in == (* src = "S.v:12" *) 3'h5;
  assign _170_ = in == (* src = "S.v:12" *) 3'h4;
  assign _171_ = in == (* src = "S.v:12" *) 2'h3;
  assign _172_ = in == (* src = "S.v:12" *) 2'h2;
  assign _173_ = in == (* src = "S.v:12" *) 1'h1;
  assign _174_ = ! (* src = "S.v:12" *) in;
  assign _175_ = in == (* src = "S.v:12" *) 8'he9;
  assign _176_ = in == (* src = "S.v:12" *) 8'he8;
  assign _177_ = in == (* src = "S.v:12" *) 8'he7;
  assign _178_ = in == (* src = "S.v:12" *) 8'he6;
  assign _179_ = in == (* src = "S.v:12" *) 8'he5;
  assign _180_ = in == (* src = "S.v:12" *) 8'he4;
  assign _181_ = in == (* src = "S.v:12" *) 8'he3;
  assign _182_ = in == (* src = "S.v:12" *) 8'he2;
  assign _183_ = in == (* src = "S.v:12" *) 8'he1;
  assign _184_ = in == (* src = "S.v:12" *) 8'he0;
  assign _185_ = in == (* src = "S.v:12" *) 8'hdf;
  assign _186_ = in == (* src = "S.v:12" *) 8'hde;
  assign _187_ = in == (* src = "S.v:12" *) 8'hdd;
  assign _188_ = in == (* src = "S.v:12" *) 8'hdc;
  assign _189_ = in == (* src = "S.v:12" *) 8'hdb;
  assign _190_ = in == (* src = "S.v:12" *) 8'hff;
  assign _191_ = in == (* src = "S.v:12" *) 8'hda;
  assign _192_ = in == (* src = "S.v:12" *) 8'hd9;
  assign _193_ = in == (* src = "S.v:12" *) 8'hd8;
  assign _194_ = in == (* src = "S.v:12" *) 8'hd7;
  assign _195_ = in == (* src = "S.v:12" *) 8'hd6;
  assign _196_ = in == (* src = "S.v:12" *) 8'hd5;
  assign _197_ = in == (* src = "S.v:12" *) 8'hd4;
  assign _198_ = in == (* src = "S.v:12" *) 8'hd3;
  assign _199_ = in == (* src = "S.v:12" *) 8'hd2;
  assign _200_ = in == (* src = "S.v:12" *) 8'hd1;
  assign _201_ = in == (* src = "S.v:12" *) 8'hfe;
  assign _202_ = in == (* src = "S.v:12" *) 8'hd0;
  assign _203_ = in == (* src = "S.v:12" *) 8'hcf;
  assign _204_ = in == (* src = "S.v:12" *) 8'hce;
  assign _205_ = in == (* src = "S.v:12" *) 8'hcd;
  assign _206_ = in == (* src = "S.v:12" *) 8'hcc;
  assign _207_ = in == (* src = "S.v:12" *) 8'hcb;
  assign _208_ = in == (* src = "S.v:12" *) 8'hca;
  assign _209_ = in == (* src = "S.v:12" *) 8'hc9;
  assign _210_ = in == (* src = "S.v:12" *) 8'hc8;
  assign _211_ = in == (* src = "S.v:12" *) 8'hc7;
  assign _212_ = in == (* src = "S.v:12" *) 8'hfd;
  assign _213_ = in == (* src = "S.v:12" *) 8'hc6;
  assign _214_ = in == (* src = "S.v:12" *) 8'hc5;
  assign _215_ = in == (* src = "S.v:12" *) 8'hc4;
  assign _216_ = in == (* src = "S.v:12" *) 8'hc3;
  assign _217_ = in == (* src = "S.v:12" *) 8'hc2;
  assign _218_ = in == (* src = "S.v:12" *) 8'hc1;
  assign _219_ = in == (* src = "S.v:12" *) 8'hc0;
  assign _220_ = in == (* src = "S.v:12" *) 8'hbf;
  assign _221_ = in == (* src = "S.v:12" *) 8'hbe;
  assign _222_ = in == (* src = "S.v:12" *) 8'hbd;
  assign _223_ = in == (* src = "S.v:12" *) 8'hfc;
  assign _224_ = in == (* src = "S.v:12" *) 8'hbc;
  assign _225_ = in == (* src = "S.v:12" *) 8'hbb;
  assign _226_ = in == (* src = "S.v:12" *) 8'hba;
  assign _227_ = in == (* src = "S.v:12" *) 8'hb9;
  assign _228_ = in == (* src = "S.v:12" *) 8'hb8;
  assign _229_ = in == (* src = "S.v:12" *) 8'hb7;
  assign _230_ = in == (* src = "S.v:12" *) 8'hb6;
  assign _231_ = in == (* src = "S.v:12" *) 8'hb5;
  assign _232_ = in == (* src = "S.v:12" *) 8'hb4;
  assign _233_ = in == (* src = "S.v:12" *) 8'hb3;
  assign _234_ = in == (* src = "S.v:12" *) 8'hfb;
  assign _235_ = in == (* src = "S.v:12" *) 8'hb2;
  assign _236_ = in == (* src = "S.v:12" *) 8'hb1;
  assign _237_ = in == (* src = "S.v:12" *) 8'hb0;
  assign _238_ = in == (* src = "S.v:12" *) 8'haf;
  assign _239_ = in == (* src = "S.v:12" *) 8'hae;
  assign _240_ = in == (* src = "S.v:12" *) 8'had;
  assign _241_ = in == (* src = "S.v:12" *) 8'hac;
  assign _242_ = in == (* src = "S.v:12" *) 8'hab;
  assign _243_ = in == (* src = "S.v:12" *) 8'haa;
  assign _244_ = in == (* src = "S.v:12" *) 8'ha9;
  assign _245_ = in == (* src = "S.v:12" *) 8'hfa;
  assign _246_ = in == (* src = "S.v:12" *) 8'ha8;
  assign _247_ = in == (* src = "S.v:12" *) 8'ha7;
  assign _248_ = in == (* src = "S.v:12" *) 8'ha6;
  assign _249_ = in == (* src = "S.v:12" *) 8'ha5;
  assign _250_ = in == (* src = "S.v:12" *) 8'ha4;
  assign _251_ = in == (* src = "S.v:12" *) 8'ha3;
  assign _252_ = in == (* src = "S.v:12" *) 8'ha2;
  assign _253_ = in == (* src = "S.v:12" *) 8'ha1;
  assign _254_ = in == (* src = "S.v:12" *) 8'ha0;
  assign _255_ = in == (* src = "S.v:12" *) 8'h9f;
  assign _256_ = in == (* src = "S.v:12" *) 8'hf9;
endmodule
