module FP17_ADD_chn_o_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_add.v:277" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:278" *)
  output outsig;
  assign outsig = in_0;
endmodule
