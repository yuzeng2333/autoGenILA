module FP17_MUL_chn_o_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_mul.v:74" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_mul.v:75" *)
  output outsig;
  assign outsig = in_0;
endmodule
