module NV_NVDLA_CACC_calculator(nvdla_core_clk, nvdla_core_rstn, abuf_rd_data_0, abuf_rd_data_1, abuf_rd_data_2, abuf_rd_data_3, abuf_rd_data_4, abuf_rd_data_5, abuf_rd_data_6, abuf_rd_data_7, accu_ctrl_pd, accu_ctrl_ram_valid, accu_ctrl_valid, cfg_in_en_mask, cfg_is_fp, cfg_is_int, cfg_is_int8, cfg_is_wg, cfg_truncate, mac_a2accu_data0, mac_a2accu_data1, mac_a2accu_data2, mac_a2accu_data3, mac_a2accu_data4, mac_a2accu_data5, mac_a2accu_data6, mac_a2accu_data7, mac_a2accu_mask, mac_a2accu_mode, mac_a2accu_pvld, mac_b2accu_data0, mac_b2accu_data1, mac_b2accu_data2, mac_b2accu_data3, mac_b2accu_data4, mac_b2accu_data5, mac_b2accu_data6, mac_b2accu_data7, mac_b2accu_mask, mac_b2accu_mode, mac_b2accu_pvld, nvdla_cell_clk_0, nvdla_cell_clk_1, nvdla_cell_clk_2, nvdla_cell_clk_3, abuf_wr_addr, abuf_wr_data_0, abuf_wr_data_1, abuf_wr_data_2, abuf_wr_data_3, abuf_wr_data_4, abuf_wr_data_5, abuf_wr_data_6, abuf_wr_data_7, abuf_wr_en, dlv_data_0, dlv_data_1, dlv_data_2, dlv_data_3, dlv_data_4, dlv_data_5, dlv_data_6, dlv_data_7, dlv_mask, dlv_pd, dlv_valid, dp2reg_sat_count);
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12584" *)
  wire [4:0] _0000_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12645" *)
  wire [767:0] _0001_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12655" *)
  wire [767:0] _0002_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12665" *)
  wire [767:0] _0003_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12675" *)
  wire [767:0] _0004_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12685" *)
  wire [543:0] _0005_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12695" *)
  wire [543:0] _0006_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12705" *)
  wire [543:0] _0007_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12715" *)
  wire [543:0] _0008_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7137" *)
  wire [4:0] _0009_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10581" *)
  wire [4:0] _0010_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10710" *)
  wire [4:0] _0011_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10839" *)
  wire [4:0] _0012_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2279" *)
  wire [131:0] _0013_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2269" *)
  wire [43:0] _0014_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2479" *)
  wire [131:0] _0015_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2469" *)
  wire [43:0] _0016_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2499" *)
  wire [131:0] _0017_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2489" *)
  wire [43:0] _0018_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2519" *)
  wire [131:0] _0019_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2509" *)
  wire [43:0] _0020_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2539" *)
  wire [131:0] _0021_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2529" *)
  wire [43:0] _0022_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2559" *)
  wire [131:0] _0023_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2549" *)
  wire [43:0] _0024_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2579" *)
  wire [131:0] _0025_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2569" *)
  wire [43:0] _0026_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2299" *)
  wire [131:0] _0027_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2289" *)
  wire [43:0] _0028_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2319" *)
  wire [131:0] _0029_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2309" *)
  wire [43:0] _0030_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2339" *)
  wire [131:0] _0031_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2329" *)
  wire [43:0] _0032_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2359" *)
  wire [131:0] _0033_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2349" *)
  wire [43:0] _0034_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2379" *)
  wire [131:0] _0035_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2369" *)
  wire [43:0] _0036_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2399" *)
  wire [131:0] _0037_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2389" *)
  wire [43:0] _0038_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2419" *)
  wire [131:0] _0039_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2409" *)
  wire [43:0] _0040_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2439" *)
  wire [131:0] _0041_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2429" *)
  wire [43:0] _0042_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2459" *)
  wire [131:0] _0043_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2449" *)
  wire [43:0] _0044_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7205" *)
  wire [7:0] _0045_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10913" *)
  wire [7:0] _0046_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11103" *)
  wire [7:0] _0047_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11293" *)
  wire [7:0] _0048_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11483" *)
  wire [7:0] _0049_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7693" *)
  wire [63:0] _0050_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7632" *)
  wire [127:0] _0051_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2612" *)
  wire [191:0] _0052_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7327" *)
  wire _0053_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11035" *)
  wire _0054_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11225" *)
  wire _0055_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11415" *)
  wire _0056_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11605" *)
  wire _0057_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4509" *)
  wire [43:0] _0058_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4609" *)
  wire [43:0] _0059_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4619" *)
  wire [43:0] _0060_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4629" *)
  wire [43:0] _0061_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4639" *)
  wire [43:0] _0062_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4649" *)
  wire [43:0] _0063_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4659" *)
  wire [43:0] _0064_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4669" *)
  wire [43:0] _0065_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4679" *)
  wire [43:0] _0066_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4689" *)
  wire [43:0] _0067_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4699" *)
  wire [43:0] _0068_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4519" *)
  wire [43:0] _0069_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4709" *)
  wire [43:0] _0070_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4719" *)
  wire [43:0] _0071_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4729" *)
  wire [43:0] _0072_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4739" *)
  wire [43:0] _0073_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4749" *)
  wire [43:0] _0074_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4759" *)
  wire [43:0] _0075_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4769" *)
  wire [43:0] _0076_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4779" *)
  wire [43:0] _0077_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4789" *)
  wire [43:0] _0078_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4799" *)
  wire [43:0] _0079_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4529" *)
  wire [43:0] _0080_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4809" *)
  wire [43:0] _0081_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4819" *)
  wire [43:0] _0082_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4829" *)
  wire [43:0] _0083_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4839" *)
  wire [43:0] _0084_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4849" *)
  wire [43:0] _0085_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4859" *)
  wire [43:0] _0086_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4869" *)
  wire [43:0] _0087_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4879" *)
  wire [43:0] _0088_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4889" *)
  wire [43:0] _0089_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4899" *)
  wire [43:0] _0090_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4539" *)
  wire [43:0] _0091_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4909" *)
  wire [43:0] _0092_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4919" *)
  wire [43:0] _0093_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4929" *)
  wire [43:0] _0094_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4939" *)
  wire [43:0] _0095_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4949" *)
  wire [43:0] _0096_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4959" *)
  wire [43:0] _0097_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4969" *)
  wire [43:0] _0098_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4979" *)
  wire [43:0] _0099_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4989" *)
  wire [43:0] _0100_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4999" *)
  wire [43:0] _0101_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4549" *)
  wire [43:0] _0102_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5009" *)
  wire [43:0] _0103_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5019" *)
  wire [43:0] _0104_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5029" *)
  wire [43:0] _0105_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5039" *)
  wire [43:0] _0106_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5049" *)
  wire [43:0] _0107_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5059" *)
  wire [43:0] _0108_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5069" *)
  wire [43:0] _0109_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5079" *)
  wire [43:0] _0110_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5089" *)
  wire [43:0] _0111_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5099" *)
  wire [43:0] _0112_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4559" *)
  wire [43:0] _0113_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5109" *)
  wire [43:0] _0114_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5119" *)
  wire [43:0] _0115_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5129" *)
  wire [43:0] _0116_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5139" *)
  wire [43:0] _0117_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4569" *)
  wire [43:0] _0118_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4579" *)
  wire [43:0] _0119_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4589" *)
  wire [43:0] _0120_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4599" *)
  wire [43:0] _0121_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3229" *)
  wire [37:0] _0122_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4229" *)
  wire [21:0] _0123_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4239" *)
  wire [21:0] _0124_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4249" *)
  wire [21:0] _0125_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4259" *)
  wire [21:0] _0126_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4269" *)
  wire [21:0] _0127_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4279" *)
  wire [21:0] _0128_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4289" *)
  wire [21:0] _0129_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4299" *)
  wire [21:0] _0130_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4309" *)
  wire [21:0] _0131_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4319" *)
  wire [21:0] _0132_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3329" *)
  wire [37:0] _0133_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4329" *)
  wire [21:0] _0134_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4339" *)
  wire [21:0] _0135_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4349" *)
  wire [21:0] _0136_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4359" *)
  wire [21:0] _0137_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4369" *)
  wire [21:0] _0138_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4379" *)
  wire [21:0] _0139_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4389" *)
  wire [21:0] _0140_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4399" *)
  wire [21:0] _0141_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4409" *)
  wire [21:0] _0142_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4419" *)
  wire [21:0] _0143_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3339" *)
  wire [37:0] _0144_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4429" *)
  wire [21:0] _0145_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4439" *)
  wire [21:0] _0146_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4449" *)
  wire [21:0] _0147_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4459" *)
  wire [21:0] _0148_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4469" *)
  wire [21:0] _0149_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4479" *)
  wire [21:0] _0150_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4489" *)
  wire [21:0] _0151_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4499" *)
  wire [21:0] _0152_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3349" *)
  wire [37:0] _0153_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3359" *)
  wire [37:0] _0154_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3369" *)
  wire [37:0] _0155_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3379" *)
  wire [37:0] _0156_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3389" *)
  wire [37:0] _0157_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3399" *)
  wire [37:0] _0158_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3409" *)
  wire [37:0] _0159_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3419" *)
  wire [37:0] _0160_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3239" *)
  wire [37:0] _0161_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3429" *)
  wire [37:0] _0162_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3439" *)
  wire [37:0] _0163_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3449" *)
  wire [37:0] _0164_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3459" *)
  wire [37:0] _0165_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3469" *)
  wire [37:0] _0166_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3479" *)
  wire [37:0] _0167_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3489" *)
  wire [37:0] _0168_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3499" *)
  wire [37:0] _0169_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3509" *)
  wire [37:0] _0170_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3519" *)
  wire [37:0] _0171_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3249" *)
  wire [37:0] _0172_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3529" *)
  wire [37:0] _0173_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3539" *)
  wire [37:0] _0174_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3549" *)
  wire [37:0] _0175_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3559" *)
  wire [37:0] _0176_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3569" *)
  wire [37:0] _0177_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3579" *)
  wire [37:0] _0178_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3589" *)
  wire [37:0] _0179_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3599" *)
  wire [37:0] _0180_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3609" *)
  wire [37:0] _0181_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3619" *)
  wire [37:0] _0182_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3259" *)
  wire [37:0] _0183_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3629" *)
  wire [37:0] _0184_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3639" *)
  wire [37:0] _0185_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3649" *)
  wire [37:0] _0186_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3659" *)
  wire [37:0] _0187_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3669" *)
  wire [37:0] _0188_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3679" *)
  wire [37:0] _0189_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3689" *)
  wire [37:0] _0190_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3699" *)
  wire [37:0] _0191_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3709" *)
  wire [37:0] _0192_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3719" *)
  wire [37:0] _0193_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3269" *)
  wire [37:0] _0194_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3729" *)
  wire [37:0] _0195_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3739" *)
  wire [37:0] _0196_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3749" *)
  wire [37:0] _0197_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3759" *)
  wire [37:0] _0198_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3769" *)
  wire [37:0] _0199_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3779" *)
  wire [37:0] _0200_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3789" *)
  wire [37:0] _0201_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3799" *)
  wire [37:0] _0202_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3809" *)
  wire [37:0] _0203_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3819" *)
  wire [37:0] _0204_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3279" *)
  wire [37:0] _0205_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3829" *)
  wire [37:0] _0206_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3839" *)
  wire [37:0] _0207_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3849" *)
  wire [37:0] _0208_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3859" *)
  wire [37:0] _0209_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3869" *)
  wire [21:0] _0210_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3879" *)
  wire [21:0] _0211_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3889" *)
  wire [21:0] _0212_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3899" *)
  wire [21:0] _0213_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3909" *)
  wire [21:0] _0214_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3919" *)
  wire [21:0] _0215_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3289" *)
  wire [37:0] _0216_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3929" *)
  wire [21:0] _0217_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3939" *)
  wire [21:0] _0218_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3949" *)
  wire [21:0] _0219_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3959" *)
  wire [21:0] _0220_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3969" *)
  wire [21:0] _0221_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3979" *)
  wire [21:0] _0222_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3989" *)
  wire [21:0] _0223_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3999" *)
  wire [21:0] _0224_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4009" *)
  wire [21:0] _0225_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4019" *)
  wire [21:0] _0226_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3299" *)
  wire [37:0] _0227_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4029" *)
  wire [21:0] _0228_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4039" *)
  wire [21:0] _0229_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4049" *)
  wire [21:0] _0230_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4059" *)
  wire [21:0] _0231_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4069" *)
  wire [21:0] _0232_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4079" *)
  wire [21:0] _0233_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4089" *)
  wire [21:0] _0234_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4099" *)
  wire [21:0] _0235_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4109" *)
  wire [21:0] _0236_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4119" *)
  wire [21:0] _0237_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3309" *)
  wire [37:0] _0238_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4129" *)
  wire [21:0] _0239_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4139" *)
  wire [21:0] _0240_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4149" *)
  wire [21:0] _0241_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4159" *)
  wire [21:0] _0242_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4169" *)
  wire [21:0] _0243_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4179" *)
  wire [21:0] _0244_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4189" *)
  wire [21:0] _0245_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4199" *)
  wire [21:0] _0246_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4209" *)
  wire [21:0] _0247_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4219" *)
  wire [21:0] _0248_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3319" *)
  wire [37:0] _0249_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6429" *)
  wire [47:0] _0250_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6529" *)
  wire [47:0] _0251_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6539" *)
  wire [47:0] _0252_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6549" *)
  wire [47:0] _0253_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6559" *)
  wire [47:0] _0254_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6569" *)
  wire [47:0] _0255_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6579" *)
  wire [47:0] _0256_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6589" *)
  wire [47:0] _0257_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6599" *)
  wire [47:0] _0258_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6609" *)
  wire [47:0] _0259_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6619" *)
  wire [47:0] _0260_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6439" *)
  wire [47:0] _0261_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6629" *)
  wire [47:0] _0262_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6639" *)
  wire [47:0] _0263_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6649" *)
  wire [47:0] _0264_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6659" *)
  wire [47:0] _0265_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6669" *)
  wire [47:0] _0266_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6679" *)
  wire [47:0] _0267_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6689" *)
  wire [47:0] _0268_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6699" *)
  wire [47:0] _0269_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6709" *)
  wire [47:0] _0270_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6719" *)
  wire [47:0] _0271_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6449" *)
  wire [47:0] _0272_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6729" *)
  wire [47:0] _0273_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6739" *)
  wire [47:0] _0274_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6749" *)
  wire [47:0] _0275_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6759" *)
  wire [47:0] _0276_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6769" *)
  wire [47:0] _0277_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6779" *)
  wire [47:0] _0278_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6789" *)
  wire [47:0] _0279_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6799" *)
  wire [47:0] _0280_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6809" *)
  wire [47:0] _0281_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6819" *)
  wire [47:0] _0282_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6459" *)
  wire [47:0] _0283_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6829" *)
  wire [47:0] _0284_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6839" *)
  wire [47:0] _0285_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6849" *)
  wire [47:0] _0286_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6859" *)
  wire [47:0] _0287_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6869" *)
  wire [47:0] _0288_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6879" *)
  wire [47:0] _0289_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6889" *)
  wire [47:0] _0290_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6899" *)
  wire [47:0] _0291_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6909" *)
  wire [47:0] _0292_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6919" *)
  wire [47:0] _0293_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6469" *)
  wire [47:0] _0294_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6929" *)
  wire [47:0] _0295_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6939" *)
  wire [47:0] _0296_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6949" *)
  wire [47:0] _0297_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6959" *)
  wire [47:0] _0298_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6969" *)
  wire [47:0] _0299_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6979" *)
  wire [47:0] _0300_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6989" *)
  wire [47:0] _0301_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6999" *)
  wire [47:0] _0302_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7009" *)
  wire [47:0] _0303_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7019" *)
  wire [47:0] _0304_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6479" *)
  wire [47:0] _0305_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7029" *)
  wire [47:0] _0306_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7039" *)
  wire [47:0] _0307_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7049" *)
  wire [47:0] _0308_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7059" *)
  wire [47:0] _0309_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6489" *)
  wire [47:0] _0310_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6499" *)
  wire [47:0] _0311_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6509" *)
  wire [47:0] _0312_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6519" *)
  wire [47:0] _0313_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5149" *)
  wire [47:0] _0314_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6149" *)
  wire [33:0] _0315_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6159" *)
  wire [33:0] _0316_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6169" *)
  wire [33:0] _0317_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6179" *)
  wire [33:0] _0318_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6189" *)
  wire [33:0] _0319_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6199" *)
  wire [33:0] _0320_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6209" *)
  wire [33:0] _0321_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6219" *)
  wire [33:0] _0322_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6229" *)
  wire [33:0] _0323_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6239" *)
  wire [33:0] _0324_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5249" *)
  wire [47:0] _0325_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6249" *)
  wire [33:0] _0326_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6259" *)
  wire [33:0] _0327_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6269" *)
  wire [33:0] _0328_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6279" *)
  wire [33:0] _0329_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6289" *)
  wire [33:0] _0330_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6299" *)
  wire [33:0] _0331_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6309" *)
  wire [33:0] _0332_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6319" *)
  wire [33:0] _0333_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6329" *)
  wire [33:0] _0334_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6339" *)
  wire [33:0] _0335_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5259" *)
  wire [47:0] _0336_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6349" *)
  wire [33:0] _0337_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6359" *)
  wire [33:0] _0338_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6369" *)
  wire [33:0] _0339_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6379" *)
  wire [33:0] _0340_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6389" *)
  wire [33:0] _0341_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6399" *)
  wire [33:0] _0342_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6409" *)
  wire [33:0] _0343_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6419" *)
  wire [33:0] _0344_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5269" *)
  wire [47:0] _0345_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5279" *)
  wire [47:0] _0346_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5289" *)
  wire [47:0] _0347_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5299" *)
  wire [47:0] _0348_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5309" *)
  wire [47:0] _0349_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5319" *)
  wire [47:0] _0350_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5329" *)
  wire [47:0] _0351_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5339" *)
  wire [47:0] _0352_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5159" *)
  wire [47:0] _0353_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5349" *)
  wire [47:0] _0354_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5359" *)
  wire [47:0] _0355_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5369" *)
  wire [47:0] _0356_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5379" *)
  wire [47:0] _0357_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5389" *)
  wire [47:0] _0358_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5399" *)
  wire [47:0] _0359_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5409" *)
  wire [47:0] _0360_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5419" *)
  wire [47:0] _0361_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5429" *)
  wire [47:0] _0362_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5439" *)
  wire [47:0] _0363_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5169" *)
  wire [47:0] _0364_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5449" *)
  wire [47:0] _0365_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5459" *)
  wire [47:0] _0366_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5469" *)
  wire [47:0] _0367_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5479" *)
  wire [47:0] _0368_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5489" *)
  wire [47:0] _0369_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5499" *)
  wire [47:0] _0370_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5509" *)
  wire [47:0] _0371_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5519" *)
  wire [47:0] _0372_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5529" *)
  wire [47:0] _0373_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5539" *)
  wire [47:0] _0374_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5179" *)
  wire [47:0] _0375_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5549" *)
  wire [47:0] _0376_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5559" *)
  wire [47:0] _0377_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5569" *)
  wire [47:0] _0378_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5579" *)
  wire [47:0] _0379_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5589" *)
  wire [47:0] _0380_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5599" *)
  wire [47:0] _0381_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5609" *)
  wire [47:0] _0382_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5619" *)
  wire [47:0] _0383_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5629" *)
  wire [47:0] _0384_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5639" *)
  wire [47:0] _0385_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5189" *)
  wire [47:0] _0386_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5649" *)
  wire [47:0] _0387_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5659" *)
  wire [47:0] _0388_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5669" *)
  wire [47:0] _0389_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5679" *)
  wire [47:0] _0390_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5689" *)
  wire [47:0] _0391_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5699" *)
  wire [47:0] _0392_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5709" *)
  wire [47:0] _0393_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5719" *)
  wire [47:0] _0394_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5729" *)
  wire [47:0] _0395_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5739" *)
  wire [47:0] _0396_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5199" *)
  wire [47:0] _0397_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5749" *)
  wire [47:0] _0398_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5759" *)
  wire [47:0] _0399_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5769" *)
  wire [47:0] _0400_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5779" *)
  wire [47:0] _0401_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5789" *)
  wire [33:0] _0402_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5799" *)
  wire [33:0] _0403_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5809" *)
  wire [33:0] _0404_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5819" *)
  wire [33:0] _0405_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5829" *)
  wire [33:0] _0406_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5839" *)
  wire [33:0] _0407_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5209" *)
  wire [47:0] _0408_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5849" *)
  wire [33:0] _0409_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5859" *)
  wire [33:0] _0410_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5869" *)
  wire [33:0] _0411_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5879" *)
  wire [33:0] _0412_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5889" *)
  wire [33:0] _0413_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5899" *)
  wire [33:0] _0414_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5909" *)
  wire [33:0] _0415_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5919" *)
  wire [33:0] _0416_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5929" *)
  wire [33:0] _0417_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5939" *)
  wire [33:0] _0418_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5219" *)
  wire [47:0] _0419_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5949" *)
  wire [33:0] _0420_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5959" *)
  wire [33:0] _0421_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5969" *)
  wire [33:0] _0422_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5979" *)
  wire [33:0] _0423_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5989" *)
  wire [33:0] _0424_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5999" *)
  wire [33:0] _0425_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6009" *)
  wire [33:0] _0426_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6019" *)
  wire [33:0] _0427_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6029" *)
  wire [33:0] _0428_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6039" *)
  wire [33:0] _0429_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5229" *)
  wire [47:0] _0430_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6049" *)
  wire [33:0] _0431_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6059" *)
  wire [33:0] _0432_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6069" *)
  wire [33:0] _0433_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6079" *)
  wire [33:0] _0434_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6089" *)
  wire [33:0] _0435_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6099" *)
  wire [33:0] _0436_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6109" *)
  wire [33:0] _0437_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6119" *)
  wire [33:0] _0438_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6129" *)
  wire [33:0] _0439_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6139" *)
  wire [33:0] _0440_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5239" *)
  wire [47:0] _0441_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7571" *)
  wire [63:0] _0442_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7510" *)
  wire [127:0] _0443_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7449" *)
  wire [63:0] _0444_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7388" *)
  wire [127:0] _0445_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7266" *)
  wire _0446_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10974" *)
  wire _0447_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11164" *)
  wire _0448_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11354" *)
  wire _0449_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11544" *)
  wire _0450_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7076" *)
  wire [7:0] _0451_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10520" *)
  wire [7:0] _0452_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10649" *)
  wire [7:0] _0453_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10778" *)
  wire [7:0] _0454_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12989" *)
  wire [511:0] _0455_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12999" *)
  wire [511:0] _0456_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13009" *)
  wire [511:0] _0457_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13019" *)
  wire [511:0] _0458_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13029" *)
  wire [511:0] _0459_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13039" *)
  wire [511:0] _0460_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13049" *)
  wire [511:0] _0461_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13059" *)
  wire [511:0] _0462_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13198" *)
  wire _0463_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13076" *)
  wire [7:0] _0464_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13336" *)
  wire [127:0] _0465_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13275" *)
  wire _0466_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13137" *)
  wire _0467_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13421" *)
  wire [31:0] _0468_;
  wire [1:0] _0469_;
  wire [2:0] _0470_;
  wire [3:0] _0471_;
  wire [4:0] _0472_;
  wire [5:0] _0473_;
  wire [6:0] _0474_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0475_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0476_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0477_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0478_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0479_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0480_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0481_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0482_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0483_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0484_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0485_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0486_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0487_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0488_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0489_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0490_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0491_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0492_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0493_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0494_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0495_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0496_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0497_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0498_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0499_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0500_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0501_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0502_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0503_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0504_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0505_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0506_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0507_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0508_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0509_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0510_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0511_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0512_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0513_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0514_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0515_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0516_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0517_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0518_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0519_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0520_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0521_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0522_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0523_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0524_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0525_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0526_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0527_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0528_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0529_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0530_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0531_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0532_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0533_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0534_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0535_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0536_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0537_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0538_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0539_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0540_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0541_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0542_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0543_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0544_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0545_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0546_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0547_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0548_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0549_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0550_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0551_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0552_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0553_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0554_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0555_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0556_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0557_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0558_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0559_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0560_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0561_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0562_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0563_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0564_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0565_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0566_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0567_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0568_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0569_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0570_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0571_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0572_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0573_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0574_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0575_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0576_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0577_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0578_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0579_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0580_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0581_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0582_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0583_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0584_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0585_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0586_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0587_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0588_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0589_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0590_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0591_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0592_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0593_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *)
  wire [7:0] _0594_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10902" *)
  wire [7:0] _0595_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10903" *)
  wire [7:0] _0596_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10904" *)
  wire [4:0] _0597_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10905" *)
  wire [4:0] _0598_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11666" *)
  wire _0599_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11667" *)
  wire _0600_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11668" *)
  wire [7:0] _0601_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11669" *)
  wire [7:0] _0602_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11670" *)
  wire _0603_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11671" *)
  wire _0604_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11672" *)
  wire _0605_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11673" *)
  wire _0606_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11741" *)
  wire [47:0] _0607_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11742" *)
  wire [47:0] _0608_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11743" *)
  wire [47:0] _0609_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11744" *)
  wire [47:0] _0610_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11745" *)
  wire [47:0] _0611_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11746" *)
  wire [47:0] _0612_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11747" *)
  wire [47:0] _0613_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11748" *)
  wire [47:0] _0614_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11749" *)
  wire [47:0] _0615_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11750" *)
  wire [47:0] _0616_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11751" *)
  wire [47:0] _0617_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11752" *)
  wire [47:0] _0618_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11753" *)
  wire [47:0] _0619_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11754" *)
  wire [47:0] _0620_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11755" *)
  wire [47:0] _0621_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11756" *)
  wire [47:0] _0622_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11757" *)
  wire [47:0] _0623_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11758" *)
  wire [47:0] _0624_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11759" *)
  wire [47:0] _0625_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11760" *)
  wire [47:0] _0626_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11761" *)
  wire [47:0] _0627_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11762" *)
  wire [47:0] _0628_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11763" *)
  wire [47:0] _0629_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11764" *)
  wire [47:0] _0630_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11765" *)
  wire [47:0] _0631_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11766" *)
  wire [47:0] _0632_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11767" *)
  wire [47:0] _0633_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11768" *)
  wire [47:0] _0634_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11769" *)
  wire [47:0] _0635_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11770" *)
  wire [47:0] _0636_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11771" *)
  wire [47:0] _0637_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11772" *)
  wire [47:0] _0638_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11773" *)
  wire [47:0] _0639_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11774" *)
  wire [47:0] _0640_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11775" *)
  wire [47:0] _0641_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11776" *)
  wire [47:0] _0642_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11777" *)
  wire [47:0] _0643_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11778" *)
  wire [47:0] _0644_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11779" *)
  wire [47:0] _0645_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11780" *)
  wire [47:0] _0646_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11781" *)
  wire [47:0] _0647_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11782" *)
  wire [47:0] _0648_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11783" *)
  wire [47:0] _0649_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11784" *)
  wire [47:0] _0650_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11785" *)
  wire [47:0] _0651_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11786" *)
  wire [47:0] _0652_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11787" *)
  wire [47:0] _0653_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11788" *)
  wire [47:0] _0654_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11789" *)
  wire [47:0] _0655_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11790" *)
  wire [47:0] _0656_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11791" *)
  wire [47:0] _0657_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11792" *)
  wire [47:0] _0658_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11793" *)
  wire [47:0] _0659_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11794" *)
  wire [47:0] _0660_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11795" *)
  wire [47:0] _0661_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11796" *)
  wire [47:0] _0662_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11797" *)
  wire [47:0] _0663_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11798" *)
  wire [47:0] _0664_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11799" *)
  wire [47:0] _0665_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11800" *)
  wire [47:0] _0666_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11801" *)
  wire [47:0] _0667_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11802" *)
  wire [47:0] _0668_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11803" *)
  wire [47:0] _0669_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11804" *)
  wire [47:0] _0670_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11805" *)
  wire [47:0] _0671_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11806" *)
  wire [47:0] _0672_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11807" *)
  wire [47:0] _0673_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11808" *)
  wire [47:0] _0674_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11809" *)
  wire [47:0] _0675_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11810" *)
  wire [47:0] _0676_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11811" *)
  wire [47:0] _0677_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11812" *)
  wire [47:0] _0678_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11813" *)
  wire [47:0] _0679_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11814" *)
  wire [47:0] _0680_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11815" *)
  wire [47:0] _0681_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11816" *)
  wire [47:0] _0682_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11817" *)
  wire [47:0] _0683_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11818" *)
  wire [47:0] _0684_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11819" *)
  wire [47:0] _0685_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11820" *)
  wire [47:0] _0686_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11821" *)
  wire [47:0] _0687_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11822" *)
  wire [47:0] _0688_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11823" *)
  wire [47:0] _0689_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11824" *)
  wire [47:0] _0690_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11825" *)
  wire [47:0] _0691_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11826" *)
  wire [47:0] _0692_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11827" *)
  wire [47:0] _0693_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11828" *)
  wire [47:0] _0694_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11829" *)
  wire [47:0] _0695_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11830" *)
  wire [47:0] _0696_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11831" *)
  wire [47:0] _0697_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11832" *)
  wire [47:0] _0698_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11833" *)
  wire [47:0] _0699_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11834" *)
  wire [47:0] _0700_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11835" *)
  wire [47:0] _0701_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11836" *)
  wire [47:0] _0702_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11837" *)
  wire [47:0] _0703_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11838" *)
  wire [47:0] _0704_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11839" *)
  wire [47:0] _0705_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11840" *)
  wire [47:0] _0706_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11841" *)
  wire [47:0] _0707_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11842" *)
  wire [47:0] _0708_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11843" *)
  wire [47:0] _0709_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11844" *)
  wire [47:0] _0710_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11845" *)
  wire [47:0] _0711_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11846" *)
  wire [47:0] _0712_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11847" *)
  wire [47:0] _0713_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11848" *)
  wire [47:0] _0714_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11849" *)
  wire [47:0] _0715_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11850" *)
  wire [47:0] _0716_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11851" *)
  wire [47:0] _0717_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11852" *)
  wire [47:0] _0718_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11853" *)
  wire [47:0] _0719_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11854" *)
  wire [47:0] _0720_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11855" *)
  wire [47:0] _0721_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11856" *)
  wire [47:0] _0722_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11857" *)
  wire [47:0] _0723_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11858" *)
  wire [47:0] _0724_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11859" *)
  wire [47:0] _0725_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11860" *)
  wire [47:0] _0726_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11861" *)
  wire [47:0] _0727_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11862" *)
  wire [47:0] _0728_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11863" *)
  wire [47:0] _0729_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11864" *)
  wire [47:0] _0730_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11865" *)
  wire [47:0] _0731_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11866" *)
  wire [47:0] _0732_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11867" *)
  wire [47:0] _0733_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11868" *)
  wire [47:0] _0734_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11933" *)
  wire [31:0] _0735_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11934" *)
  wire [31:0] _0736_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11935" *)
  wire [31:0] _0737_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11936" *)
  wire [31:0] _0738_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11937" *)
  wire [31:0] _0739_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11938" *)
  wire [31:0] _0740_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11939" *)
  wire [31:0] _0741_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11940" *)
  wire [31:0] _0742_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11941" *)
  wire [31:0] _0743_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11942" *)
  wire [31:0] _0744_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11943" *)
  wire [31:0] _0745_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11944" *)
  wire [31:0] _0746_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11945" *)
  wire [31:0] _0747_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11946" *)
  wire [31:0] _0748_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11947" *)
  wire [31:0] _0749_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11948" *)
  wire [31:0] _0750_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11949" *)
  wire [31:0] _0751_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11950" *)
  wire [31:0] _0752_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11951" *)
  wire [31:0] _0753_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11952" *)
  wire [31:0] _0754_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11953" *)
  wire [31:0] _0755_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11954" *)
  wire [31:0] _0756_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11955" *)
  wire [31:0] _0757_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11956" *)
  wire [31:0] _0758_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11957" *)
  wire [31:0] _0759_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11958" *)
  wire [31:0] _0760_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11959" *)
  wire [31:0] _0761_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11960" *)
  wire [31:0] _0762_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11961" *)
  wire [31:0] _0763_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11962" *)
  wire [31:0] _0764_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11963" *)
  wire [31:0] _0765_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11964" *)
  wire [31:0] _0766_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11965" *)
  wire [31:0] _0767_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11966" *)
  wire [31:0] _0768_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11967" *)
  wire [31:0] _0769_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11968" *)
  wire [31:0] _0770_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11969" *)
  wire [31:0] _0771_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11970" *)
  wire [31:0] _0772_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11971" *)
  wire [31:0] _0773_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11972" *)
  wire [31:0] _0774_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11973" *)
  wire [31:0] _0775_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11974" *)
  wire [31:0] _0776_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11975" *)
  wire [31:0] _0777_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11976" *)
  wire [31:0] _0778_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11977" *)
  wire [31:0] _0779_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11978" *)
  wire [31:0] _0780_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11979" *)
  wire [31:0] _0781_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11980" *)
  wire [31:0] _0782_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11981" *)
  wire [31:0] _0783_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11982" *)
  wire [31:0] _0784_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11983" *)
  wire [31:0] _0785_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11984" *)
  wire [31:0] _0786_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11985" *)
  wire [31:0] _0787_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11986" *)
  wire [31:0] _0788_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11987" *)
  wire [31:0] _0789_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11988" *)
  wire [31:0] _0790_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11989" *)
  wire [31:0] _0791_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11990" *)
  wire [31:0] _0792_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11991" *)
  wire [31:0] _0793_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11992" *)
  wire [31:0] _0794_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11993" *)
  wire [31:0] _0795_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11994" *)
  wire [31:0] _0796_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11995" *)
  wire [31:0] _0797_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11996" *)
  wire [31:0] _0798_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11997" *)
  wire [31:0] _0799_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11998" *)
  wire [31:0] _0800_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11999" *)
  wire [31:0] _0801_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12000" *)
  wire [31:0] _0802_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12001" *)
  wire [31:0] _0803_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12002" *)
  wire [31:0] _0804_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12003" *)
  wire [31:0] _0805_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12004" *)
  wire [31:0] _0806_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12005" *)
  wire [31:0] _0807_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12006" *)
  wire [31:0] _0808_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12007" *)
  wire [31:0] _0809_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12008" *)
  wire [31:0] _0810_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12009" *)
  wire [31:0] _0811_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12010" *)
  wire [31:0] _0812_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12011" *)
  wire [31:0] _0813_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12012" *)
  wire [31:0] _0814_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12013" *)
  wire [31:0] _0815_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12014" *)
  wire [31:0] _0816_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12015" *)
  wire [31:0] _0817_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12016" *)
  wire [31:0] _0818_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12017" *)
  wire [31:0] _0819_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12018" *)
  wire [31:0] _0820_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12019" *)
  wire [31:0] _0821_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12020" *)
  wire [31:0] _0822_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12021" *)
  wire [31:0] _0823_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12022" *)
  wire [31:0] _0824_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12023" *)
  wire [31:0] _0825_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12024" *)
  wire [31:0] _0826_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12025" *)
  wire [31:0] _0827_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12026" *)
  wire [31:0] _0828_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12027" *)
  wire [31:0] _0829_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12028" *)
  wire [31:0] _0830_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12029" *)
  wire [31:0] _0831_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12030" *)
  wire [31:0] _0832_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12031" *)
  wire [31:0] _0833_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12032" *)
  wire [31:0] _0834_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12033" *)
  wire [31:0] _0835_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12034" *)
  wire [31:0] _0836_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12035" *)
  wire [31:0] _0837_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12036" *)
  wire [31:0] _0838_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12037" *)
  wire [31:0] _0839_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12038" *)
  wire [31:0] _0840_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12039" *)
  wire [31:0] _0841_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12040" *)
  wire [31:0] _0842_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12041" *)
  wire [31:0] _0843_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12042" *)
  wire [31:0] _0844_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12043" *)
  wire [31:0] _0845_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12044" *)
  wire [31:0] _0846_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12045" *)
  wire [31:0] _0847_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12046" *)
  wire [31:0] _0848_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12047" *)
  wire [31:0] _0849_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12048" *)
  wire [31:0] _0850_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12049" *)
  wire [31:0] _0851_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12050" *)
  wire [31:0] _0852_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12051" *)
  wire [31:0] _0853_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12052" *)
  wire [31:0] _0854_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12053" *)
  wire [31:0] _0855_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12054" *)
  wire [31:0] _0856_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12055" *)
  wire [31:0] _0857_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12056" *)
  wire [31:0] _0858_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12057" *)
  wire [31:0] _0859_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12058" *)
  wire [31:0] _0860_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12059" *)
  wire [31:0] _0861_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12060" *)
  wire [31:0] _0862_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13267" *)
  wire _0863_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2280" *)
  wire _0864_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2300" *)
  wire _0865_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2320" *)
  wire _0866_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2340" *)
  wire _0867_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2360" *)
  wire _0868_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2380" *)
  wire _0869_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2400" *)
  wire _0870_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2420" *)
  wire _0871_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2440" *)
  wire _0872_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2460" *)
  wire _0873_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2480" *)
  wire _0874_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2500" *)
  wire _0875_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2520" *)
  wire _0876_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2540" *)
  wire _0877_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2560" *)
  wire _0878_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2580" *)
  wire _0879_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3138" *)
  wire [767:0] _0880_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3139" *)
  wire [767:0] _0881_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3140" *)
  wire [767:0] _0882_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3141" *)
  wire [767:0] _0883_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3162" *)
  wire [543:0] _0884_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3163" *)
  wire [543:0] _0885_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3164" *)
  wire [543:0] _0886_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3165" *)
  wire [543:0] _0887_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10524" *)
  wire _0888_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10653" *)
  wire _0889_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10782" *)
  wire _0890_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10917" *)
  wire _0891_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11107" *)
  wire _0892_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11297" *)
  wire _0893_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11487" *)
  wire _0894_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12588" *)
  wire _0895_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2616" *)
  wire _0896_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7080" *)
  wire _0897_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13267" *)
  wire _0898_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3205" *)
  wire _0899_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3205" *)
  wire _0900_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3216" *)
  wire _0901_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13420" *)
  wire _0902_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3139" *)
  wire [767:0] _0903_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3140" *)
  wire [767:0] _0904_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3163" *)
  wire [543:0] _0905_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3164" *)
  wire [543:0] _0906_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3205" *)
  wire _0907_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3216" *)
  wire _0908_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13420" *)
  wire _0909_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13419" *)
  wire [31:0] _0910_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *)
  wire [7:0] _0911_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *)
  wire [7:0] _0912_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *)
  wire [7:0] _0913_;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1606" *)
  wire [47:0] abuf_in_data_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1607" *)
  wire [47:0] abuf_in_data_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1608" *)
  wire [47:0] abuf_in_data_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1609" *)
  wire [33:0] abuf_in_data_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1610" *)
  wire [33:0] abuf_in_data_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1611" *)
  wire [33:0] abuf_in_data_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1612" *)
  wire [33:0] abuf_in_data_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1613" *)
  wire [33:0] abuf_in_data_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1614" *)
  wire [33:0] abuf_in_data_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1615" *)
  wire [33:0] abuf_in_data_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1616" *)
  wire [33:0] abuf_in_data_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1617" *)
  wire [33:0] abuf_in_data_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1618" *)
  wire [33:0] abuf_in_data_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1619" *)
  wire [47:0] abuf_in_data_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1620" *)
  wire [33:0] abuf_in_data_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1621" *)
  wire [33:0] abuf_in_data_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1622" *)
  wire [33:0] abuf_in_data_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1623" *)
  wire [33:0] abuf_in_data_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1624" *)
  wire [33:0] abuf_in_data_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1625" *)
  wire [33:0] abuf_in_data_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1626" *)
  wire [33:0] abuf_in_data_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1627" *)
  wire [33:0] abuf_in_data_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1628" *)
  wire [33:0] abuf_in_data_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1629" *)
  wire [33:0] abuf_in_data_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1630" *)
  wire [47:0] abuf_in_data_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1631" *)
  wire [33:0] abuf_in_data_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1632" *)
  wire [33:0] abuf_in_data_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1633" *)
  wire [33:0] abuf_in_data_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1634" *)
  wire [33:0] abuf_in_data_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1635" *)
  wire [33:0] abuf_in_data_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1636" *)
  wire [33:0] abuf_in_data_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1637" *)
  wire [33:0] abuf_in_data_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1638" *)
  wire [33:0] abuf_in_data_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1639" *)
  wire [47:0] abuf_in_data_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1640" *)
  wire [47:0] abuf_in_data_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1641" *)
  wire [47:0] abuf_in_data_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1642" *)
  wire [47:0] abuf_in_data_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1643" *)
  wire [47:0] abuf_in_data_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1644" *)
  wire [47:0] abuf_in_data_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1645" *)
  wire [47:0] abuf_in_data_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1646" *)
  wire [47:0] abuf_in_data_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1647" *)
  wire [47:0] abuf_in_data_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1648" *)
  wire [47:0] abuf_in_data_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1649" *)
  wire [47:0] abuf_in_data_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1650" *)
  wire [47:0] abuf_in_data_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1651" *)
  wire [47:0] abuf_in_data_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1652" *)
  wire [47:0] abuf_in_data_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1653" *)
  wire [47:0] abuf_in_data_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1654" *)
  wire [47:0] abuf_in_data_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1655" *)
  wire [47:0] abuf_in_data_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1656" *)
  wire [47:0] abuf_in_data_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1657" *)
  wire [47:0] abuf_in_data_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1658" *)
  wire [47:0] abuf_in_data_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1659" *)
  wire [47:0] abuf_in_data_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1660" *)
  wire [47:0] abuf_in_data_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1661" *)
  wire [47:0] abuf_in_data_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1662" *)
  wire [47:0] abuf_in_data_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1663" *)
  wire [47:0] abuf_in_data_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1664" *)
  wire [47:0] abuf_in_data_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1665" *)
  wire [47:0] abuf_in_data_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1666" *)
  wire [47:0] abuf_in_data_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1667" *)
  wire [47:0] abuf_in_data_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1668" *)
  wire [47:0] abuf_in_data_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1669" *)
  wire [47:0] abuf_in_data_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1670" *)
  wire [47:0] abuf_in_data_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1671" *)
  wire [47:0] abuf_in_data_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1672" *)
  wire [47:0] abuf_in_data_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1673" *)
  wire [47:0] abuf_in_data_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1674" *)
  wire [47:0] abuf_in_data_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1675" *)
  wire [47:0] abuf_in_data_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1676" *)
  wire [47:0] abuf_in_data_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1677" *)
  wire [47:0] abuf_in_data_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1678" *)
  wire [47:0] abuf_in_data_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1679" *)
  wire [47:0] abuf_in_data_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1680" *)
  wire [47:0] abuf_in_data_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1681" *)
  wire [47:0] abuf_in_data_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1682" *)
  wire [47:0] abuf_in_data_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1683" *)
  wire [47:0] abuf_in_data_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1684" *)
  wire [47:0] abuf_in_data_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1685" *)
  wire [47:0] abuf_in_data_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1686" *)
  wire [47:0] abuf_in_data_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1687" *)
  wire [47:0] abuf_in_data_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1688" *)
  wire [47:0] abuf_in_data_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1689" *)
  wire [47:0] abuf_in_data_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1690" *)
  wire [47:0] abuf_in_data_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1691" *)
  wire [47:0] abuf_in_data_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1692" *)
  wire [47:0] abuf_in_data_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1693" *)
  wire [47:0] abuf_in_data_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1694" *)
  wire [47:0] abuf_in_data_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1695" *)
  wire [33:0] abuf_in_data_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1696" *)
  wire [33:0] abuf_in_data_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1697" *)
  wire [33:0] abuf_in_data_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1698" *)
  wire [33:0] abuf_in_data_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1699" *)
  wire [33:0] abuf_in_data_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1700" *)
  wire [33:0] abuf_in_data_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1701" *)
  wire [47:0] abuf_in_data_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1702" *)
  wire [33:0] abuf_in_data_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1703" *)
  wire [33:0] abuf_in_data_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1704" *)
  wire [33:0] abuf_in_data_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1705" *)
  wire [33:0] abuf_in_data_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1706" *)
  wire [33:0] abuf_in_data_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1707" *)
  wire [33:0] abuf_in_data_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1708" *)
  wire [33:0] abuf_in_data_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1709" *)
  wire [33:0] abuf_in_data_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1710" *)
  wire [33:0] abuf_in_data_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1711" *)
  wire [33:0] abuf_in_data_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1712" *)
  wire [47:0] abuf_in_data_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1713" *)
  wire [33:0] abuf_in_data_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1714" *)
  wire [33:0] abuf_in_data_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1715" *)
  wire [33:0] abuf_in_data_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1716" *)
  wire [33:0] abuf_in_data_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1717" *)
  wire [33:0] abuf_in_data_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1718" *)
  wire [33:0] abuf_in_data_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1719" *)
  wire [33:0] abuf_in_data_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1720" *)
  wire [33:0] abuf_in_data_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1721" *)
  wire [33:0] abuf_in_data_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1722" *)
  wire [33:0] abuf_in_data_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1723" *)
  wire [47:0] abuf_in_data_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1724" *)
  wire [33:0] abuf_in_data_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1725" *)
  wire [33:0] abuf_in_data_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1726" *)
  wire [33:0] abuf_in_data_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1727" *)
  wire [33:0] abuf_in_data_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1728" *)
  wire [33:0] abuf_in_data_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1729" *)
  wire [33:0] abuf_in_data_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1730" *)
  wire [33:0] abuf_in_data_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1731" *)
  wire [33:0] abuf_in_data_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1732" *)
  wire [33:0] abuf_in_data_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1733" *)
  wire [33:0] abuf_in_data_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:84" *)
  input [767:0] abuf_rd_data_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1734" *)
  wire [767:0] abuf_rd_data_0_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:85" *)
  input [767:0] abuf_rd_data_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1735" *)
  wire [767:0] abuf_rd_data_1_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:86" *)
  input [767:0] abuf_rd_data_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1736" *)
  wire [767:0] abuf_rd_data_2_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:87" *)
  input [767:0] abuf_rd_data_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1737" *)
  wire [767:0] abuf_rd_data_3_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:88" *)
  input [543:0] abuf_rd_data_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1738" *)
  wire [543:0] abuf_rd_data_4_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:89" *)
  input [543:0] abuf_rd_data_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1739" *)
  wire [543:0] abuf_rd_data_5_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:90" *)
  input [543:0] abuf_rd_data_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1740" *)
  wire [543:0] abuf_rd_data_6_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:91" *)
  input [543:0] abuf_rd_data_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1741" *)
  wire [543:0] abuf_rd_data_7_sft;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:123" *)
  output [4:0] abuf_wr_addr;
  reg [4:0] abuf_wr_addr;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:124" *)
  output [767:0] abuf_wr_data_0;
  reg [767:0] abuf_wr_data_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1744" *)
  wire [767:0] abuf_wr_data_0_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:125" *)
  output [767:0] abuf_wr_data_1;
  reg [767:0] abuf_wr_data_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1746" *)
  wire [767:0] abuf_wr_data_1_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:126" *)
  output [767:0] abuf_wr_data_2;
  reg [767:0] abuf_wr_data_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1748" *)
  wire [767:0] abuf_wr_data_2_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:127" *)
  output [767:0] abuf_wr_data_3;
  reg [767:0] abuf_wr_data_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1750" *)
  wire [767:0] abuf_wr_data_3_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:128" *)
  output [543:0] abuf_wr_data_4;
  reg [543:0] abuf_wr_data_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1752" *)
  wire [543:0] abuf_wr_data_4_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:129" *)
  output [543:0] abuf_wr_data_5;
  reg [543:0] abuf_wr_data_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1754" *)
  wire [543:0] abuf_wr_data_5_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:130" *)
  output [543:0] abuf_wr_data_6;
  reg [543:0] abuf_wr_data_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1756" *)
  wire [543:0] abuf_wr_data_6_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:131" *)
  output [543:0] abuf_wr_data_7;
  reg [543:0] abuf_wr_data_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1758" *)
  wire [543:0] abuf_wr_data_7_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:145" *)
  wire [47:0] abuf_wr_elem_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:146" *)
  wire [47:0] abuf_wr_elem_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:147" *)
  wire [47:0] abuf_wr_elem_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:148" *)
  wire [33:0] abuf_wr_elem_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:149" *)
  wire [33:0] abuf_wr_elem_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:150" *)
  wire [33:0] abuf_wr_elem_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:151" *)
  wire [33:0] abuf_wr_elem_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:152" *)
  wire [33:0] abuf_wr_elem_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:153" *)
  wire [33:0] abuf_wr_elem_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:154" *)
  wire [33:0] abuf_wr_elem_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:155" *)
  wire [33:0] abuf_wr_elem_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:156" *)
  wire [33:0] abuf_wr_elem_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:157" *)
  wire [33:0] abuf_wr_elem_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:158" *)
  wire [47:0] abuf_wr_elem_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:159" *)
  wire [33:0] abuf_wr_elem_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:160" *)
  wire [33:0] abuf_wr_elem_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:161" *)
  wire [33:0] abuf_wr_elem_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:162" *)
  wire [33:0] abuf_wr_elem_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:163" *)
  wire [33:0] abuf_wr_elem_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:164" *)
  wire [33:0] abuf_wr_elem_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:165" *)
  wire [33:0] abuf_wr_elem_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:166" *)
  wire [33:0] abuf_wr_elem_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:167" *)
  wire [33:0] abuf_wr_elem_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:168" *)
  wire [33:0] abuf_wr_elem_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:169" *)
  wire [47:0] abuf_wr_elem_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:170" *)
  wire [33:0] abuf_wr_elem_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:171" *)
  wire [33:0] abuf_wr_elem_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:172" *)
  wire [33:0] abuf_wr_elem_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:173" *)
  wire [33:0] abuf_wr_elem_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:174" *)
  wire [33:0] abuf_wr_elem_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:175" *)
  wire [33:0] abuf_wr_elem_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:176" *)
  wire [33:0] abuf_wr_elem_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:177" *)
  wire [33:0] abuf_wr_elem_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:178" *)
  wire [47:0] abuf_wr_elem_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:179" *)
  wire [47:0] abuf_wr_elem_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:180" *)
  wire [47:0] abuf_wr_elem_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:181" *)
  wire [47:0] abuf_wr_elem_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:182" *)
  wire [47:0] abuf_wr_elem_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:183" *)
  wire [47:0] abuf_wr_elem_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:184" *)
  wire [47:0] abuf_wr_elem_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:185" *)
  wire [47:0] abuf_wr_elem_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:186" *)
  wire [47:0] abuf_wr_elem_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:187" *)
  wire [47:0] abuf_wr_elem_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:188" *)
  wire [47:0] abuf_wr_elem_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:189" *)
  wire [47:0] abuf_wr_elem_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:190" *)
  wire [47:0] abuf_wr_elem_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:191" *)
  wire [47:0] abuf_wr_elem_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:192" *)
  wire [47:0] abuf_wr_elem_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:193" *)
  wire [47:0] abuf_wr_elem_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:194" *)
  wire [47:0] abuf_wr_elem_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:195" *)
  wire [47:0] abuf_wr_elem_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:196" *)
  wire [47:0] abuf_wr_elem_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:197" *)
  wire [47:0] abuf_wr_elem_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:198" *)
  wire [47:0] abuf_wr_elem_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:199" *)
  wire [47:0] abuf_wr_elem_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:200" *)
  wire [47:0] abuf_wr_elem_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:201" *)
  wire [47:0] abuf_wr_elem_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:202" *)
  wire [47:0] abuf_wr_elem_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:203" *)
  wire [47:0] abuf_wr_elem_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:204" *)
  wire [47:0] abuf_wr_elem_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:205" *)
  wire [47:0] abuf_wr_elem_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:206" *)
  wire [47:0] abuf_wr_elem_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:207" *)
  wire [47:0] abuf_wr_elem_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:208" *)
  wire [47:0] abuf_wr_elem_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:209" *)
  wire [47:0] abuf_wr_elem_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:210" *)
  wire [47:0] abuf_wr_elem_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:211" *)
  wire [47:0] abuf_wr_elem_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:212" *)
  wire [47:0] abuf_wr_elem_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:213" *)
  wire [47:0] abuf_wr_elem_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:214" *)
  wire [47:0] abuf_wr_elem_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:215" *)
  wire [47:0] abuf_wr_elem_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:216" *)
  wire [47:0] abuf_wr_elem_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:217" *)
  wire [47:0] abuf_wr_elem_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:218" *)
  wire [47:0] abuf_wr_elem_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:219" *)
  wire [47:0] abuf_wr_elem_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:220" *)
  wire [47:0] abuf_wr_elem_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:221" *)
  wire [47:0] abuf_wr_elem_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:222" *)
  wire [47:0] abuf_wr_elem_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:223" *)
  wire [47:0] abuf_wr_elem_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:224" *)
  wire [47:0] abuf_wr_elem_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:225" *)
  wire [47:0] abuf_wr_elem_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:226" *)
  wire [47:0] abuf_wr_elem_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:227" *)
  wire [47:0] abuf_wr_elem_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:228" *)
  wire [47:0] abuf_wr_elem_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:229" *)
  wire [47:0] abuf_wr_elem_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:230" *)
  wire [47:0] abuf_wr_elem_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:231" *)
  wire [47:0] abuf_wr_elem_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:232" *)
  wire [47:0] abuf_wr_elem_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:233" *)
  wire [47:0] abuf_wr_elem_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:234" *)
  wire [33:0] abuf_wr_elem_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:235" *)
  wire [33:0] abuf_wr_elem_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:236" *)
  wire [33:0] abuf_wr_elem_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:237" *)
  wire [33:0] abuf_wr_elem_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:238" *)
  wire [33:0] abuf_wr_elem_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:239" *)
  wire [33:0] abuf_wr_elem_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:240" *)
  wire [47:0] abuf_wr_elem_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:241" *)
  wire [33:0] abuf_wr_elem_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:242" *)
  wire [33:0] abuf_wr_elem_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:243" *)
  wire [33:0] abuf_wr_elem_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:244" *)
  wire [33:0] abuf_wr_elem_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:245" *)
  wire [33:0] abuf_wr_elem_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:246" *)
  wire [33:0] abuf_wr_elem_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:247" *)
  wire [33:0] abuf_wr_elem_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:248" *)
  wire [33:0] abuf_wr_elem_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:249" *)
  wire [33:0] abuf_wr_elem_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:250" *)
  wire [33:0] abuf_wr_elem_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:251" *)
  wire [47:0] abuf_wr_elem_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:252" *)
  wire [33:0] abuf_wr_elem_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:253" *)
  wire [33:0] abuf_wr_elem_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:254" *)
  wire [33:0] abuf_wr_elem_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:255" *)
  wire [33:0] abuf_wr_elem_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:256" *)
  wire [33:0] abuf_wr_elem_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:257" *)
  wire [33:0] abuf_wr_elem_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:258" *)
  wire [33:0] abuf_wr_elem_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:259" *)
  wire [33:0] abuf_wr_elem_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:260" *)
  wire [33:0] abuf_wr_elem_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:261" *)
  wire [33:0] abuf_wr_elem_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:262" *)
  wire [47:0] abuf_wr_elem_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:263" *)
  wire [33:0] abuf_wr_elem_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:264" *)
  wire [33:0] abuf_wr_elem_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:265" *)
  wire [33:0] abuf_wr_elem_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:266" *)
  wire [33:0] abuf_wr_elem_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:267" *)
  wire [33:0] abuf_wr_elem_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:268" *)
  wire [33:0] abuf_wr_elem_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:269" *)
  wire [33:0] abuf_wr_elem_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:270" *)
  wire [33:0] abuf_wr_elem_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:271" *)
  wire [33:0] abuf_wr_elem_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:272" *)
  wire [33:0] abuf_wr_elem_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:132" *)
  output [7:0] abuf_wr_en;
  reg [7:0] abuf_wr_en;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:92" *)
  input [339:0] accu_ctrl_pd;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:93" *)
  input [191:0] accu_ctrl_ram_valid;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:94" *)
  input accu_ctrl_valid;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:273" *)
  wire [4:0] calc_addr;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1760" *)
  reg [4:0] calc_addr_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1761" *)
  reg [4:0] calc_addr_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1762" *)
  reg [4:0] calc_addr_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1763" *)
  reg [4:0] calc_addr_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:274" *)
  wire [4:0] calc_addr_out;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:275" *)
  wire calc_channel_end;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1764" *)
  reg [175:0] calc_data_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1765" *)
  reg [175:0] calc_data_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1766" *)
  reg [175:0] calc_data_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1767" *)
  reg [175:0] calc_data_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1768" *)
  reg [175:0] calc_data_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1769" *)
  reg [175:0] calc_data_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1770" *)
  reg [175:0] calc_data_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1771" *)
  reg [175:0] calc_data_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:276" *)
  wire [43:0] calc_data_16_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:277" *)
  wire [43:0] calc_data_16_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:278" *)
  wire [43:0] calc_data_16_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:279" *)
  wire [43:0] calc_data_16_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:280" *)
  wire [43:0] calc_data_16_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:281" *)
  wire [43:0] calc_data_16_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:282" *)
  wire [43:0] calc_data_16_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:283" *)
  wire [43:0] calc_data_16_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:284" *)
  wire [43:0] calc_data_16_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:285" *)
  wire [43:0] calc_data_16_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:286" *)
  wire [43:0] calc_data_16_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:287" *)
  wire [43:0] calc_data_16_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:288" *)
  wire [43:0] calc_data_16_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:289" *)
  wire [43:0] calc_data_16_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:290" *)
  wire [43:0] calc_data_16_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:291" *)
  wire [43:0] calc_data_16_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:292" *)
  wire [43:0] calc_data_16_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:293" *)
  wire [43:0] calc_data_16_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:294" *)
  wire [43:0] calc_data_16_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:295" *)
  wire [43:0] calc_data_16_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:296" *)
  wire [43:0] calc_data_16_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:297" *)
  wire [43:0] calc_data_16_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:298" *)
  wire [43:0] calc_data_16_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:299" *)
  wire [43:0] calc_data_16_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:300" *)
  wire [43:0] calc_data_16_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:301" *)
  wire [43:0] calc_data_16_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:302" *)
  wire [43:0] calc_data_16_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:303" *)
  wire [43:0] calc_data_16_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:304" *)
  wire [43:0] calc_data_16_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:305" *)
  wire [43:0] calc_data_16_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:306" *)
  wire [43:0] calc_data_16_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:307" *)
  wire [43:0] calc_data_16_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:308" *)
  wire [43:0] calc_data_16_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:309" *)
  wire [43:0] calc_data_16_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:310" *)
  wire [43:0] calc_data_16_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:311" *)
  wire [43:0] calc_data_16_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:312" *)
  wire [43:0] calc_data_16_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:313" *)
  wire [43:0] calc_data_16_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:314" *)
  wire [43:0] calc_data_16_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:315" *)
  wire [43:0] calc_data_16_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:316" *)
  wire [43:0] calc_data_16_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:317" *)
  wire [43:0] calc_data_16_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:318" *)
  wire [43:0] calc_data_16_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:319" *)
  wire [43:0] calc_data_16_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:320" *)
  wire [43:0] calc_data_16_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:321" *)
  wire [43:0] calc_data_16_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:322" *)
  wire [43:0] calc_data_16_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:323" *)
  wire [43:0] calc_data_16_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:324" *)
  wire [43:0] calc_data_16_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:325" *)
  wire [43:0] calc_data_16_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:326" *)
  wire [43:0] calc_data_16_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:327" *)
  wire [43:0] calc_data_16_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:328" *)
  wire [43:0] calc_data_16_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:329" *)
  wire [43:0] calc_data_16_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:330" *)
  wire [43:0] calc_data_16_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:331" *)
  wire [43:0] calc_data_16_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:332" *)
  wire [43:0] calc_data_16_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:333" *)
  wire [43:0] calc_data_16_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:334" *)
  wire [43:0] calc_data_16_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:335" *)
  wire [43:0] calc_data_16_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:336" *)
  wire [43:0] calc_data_16_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:337" *)
  wire [43:0] calc_data_16_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:338" *)
  wire [43:0] calc_data_16_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:339" *)
  wire [43:0] calc_data_16_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1772" *)
  reg [175:0] calc_data_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1773" *)
  reg [175:0] calc_data_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1774" *)
  reg [175:0] calc_data_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1775" *)
  reg [175:0] calc_data_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1776" *)
  reg [175:0] calc_data_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1777" *)
  reg [175:0] calc_data_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1778" *)
  reg [175:0] calc_data_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:340" *)
  wire [43:0] calc_data_8_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:341" *)
  wire [21:0] calc_data_8_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:342" *)
  wire [43:0] calc_data_8_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:343" *)
  wire [43:0] calc_data_8_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:344" *)
  wire [21:0] calc_data_8_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:345" *)
  wire [43:0] calc_data_8_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:346" *)
  wire [21:0] calc_data_8_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:347" *)
  wire [43:0] calc_data_8_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:348" *)
  wire [21:0] calc_data_8_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:349" *)
  wire [43:0] calc_data_8_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:350" *)
  wire [21:0] calc_data_8_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:351" *)
  wire [43:0] calc_data_8_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:352" *)
  wire [21:0] calc_data_8_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:353" *)
  wire [21:0] calc_data_8_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:354" *)
  wire [43:0] calc_data_8_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:355" *)
  wire [21:0] calc_data_8_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:356" *)
  wire [43:0] calc_data_8_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:357" *)
  wire [21:0] calc_data_8_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:358" *)
  wire [43:0] calc_data_8_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:359" *)
  wire [21:0] calc_data_8_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:360" *)
  wire [43:0] calc_data_8_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:361" *)
  wire [21:0] calc_data_8_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:362" *)
  wire [43:0] calc_data_8_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:363" *)
  wire [21:0] calc_data_8_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:364" *)
  wire [43:0] calc_data_8_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:365" *)
  wire [43:0] calc_data_8_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:366" *)
  wire [21:0] calc_data_8_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:367" *)
  wire [43:0] calc_data_8_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:368" *)
  wire [21:0] calc_data_8_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:369" *)
  wire [43:0] calc_data_8_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:370" *)
  wire [21:0] calc_data_8_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:371" *)
  wire [43:0] calc_data_8_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:372" *)
  wire [21:0] calc_data_8_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:373" *)
  wire [21:0] calc_data_8_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:374" *)
  wire [43:0] calc_data_8_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:375" *)
  wire [21:0] calc_data_8_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:376" *)
  wire [43:0] calc_data_8_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:377" *)
  wire [21:0] calc_data_8_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:378" *)
  wire [43:0] calc_data_8_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:379" *)
  wire [21:0] calc_data_8_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:380" *)
  wire [43:0] calc_data_8_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:381" *)
  wire [43:0] calc_data_8_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:382" *)
  wire [21:0] calc_data_8_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:383" *)
  wire [43:0] calc_data_8_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:384" *)
  wire [21:0] calc_data_8_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:385" *)
  wire [43:0] calc_data_8_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:386" *)
  wire [21:0] calc_data_8_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:387" *)
  wire [43:0] calc_data_8_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:388" *)
  wire [21:0] calc_data_8_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:389" *)
  wire [43:0] calc_data_8_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:390" *)
  wire [21:0] calc_data_8_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:391" *)
  wire [21:0] calc_data_8_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:392" *)
  wire [43:0] calc_data_8_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:393" *)
  wire [21:0] calc_data_8_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:394" *)
  wire [43:0] calc_data_8_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:395" *)
  wire [21:0] calc_data_8_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:396" *)
  wire [43:0] calc_data_8_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:397" *)
  wire [21:0] calc_data_8_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:398" *)
  wire [43:0] calc_data_8_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:399" *)
  wire [21:0] calc_data_8_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:400" *)
  wire [43:0] calc_data_8_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:401" *)
  wire [21:0] calc_data_8_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:402" *)
  wire [43:0] calc_data_8_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:403" *)
  wire [43:0] calc_data_8_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:404" *)
  wire [21:0] calc_data_8_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:405" *)
  wire [43:0] calc_data_8_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:406" *)
  wire [21:0] calc_data_8_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:407" *)
  wire [43:0] calc_data_8_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:408" *)
  wire [21:0] calc_data_8_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:409" *)
  wire [43:0] calc_data_8_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:410" *)
  wire [21:0] calc_data_8_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:411" *)
  wire [43:0] calc_data_8_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:412" *)
  wire [21:0] calc_data_8_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:413" *)
  wire [21:0] calc_data_8_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:414" *)
  wire [43:0] calc_data_8_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:415" *)
  wire [21:0] calc_data_8_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:416" *)
  wire [43:0] calc_data_8_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:417" *)
  wire [21:0] calc_data_8_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:418" *)
  wire [43:0] calc_data_8_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:419" *)
  wire [21:0] calc_data_8_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:420" *)
  wire [43:0] calc_data_8_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:421" *)
  wire [21:0] calc_data_8_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:422" *)
  wire [43:0] calc_data_8_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:423" *)
  wire [21:0] calc_data_8_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:424" *)
  wire [43:0] calc_data_8_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:425" *)
  wire [43:0] calc_data_8_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:426" *)
  wire [21:0] calc_data_8_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:427" *)
  wire [43:0] calc_data_8_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:428" *)
  wire [21:0] calc_data_8_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:429" *)
  wire [43:0] calc_data_8_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:430" *)
  wire [21:0] calc_data_8_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:431" *)
  wire [43:0] calc_data_8_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:432" *)
  wire [21:0] calc_data_8_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:433" *)
  wire [43:0] calc_data_8_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:434" *)
  wire [21:0] calc_data_8_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:435" *)
  wire [21:0] calc_data_8_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:436" *)
  wire [43:0] calc_data_8_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:437" *)
  wire [21:0] calc_data_8_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:438" *)
  wire [43:0] calc_data_8_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:439" *)
  wire [21:0] calc_data_8_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:440" *)
  wire [43:0] calc_data_8_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:441" *)
  wire [21:0] calc_data_8_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:442" *)
  wire [43:0] calc_data_8_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:443" *)
  wire [21:0] calc_data_8_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:444" *)
  wire [43:0] calc_data_8_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:445" *)
  wire [21:0] calc_data_8_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:446" *)
  wire [43:0] calc_data_8_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:447" *)
  wire [43:0] calc_data_8_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:448" *)
  wire [21:0] calc_data_8_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:449" *)
  wire [43:0] calc_data_8_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:450" *)
  wire [21:0] calc_data_8_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:451" *)
  wire [43:0] calc_data_8_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:452" *)
  wire [21:0] calc_data_8_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:453" *)
  wire [43:0] calc_data_8_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:454" *)
  wire [21:0] calc_data_8_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:455" *)
  wire [43:0] calc_data_8_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:456" *)
  wire [21:0] calc_data_8_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:457" *)
  wire [21:0] calc_data_8_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:458" *)
  wire [43:0] calc_data_8_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:459" *)
  wire [21:0] calc_data_8_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:460" *)
  wire [43:0] calc_data_8_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:461" *)
  wire [21:0] calc_data_8_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:462" *)
  wire [43:0] calc_data_8_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:463" *)
  wire [21:0] calc_data_8_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:464" *)
  wire [43:0] calc_data_8_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:465" *)
  wire [21:0] calc_data_8_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:466" *)
  wire [43:0] calc_data_8_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:467" *)
  wire [21:0] calc_data_8_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1779" *)
  reg [175:0] calc_data_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:468" *)
  wire [2815:0] calc_data_all;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:469" *)
  wire [31:0] calc_dlv_elem_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:470" *)
  wire [31:0] calc_dlv_elem_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:471" *)
  wire [31:0] calc_dlv_elem_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:472" *)
  wire [31:0] calc_dlv_elem_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:473" *)
  wire [31:0] calc_dlv_elem_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:474" *)
  wire [31:0] calc_dlv_elem_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:475" *)
  wire [31:0] calc_dlv_elem_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:476" *)
  wire [31:0] calc_dlv_elem_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:477" *)
  wire [31:0] calc_dlv_elem_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:478" *)
  wire [31:0] calc_dlv_elem_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:479" *)
  wire [31:0] calc_dlv_elem_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:480" *)
  wire [31:0] calc_dlv_elem_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:481" *)
  wire [31:0] calc_dlv_elem_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:482" *)
  wire [31:0] calc_dlv_elem_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:483" *)
  wire [31:0] calc_dlv_elem_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:484" *)
  wire [31:0] calc_dlv_elem_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:485" *)
  wire [31:0] calc_dlv_elem_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:486" *)
  wire [31:0] calc_dlv_elem_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:487" *)
  wire [31:0] calc_dlv_elem_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:488" *)
  wire [31:0] calc_dlv_elem_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:489" *)
  wire [31:0] calc_dlv_elem_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:490" *)
  wire [31:0] calc_dlv_elem_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:491" *)
  wire [31:0] calc_dlv_elem_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:492" *)
  wire [31:0] calc_dlv_elem_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:493" *)
  wire [31:0] calc_dlv_elem_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:494" *)
  wire [31:0] calc_dlv_elem_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:495" *)
  wire [31:0] calc_dlv_elem_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:496" *)
  wire [31:0] calc_dlv_elem_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:497" *)
  wire [31:0] calc_dlv_elem_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:498" *)
  wire [31:0] calc_dlv_elem_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:499" *)
  wire [31:0] calc_dlv_elem_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:500" *)
  wire [31:0] calc_dlv_elem_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:501" *)
  wire [31:0] calc_dlv_elem_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:502" *)
  wire [31:0] calc_dlv_elem_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:503" *)
  wire [31:0] calc_dlv_elem_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:504" *)
  wire [31:0] calc_dlv_elem_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:505" *)
  wire [31:0] calc_dlv_elem_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:506" *)
  wire [31:0] calc_dlv_elem_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:507" *)
  wire [31:0] calc_dlv_elem_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:508" *)
  wire [31:0] calc_dlv_elem_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:509" *)
  wire [31:0] calc_dlv_elem_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:510" *)
  wire [31:0] calc_dlv_elem_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:511" *)
  wire [31:0] calc_dlv_elem_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:512" *)
  wire [31:0] calc_dlv_elem_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:513" *)
  wire [31:0] calc_dlv_elem_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:514" *)
  wire [31:0] calc_dlv_elem_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:515" *)
  wire [31:0] calc_dlv_elem_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:516" *)
  wire [31:0] calc_dlv_elem_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:517" *)
  wire [31:0] calc_dlv_elem_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:518" *)
  wire [31:0] calc_dlv_elem_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:519" *)
  wire [31:0] calc_dlv_elem_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:520" *)
  wire [31:0] calc_dlv_elem_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:521" *)
  wire [31:0] calc_dlv_elem_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:522" *)
  wire [31:0] calc_dlv_elem_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:523" *)
  wire [31:0] calc_dlv_elem_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:524" *)
  wire [31:0] calc_dlv_elem_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:525" *)
  wire [31:0] calc_dlv_elem_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:526" *)
  wire [31:0] calc_dlv_elem_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:527" *)
  wire [31:0] calc_dlv_elem_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:528" *)
  wire [31:0] calc_dlv_elem_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:529" *)
  wire [31:0] calc_dlv_elem_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:530" *)
  wire [31:0] calc_dlv_elem_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:531" *)
  wire [31:0] calc_dlv_elem_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:532" *)
  wire [31:0] calc_dlv_elem_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:533" *)
  wire [31:0] calc_dlv_elem_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:534" *)
  wire [31:0] calc_dlv_elem_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:535" *)
  wire [31:0] calc_dlv_elem_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:536" *)
  wire [31:0] calc_dlv_elem_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:537" *)
  wire [31:0] calc_dlv_elem_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:538" *)
  wire [31:0] calc_dlv_elem_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:539" *)
  wire [31:0] calc_dlv_elem_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:540" *)
  wire [31:0] calc_dlv_elem_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:541" *)
  wire [31:0] calc_dlv_elem_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:542" *)
  wire [31:0] calc_dlv_elem_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:543" *)
  wire [31:0] calc_dlv_elem_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:544" *)
  wire [31:0] calc_dlv_elem_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:545" *)
  wire [31:0] calc_dlv_elem_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:546" *)
  wire [31:0] calc_dlv_elem_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:547" *)
  wire [31:0] calc_dlv_elem_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:548" *)
  wire [31:0] calc_dlv_elem_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:549" *)
  wire [31:0] calc_dlv_elem_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:550" *)
  wire [31:0] calc_dlv_elem_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:551" *)
  wire [31:0] calc_dlv_elem_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:552" *)
  wire [31:0] calc_dlv_elem_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:553" *)
  wire [31:0] calc_dlv_elem_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:554" *)
  wire [31:0] calc_dlv_elem_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:555" *)
  wire [31:0] calc_dlv_elem_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:556" *)
  wire [31:0] calc_dlv_elem_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:557" *)
  wire [31:0] calc_dlv_elem_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:558" *)
  wire [31:0] calc_dlv_elem_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:559" *)
  wire [31:0] calc_dlv_elem_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:560" *)
  wire [31:0] calc_dlv_elem_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:561" *)
  wire [31:0] calc_dlv_elem_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:562" *)
  wire [31:0] calc_dlv_elem_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:563" *)
  wire [31:0] calc_dlv_elem_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:564" *)
  wire [31:0] calc_dlv_elem_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:565" *)
  wire [31:0] calc_dlv_elem_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:566" *)
  wire [31:0] calc_dlv_elem_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:567" *)
  wire [31:0] calc_dlv_elem_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:568" *)
  wire [31:0] calc_dlv_elem_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:569" *)
  wire [31:0] calc_dlv_elem_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:570" *)
  wire [31:0] calc_dlv_elem_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:571" *)
  wire [31:0] calc_dlv_elem_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:572" *)
  wire [31:0] calc_dlv_elem_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:573" *)
  wire [31:0] calc_dlv_elem_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:574" *)
  wire [31:0] calc_dlv_elem_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:575" *)
  wire [31:0] calc_dlv_elem_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:576" *)
  wire [31:0] calc_dlv_elem_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:577" *)
  wire [31:0] calc_dlv_elem_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:578" *)
  wire [31:0] calc_dlv_elem_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:579" *)
  wire [31:0] calc_dlv_elem_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:580" *)
  wire [31:0] calc_dlv_elem_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:581" *)
  wire [31:0] calc_dlv_elem_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:582" *)
  wire [31:0] calc_dlv_elem_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:583" *)
  wire [31:0] calc_dlv_elem_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:584" *)
  wire [31:0] calc_dlv_elem_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:585" *)
  wire [31:0] calc_dlv_elem_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:586" *)
  wire [31:0] calc_dlv_elem_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:587" *)
  wire [31:0] calc_dlv_elem_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:588" *)
  wire [31:0] calc_dlv_elem_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:589" *)
  wire [31:0] calc_dlv_elem_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:590" *)
  wire [31:0] calc_dlv_elem_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:591" *)
  wire [31:0] calc_dlv_elem_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:592" *)
  wire [31:0] calc_dlv_elem_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:593" *)
  wire [31:0] calc_dlv_elem_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:594" *)
  wire [31:0] calc_dlv_elem_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:595" *)
  wire [31:0] calc_dlv_elem_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:596" *)
  wire [31:0] calc_dlv_elem_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:597" *)
  wire [191:0] calc_dlv_elem_en;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:598" *)
  wire [191:0] calc_dlv_elem_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1780" *)
  wire [7:0] calc_dlv_en;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1781" *)
  reg [7:0] calc_dlv_en_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1782" *)
  reg [7:0] calc_dlv_en_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1783" *)
  reg [7:0] calc_dlv_en_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1784" *)
  reg [7:0] calc_dlv_en_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1785" *)
  reg [7:0] calc_dlv_en_d5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:599" *)
  wire [63:0] calc_dlv_en_fp;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1786" *)
  reg [63:0] calc_dlv_en_fp_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:600" *)
  wire [127:0] calc_dlv_en_int;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1787" *)
  reg [127:0] calc_dlv_en_int_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:601" *)
  wire [7:0] calc_dlv_en_out;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1788" *)
  wire calc_dlv_valid;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1789" *)
  reg calc_dlv_valid_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1790" *)
  reg calc_dlv_valid_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1791" *)
  reg calc_dlv_valid_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1792" *)
  reg calc_dlv_valid_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1793" *)
  reg calc_dlv_valid_d5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:602" *)
  wire calc_dlv_valid_out;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:603" *)
  wire [43:0] calc_elem_0_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:604" *)
  wire [21:0] calc_elem_100_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:605" *)
  wire [21:0] calc_elem_101_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:606" *)
  wire [21:0] calc_elem_102_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:607" *)
  wire [21:0] calc_elem_103_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:608" *)
  wire [21:0] calc_elem_104_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:609" *)
  wire [21:0] calc_elem_105_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:610" *)
  wire [21:0] calc_elem_106_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:611" *)
  wire [21:0] calc_elem_107_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:612" *)
  wire [21:0] calc_elem_108_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:613" *)
  wire [21:0] calc_elem_109_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:614" *)
  wire [43:0] calc_elem_10_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:615" *)
  wire [21:0] calc_elem_110_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:616" *)
  wire [21:0] calc_elem_111_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:617" *)
  wire [21:0] calc_elem_112_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:618" *)
  wire [21:0] calc_elem_113_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:619" *)
  wire [21:0] calc_elem_114_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:620" *)
  wire [21:0] calc_elem_115_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:621" *)
  wire [21:0] calc_elem_116_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:622" *)
  wire [21:0] calc_elem_117_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:623" *)
  wire [21:0] calc_elem_118_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:624" *)
  wire [21:0] calc_elem_119_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:625" *)
  wire [43:0] calc_elem_11_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:626" *)
  wire [21:0] calc_elem_120_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:627" *)
  wire [21:0] calc_elem_121_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:628" *)
  wire [21:0] calc_elem_122_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:629" *)
  wire [21:0] calc_elem_123_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:630" *)
  wire [21:0] calc_elem_124_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:631" *)
  wire [21:0] calc_elem_125_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:632" *)
  wire [21:0] calc_elem_126_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:633" *)
  wire [21:0] calc_elem_127_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:634" *)
  wire [43:0] calc_elem_12_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:635" *)
  wire [43:0] calc_elem_13_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:636" *)
  wire [43:0] calc_elem_14_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:637" *)
  wire [43:0] calc_elem_15_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:638" *)
  wire [43:0] calc_elem_16_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:639" *)
  wire [43:0] calc_elem_17_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:640" *)
  wire [43:0] calc_elem_18_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:641" *)
  wire [43:0] calc_elem_19_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:642" *)
  wire [43:0] calc_elem_1_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:643" *)
  wire [43:0] calc_elem_20_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:644" *)
  wire [43:0] calc_elem_21_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:645" *)
  wire [43:0] calc_elem_22_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:646" *)
  wire [43:0] calc_elem_23_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:647" *)
  wire [43:0] calc_elem_24_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:648" *)
  wire [43:0] calc_elem_25_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:649" *)
  wire [43:0] calc_elem_26_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:650" *)
  wire [43:0] calc_elem_27_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:651" *)
  wire [43:0] calc_elem_28_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:652" *)
  wire [43:0] calc_elem_29_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:653" *)
  wire [43:0] calc_elem_2_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:654" *)
  wire [43:0] calc_elem_30_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:655" *)
  wire [43:0] calc_elem_31_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:656" *)
  wire [43:0] calc_elem_32_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:657" *)
  wire [43:0] calc_elem_33_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:658" *)
  wire [43:0] calc_elem_34_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:659" *)
  wire [43:0] calc_elem_35_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:660" *)
  wire [43:0] calc_elem_36_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:661" *)
  wire [43:0] calc_elem_37_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:662" *)
  wire [43:0] calc_elem_38_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:663" *)
  wire [43:0] calc_elem_39_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:664" *)
  wire [43:0] calc_elem_3_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:665" *)
  wire [43:0] calc_elem_40_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:666" *)
  wire [43:0] calc_elem_41_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:667" *)
  wire [43:0] calc_elem_42_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:668" *)
  wire [43:0] calc_elem_43_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:669" *)
  wire [43:0] calc_elem_44_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:670" *)
  wire [43:0] calc_elem_45_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:671" *)
  wire [43:0] calc_elem_46_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:672" *)
  wire [43:0] calc_elem_47_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:673" *)
  wire [43:0] calc_elem_48_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:674" *)
  wire [43:0] calc_elem_49_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:675" *)
  wire [43:0] calc_elem_4_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:676" *)
  wire [43:0] calc_elem_50_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:677" *)
  wire [43:0] calc_elem_51_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:678" *)
  wire [43:0] calc_elem_52_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:679" *)
  wire [43:0] calc_elem_53_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:680" *)
  wire [43:0] calc_elem_54_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:681" *)
  wire [43:0] calc_elem_55_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:682" *)
  wire [43:0] calc_elem_56_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:683" *)
  wire [43:0] calc_elem_57_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:684" *)
  wire [43:0] calc_elem_58_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:685" *)
  wire [43:0] calc_elem_59_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:686" *)
  wire [43:0] calc_elem_5_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:687" *)
  wire [43:0] calc_elem_60_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:688" *)
  wire [43:0] calc_elem_61_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:689" *)
  wire [43:0] calc_elem_62_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:690" *)
  wire [43:0] calc_elem_63_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:691" *)
  wire [21:0] calc_elem_64_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:692" *)
  wire [21:0] calc_elem_65_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:693" *)
  wire [21:0] calc_elem_66_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:694" *)
  wire [21:0] calc_elem_67_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:695" *)
  wire [21:0] calc_elem_68_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:696" *)
  wire [21:0] calc_elem_69_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:697" *)
  wire [43:0] calc_elem_6_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:698" *)
  wire [21:0] calc_elem_70_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:699" *)
  wire [21:0] calc_elem_71_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:700" *)
  wire [21:0] calc_elem_72_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:701" *)
  wire [21:0] calc_elem_73_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:702" *)
  wire [21:0] calc_elem_74_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:703" *)
  wire [21:0] calc_elem_75_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:704" *)
  wire [21:0] calc_elem_76_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:705" *)
  wire [21:0] calc_elem_77_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:706" *)
  wire [21:0] calc_elem_78_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:707" *)
  wire [21:0] calc_elem_79_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:708" *)
  wire [43:0] calc_elem_7_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:709" *)
  wire [21:0] calc_elem_80_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:710" *)
  wire [21:0] calc_elem_81_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:711" *)
  wire [21:0] calc_elem_82_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:712" *)
  wire [21:0] calc_elem_83_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:713" *)
  wire [21:0] calc_elem_84_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:714" *)
  wire [21:0] calc_elem_85_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:715" *)
  wire [21:0] calc_elem_86_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:716" *)
  wire [21:0] calc_elem_87_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:717" *)
  wire [21:0] calc_elem_88_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:718" *)
  wire [21:0] calc_elem_89_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:719" *)
  wire [43:0] calc_elem_8_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:720" *)
  wire [21:0] calc_elem_90_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:721" *)
  wire [21:0] calc_elem_91_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:722" *)
  wire [21:0] calc_elem_92_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:723" *)
  wire [21:0] calc_elem_93_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:724" *)
  wire [21:0] calc_elem_94_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:725" *)
  wire [21:0] calc_elem_95_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:726" *)
  wire [21:0] calc_elem_96_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:727" *)
  wire [21:0] calc_elem_97_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:728" *)
  wire [21:0] calc_elem_98_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:729" *)
  wire [21:0] calc_elem_99_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:730" *)
  wire [43:0] calc_elem_9_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:731" *)
  wire [191:0] calc_elem_en;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:732" *)
  wire [191:0] calc_elem_op1_vld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:733" *)
  wire [31:0] calc_fout_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:734" *)
  wire [31:0] calc_fout_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:735" *)
  wire [31:0] calc_fout_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:736" *)
  wire [31:0] calc_fout_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:737" *)
  wire [31:0] calc_fout_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:738" *)
  wire [31:0] calc_fout_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:739" *)
  wire [31:0] calc_fout_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:740" *)
  wire [31:0] calc_fout_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:741" *)
  wire [31:0] calc_fout_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:742" *)
  wire [31:0] calc_fout_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:743" *)
  wire [31:0] calc_fout_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:744" *)
  wire [31:0] calc_fout_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:745" *)
  wire [31:0] calc_fout_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:746" *)
  wire [31:0] calc_fout_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:747" *)
  wire [31:0] calc_fout_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:748" *)
  wire [31:0] calc_fout_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:749" *)
  wire [31:0] calc_fout_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:750" *)
  wire [31:0] calc_fout_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:751" *)
  wire [31:0] calc_fout_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:752" *)
  wire [31:0] calc_fout_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:753" *)
  wire [31:0] calc_fout_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:754" *)
  wire [31:0] calc_fout_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:755" *)
  wire [31:0] calc_fout_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:756" *)
  wire [31:0] calc_fout_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:757" *)
  wire [31:0] calc_fout_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:758" *)
  wire [31:0] calc_fout_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:759" *)
  wire [31:0] calc_fout_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:760" *)
  wire [31:0] calc_fout_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:761" *)
  wire [31:0] calc_fout_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:762" *)
  wire [31:0] calc_fout_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:763" *)
  wire [31:0] calc_fout_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:764" *)
  wire [31:0] calc_fout_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:765" *)
  wire [31:0] calc_fout_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:766" *)
  wire [31:0] calc_fout_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:767" *)
  wire [31:0] calc_fout_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:768" *)
  wire [31:0] calc_fout_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:769" *)
  wire [31:0] calc_fout_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:770" *)
  wire [31:0] calc_fout_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:771" *)
  wire [31:0] calc_fout_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:772" *)
  wire [31:0] calc_fout_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:773" *)
  wire [31:0] calc_fout_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:774" *)
  wire [31:0] calc_fout_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:775" *)
  wire [31:0] calc_fout_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:776" *)
  wire [31:0] calc_fout_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:777" *)
  wire [31:0] calc_fout_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:778" *)
  wire [31:0] calc_fout_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:779" *)
  wire [31:0] calc_fout_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:780" *)
  wire [31:0] calc_fout_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:781" *)
  wire [31:0] calc_fout_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:782" *)
  wire [31:0] calc_fout_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:783" *)
  wire [31:0] calc_fout_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:784" *)
  wire [31:0] calc_fout_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:785" *)
  wire [31:0] calc_fout_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:786" *)
  wire [31:0] calc_fout_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:787" *)
  wire [31:0] calc_fout_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:788" *)
  wire [31:0] calc_fout_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:789" *)
  wire [31:0] calc_fout_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:790" *)
  wire [31:0] calc_fout_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:791" *)
  wire [31:0] calc_fout_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:792" *)
  wire [31:0] calc_fout_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:793" *)
  wire [31:0] calc_fout_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:794" *)
  wire [31:0] calc_fout_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:795" *)
  wire [31:0] calc_fout_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:796" *)
  wire [31:0] calc_fout_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:797" *)
  wire [31:0] calc_fout_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:798" *)
  wire [31:0] calc_fout_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:799" *)
  wire [31:0] calc_fout_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:800" *)
  wire [31:0] calc_fout_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:801" *)
  wire [31:0] calc_fout_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:802" *)
  wire [31:0] calc_fout_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:803" *)
  wire [31:0] calc_fout_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:804" *)
  wire [31:0] calc_fout_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:805" *)
  wire [31:0] calc_fout_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:806" *)
  wire [31:0] calc_fout_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:807" *)
  wire [31:0] calc_fout_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:808" *)
  wire [31:0] calc_fout_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:809" *)
  wire [31:0] calc_fout_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:810" *)
  wire [31:0] calc_fout_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:811" *)
  wire [31:0] calc_fout_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:812" *)
  wire [31:0] calc_fout_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:813" *)
  wire [31:0] calc_fout_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:814" *)
  wire [31:0] calc_fout_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:815" *)
  wire [31:0] calc_fout_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:816" *)
  wire [31:0] calc_fout_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:817" *)
  wire [31:0] calc_fout_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:818" *)
  wire [31:0] calc_fout_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:819" *)
  wire [31:0] calc_fout_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:820" *)
  wire [31:0] calc_fout_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:821" *)
  wire [31:0] calc_fout_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:822" *)
  wire [31:0] calc_fout_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:823" *)
  wire [31:0] calc_fout_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:824" *)
  wire [31:0] calc_fout_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:825" *)
  wire [31:0] calc_fout_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:826" *)
  wire [31:0] calc_fout_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:827" *)
  wire [31:0] calc_fout_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:828" *)
  wire [31:0] calc_fout_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:829" *)
  wire [31:0] calc_fout_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:830" *)
  wire [31:0] calc_fout_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:831" *)
  wire [31:0] calc_fout_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:832" *)
  wire [31:0] calc_fout_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:833" *)
  wire [31:0] calc_fout_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:834" *)
  wire [31:0] calc_fout_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:835" *)
  wire [31:0] calc_fout_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:836" *)
  wire [31:0] calc_fout_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:837" *)
  wire [31:0] calc_fout_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:838" *)
  wire [31:0] calc_fout_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:839" *)
  wire [31:0] calc_fout_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:840" *)
  wire [31:0] calc_fout_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:841" *)
  wire [31:0] calc_fout_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:842" *)
  wire [31:0] calc_fout_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:843" *)
  wire [31:0] calc_fout_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:844" *)
  wire [31:0] calc_fout_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:845" *)
  wire [31:0] calc_fout_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:846" *)
  wire [31:0] calc_fout_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:847" *)
  wire [31:0] calc_fout_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:848" *)
  wire [31:0] calc_fout_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:849" *)
  wire [31:0] calc_fout_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:850" *)
  wire [31:0] calc_fout_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:851" *)
  wire [31:0] calc_fout_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:852" *)
  wire [31:0] calc_fout_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:853" *)
  wire [31:0] calc_fout_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:854" *)
  wire [31:0] calc_fout_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:855" *)
  wire [31:0] calc_fout_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:856" *)
  wire [31:0] calc_fout_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:857" *)
  wire [31:0] calc_fout_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:858" *)
  wire [31:0] calc_fout_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:859" *)
  wire [31:0] calc_fout_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:860" *)
  wire [31:0] calc_fout_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:861" *)
  wire [31:0] calc_fout_fp_0_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:862" *)
  wire [31:0] calc_fout_fp_10_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:863" *)
  wire [31:0] calc_fout_fp_11_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:864" *)
  wire [31:0] calc_fout_fp_12_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:865" *)
  wire [31:0] calc_fout_fp_13_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:866" *)
  wire [31:0] calc_fout_fp_14_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:867" *)
  wire [31:0] calc_fout_fp_15_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:868" *)
  wire [31:0] calc_fout_fp_16_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:869" *)
  wire [31:0] calc_fout_fp_17_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:870" *)
  wire [31:0] calc_fout_fp_18_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:871" *)
  wire [31:0] calc_fout_fp_19_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:872" *)
  wire [31:0] calc_fout_fp_1_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:873" *)
  wire [31:0] calc_fout_fp_20_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:874" *)
  wire [31:0] calc_fout_fp_21_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:875" *)
  wire [31:0] calc_fout_fp_22_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:876" *)
  wire [31:0] calc_fout_fp_23_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:877" *)
  wire [31:0] calc_fout_fp_24_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:878" *)
  wire [31:0] calc_fout_fp_25_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:879" *)
  wire [31:0] calc_fout_fp_26_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:880" *)
  wire [31:0] calc_fout_fp_27_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:881" *)
  wire [31:0] calc_fout_fp_28_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:882" *)
  wire [31:0] calc_fout_fp_29_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:883" *)
  wire [31:0] calc_fout_fp_2_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:884" *)
  wire [31:0] calc_fout_fp_30_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:885" *)
  wire [31:0] calc_fout_fp_31_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:886" *)
  wire [31:0] calc_fout_fp_32_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:887" *)
  wire [31:0] calc_fout_fp_33_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:888" *)
  wire [31:0] calc_fout_fp_34_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:889" *)
  wire [31:0] calc_fout_fp_35_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:890" *)
  wire [31:0] calc_fout_fp_36_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:891" *)
  wire [31:0] calc_fout_fp_37_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:892" *)
  wire [31:0] calc_fout_fp_38_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:893" *)
  wire [31:0] calc_fout_fp_39_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:894" *)
  wire [31:0] calc_fout_fp_3_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:895" *)
  wire [31:0] calc_fout_fp_40_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:896" *)
  wire [31:0] calc_fout_fp_41_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:897" *)
  wire [31:0] calc_fout_fp_42_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:898" *)
  wire [31:0] calc_fout_fp_43_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:899" *)
  wire [31:0] calc_fout_fp_44_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:900" *)
  wire [31:0] calc_fout_fp_45_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:901" *)
  wire [31:0] calc_fout_fp_46_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:902" *)
  wire [31:0] calc_fout_fp_47_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:903" *)
  wire [31:0] calc_fout_fp_48_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:904" *)
  wire [31:0] calc_fout_fp_49_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:905" *)
  wire [31:0] calc_fout_fp_4_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:906" *)
  wire [31:0] calc_fout_fp_50_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:907" *)
  wire [31:0] calc_fout_fp_51_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:908" *)
  wire [31:0] calc_fout_fp_52_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:909" *)
  wire [31:0] calc_fout_fp_53_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:910" *)
  wire [31:0] calc_fout_fp_54_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:911" *)
  wire [31:0] calc_fout_fp_55_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:912" *)
  wire [31:0] calc_fout_fp_56_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:913" *)
  wire [31:0] calc_fout_fp_57_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:914" *)
  wire [31:0] calc_fout_fp_58_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:915" *)
  wire [31:0] calc_fout_fp_59_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:916" *)
  wire [31:0] calc_fout_fp_5_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:917" *)
  wire [31:0] calc_fout_fp_60_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:918" *)
  wire [31:0] calc_fout_fp_61_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:919" *)
  wire [31:0] calc_fout_fp_62_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:920" *)
  wire [31:0] calc_fout_fp_63_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:921" *)
  wire [31:0] calc_fout_fp_6_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:922" *)
  wire [31:0] calc_fout_fp_7_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:923" *)
  wire [31:0] calc_fout_fp_8_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:924" *)
  wire [31:0] calc_fout_fp_9_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:925" *)
  wire [63:0] calc_fout_fp_vld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:926" *)
  wire [31:0] calc_fout_int_0_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:927" *)
  wire [31:0] calc_fout_int_100_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:928" *)
  wire [31:0] calc_fout_int_101_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:929" *)
  wire [31:0] calc_fout_int_102_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:930" *)
  wire [31:0] calc_fout_int_103_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:931" *)
  wire [31:0] calc_fout_int_104_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:932" *)
  wire [31:0] calc_fout_int_105_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:933" *)
  wire [31:0] calc_fout_int_106_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:934" *)
  wire [31:0] calc_fout_int_107_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:935" *)
  wire [31:0] calc_fout_int_108_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:936" *)
  wire [31:0] calc_fout_int_109_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:937" *)
  wire [31:0] calc_fout_int_10_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:938" *)
  wire [31:0] calc_fout_int_110_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:939" *)
  wire [31:0] calc_fout_int_111_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:940" *)
  wire [31:0] calc_fout_int_112_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:941" *)
  wire [31:0] calc_fout_int_113_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:942" *)
  wire [31:0] calc_fout_int_114_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:943" *)
  wire [31:0] calc_fout_int_115_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:944" *)
  wire [31:0] calc_fout_int_116_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:945" *)
  wire [31:0] calc_fout_int_117_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:946" *)
  wire [31:0] calc_fout_int_118_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:947" *)
  wire [31:0] calc_fout_int_119_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:948" *)
  wire [31:0] calc_fout_int_11_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:949" *)
  wire [31:0] calc_fout_int_120_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:950" *)
  wire [31:0] calc_fout_int_121_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:951" *)
  wire [31:0] calc_fout_int_122_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:952" *)
  wire [31:0] calc_fout_int_123_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:953" *)
  wire [31:0] calc_fout_int_124_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:954" *)
  wire [31:0] calc_fout_int_125_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:955" *)
  wire [31:0] calc_fout_int_126_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:956" *)
  wire [31:0] calc_fout_int_127_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:957" *)
  wire [31:0] calc_fout_int_12_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:958" *)
  wire [31:0] calc_fout_int_13_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:959" *)
  wire [31:0] calc_fout_int_14_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:960" *)
  wire [31:0] calc_fout_int_15_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:961" *)
  wire [31:0] calc_fout_int_16_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:962" *)
  wire [31:0] calc_fout_int_17_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:963" *)
  wire [31:0] calc_fout_int_18_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:964" *)
  wire [31:0] calc_fout_int_19_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:965" *)
  wire [31:0] calc_fout_int_1_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:966" *)
  wire [31:0] calc_fout_int_20_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:967" *)
  wire [31:0] calc_fout_int_21_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:968" *)
  wire [31:0] calc_fout_int_22_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:969" *)
  wire [31:0] calc_fout_int_23_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:970" *)
  wire [31:0] calc_fout_int_24_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:971" *)
  wire [31:0] calc_fout_int_25_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:972" *)
  wire [31:0] calc_fout_int_26_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:973" *)
  wire [31:0] calc_fout_int_27_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:974" *)
  wire [31:0] calc_fout_int_28_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:975" *)
  wire [31:0] calc_fout_int_29_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:976" *)
  wire [31:0] calc_fout_int_2_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:977" *)
  wire [31:0] calc_fout_int_30_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:978" *)
  wire [31:0] calc_fout_int_31_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:979" *)
  wire [31:0] calc_fout_int_32_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:980" *)
  wire [31:0] calc_fout_int_33_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:981" *)
  wire [31:0] calc_fout_int_34_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:982" *)
  wire [31:0] calc_fout_int_35_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:983" *)
  wire [31:0] calc_fout_int_36_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:984" *)
  wire [31:0] calc_fout_int_37_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:985" *)
  wire [31:0] calc_fout_int_38_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:986" *)
  wire [31:0] calc_fout_int_39_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:987" *)
  wire [31:0] calc_fout_int_3_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:988" *)
  wire [31:0] calc_fout_int_40_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:989" *)
  wire [31:0] calc_fout_int_41_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:990" *)
  wire [31:0] calc_fout_int_42_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:991" *)
  wire [31:0] calc_fout_int_43_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:992" *)
  wire [31:0] calc_fout_int_44_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:993" *)
  wire [31:0] calc_fout_int_45_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:994" *)
  wire [31:0] calc_fout_int_46_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:995" *)
  wire [31:0] calc_fout_int_47_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:996" *)
  wire [31:0] calc_fout_int_48_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:997" *)
  wire [31:0] calc_fout_int_49_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:998" *)
  wire [31:0] calc_fout_int_4_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:999" *)
  wire [31:0] calc_fout_int_50_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1000" *)
  wire [31:0] calc_fout_int_51_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1001" *)
  wire [31:0] calc_fout_int_52_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1002" *)
  wire [31:0] calc_fout_int_53_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1003" *)
  wire [31:0] calc_fout_int_54_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1004" *)
  wire [31:0] calc_fout_int_55_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1005" *)
  wire [31:0] calc_fout_int_56_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1006" *)
  wire [31:0] calc_fout_int_57_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1007" *)
  wire [31:0] calc_fout_int_58_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1008" *)
  wire [31:0] calc_fout_int_59_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1009" *)
  wire [31:0] calc_fout_int_5_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1010" *)
  wire [31:0] calc_fout_int_60_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1011" *)
  wire [31:0] calc_fout_int_61_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1012" *)
  wire [31:0] calc_fout_int_62_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1013" *)
  wire [31:0] calc_fout_int_63_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1014" *)
  wire [31:0] calc_fout_int_64_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1015" *)
  wire [31:0] calc_fout_int_65_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1016" *)
  wire [31:0] calc_fout_int_66_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1017" *)
  wire [31:0] calc_fout_int_67_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1018" *)
  wire [31:0] calc_fout_int_68_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1019" *)
  wire [31:0] calc_fout_int_69_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1020" *)
  wire [31:0] calc_fout_int_6_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1021" *)
  wire [31:0] calc_fout_int_70_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1022" *)
  wire [31:0] calc_fout_int_71_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1023" *)
  wire [31:0] calc_fout_int_72_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1024" *)
  wire [31:0] calc_fout_int_73_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1025" *)
  wire [31:0] calc_fout_int_74_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1026" *)
  wire [31:0] calc_fout_int_75_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1027" *)
  wire [31:0] calc_fout_int_76_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1028" *)
  wire [31:0] calc_fout_int_77_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1029" *)
  wire [31:0] calc_fout_int_78_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1030" *)
  wire [31:0] calc_fout_int_79_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1031" *)
  wire [31:0] calc_fout_int_7_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1032" *)
  wire [31:0] calc_fout_int_80_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1033" *)
  wire [31:0] calc_fout_int_81_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1034" *)
  wire [31:0] calc_fout_int_82_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1035" *)
  wire [31:0] calc_fout_int_83_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1036" *)
  wire [31:0] calc_fout_int_84_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1037" *)
  wire [31:0] calc_fout_int_85_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1038" *)
  wire [31:0] calc_fout_int_86_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1039" *)
  wire [31:0] calc_fout_int_87_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1040" *)
  wire [31:0] calc_fout_int_88_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1041" *)
  wire [31:0] calc_fout_int_89_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1042" *)
  wire [31:0] calc_fout_int_8_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1043" *)
  wire [31:0] calc_fout_int_90_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1044" *)
  wire [31:0] calc_fout_int_91_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1045" *)
  wire [31:0] calc_fout_int_92_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1046" *)
  wire [31:0] calc_fout_int_93_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1047" *)
  wire [31:0] calc_fout_int_94_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1048" *)
  wire [31:0] calc_fout_int_95_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1049" *)
  wire [31:0] calc_fout_int_96_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1050" *)
  wire [31:0] calc_fout_int_97_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1051" *)
  wire [31:0] calc_fout_int_98_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1052" *)
  wire [31:0] calc_fout_int_99_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1053" *)
  wire [31:0] calc_fout_int_9_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1054" *)
  wire [127:0] calc_fout_int_sat;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1055" *)
  wire [127:0] calc_fout_int_vld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1794" *)
  reg [191:0] calc_in_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1056" *)
  wire calc_layer_end;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1795" *)
  reg calc_layer_end_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1796" *)
  reg calc_layer_end_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1797" *)
  reg calc_layer_end_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1798" *)
  reg calc_layer_end_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1799" *)
  reg calc_layer_end_d5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1057" *)
  wire calc_layer_end_out;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1058" *)
  (* unused_bits = "3" *)
  wire [3:0] calc_mode;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1800" *)
  reg [43:0] calc_op0_fp_0_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1801" *)
  reg [43:0] calc_op0_fp_10_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1802" *)
  reg [43:0] calc_op0_fp_11_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1803" *)
  reg [43:0] calc_op0_fp_12_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1804" *)
  reg [43:0] calc_op0_fp_13_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1805" *)
  reg [43:0] calc_op0_fp_14_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1806" *)
  reg [43:0] calc_op0_fp_15_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1807" *)
  reg [43:0] calc_op0_fp_16_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1808" *)
  reg [43:0] calc_op0_fp_17_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1809" *)
  reg [43:0] calc_op0_fp_18_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1810" *)
  reg [43:0] calc_op0_fp_19_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1811" *)
  reg [43:0] calc_op0_fp_1_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1812" *)
  reg [43:0] calc_op0_fp_20_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1813" *)
  reg [43:0] calc_op0_fp_21_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1814" *)
  reg [43:0] calc_op0_fp_22_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1815" *)
  reg [43:0] calc_op0_fp_23_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1816" *)
  reg [43:0] calc_op0_fp_24_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1817" *)
  reg [43:0] calc_op0_fp_25_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1818" *)
  reg [43:0] calc_op0_fp_26_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1819" *)
  reg [43:0] calc_op0_fp_27_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1820" *)
  reg [43:0] calc_op0_fp_28_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1821" *)
  reg [43:0] calc_op0_fp_29_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1822" *)
  reg [43:0] calc_op0_fp_2_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1823" *)
  reg [43:0] calc_op0_fp_30_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1824" *)
  reg [43:0] calc_op0_fp_31_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1825" *)
  reg [43:0] calc_op0_fp_32_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1826" *)
  reg [43:0] calc_op0_fp_33_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1827" *)
  reg [43:0] calc_op0_fp_34_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1828" *)
  reg [43:0] calc_op0_fp_35_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1829" *)
  reg [43:0] calc_op0_fp_36_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1830" *)
  reg [43:0] calc_op0_fp_37_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1831" *)
  reg [43:0] calc_op0_fp_38_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1832" *)
  reg [43:0] calc_op0_fp_39_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1833" *)
  reg [43:0] calc_op0_fp_3_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1834" *)
  reg [43:0] calc_op0_fp_40_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1835" *)
  reg [43:0] calc_op0_fp_41_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1836" *)
  reg [43:0] calc_op0_fp_42_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1837" *)
  reg [43:0] calc_op0_fp_43_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1838" *)
  reg [43:0] calc_op0_fp_44_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1839" *)
  reg [43:0] calc_op0_fp_45_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1840" *)
  reg [43:0] calc_op0_fp_46_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1841" *)
  reg [43:0] calc_op0_fp_47_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1842" *)
  reg [43:0] calc_op0_fp_48_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1843" *)
  reg [43:0] calc_op0_fp_49_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1844" *)
  reg [43:0] calc_op0_fp_4_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1845" *)
  reg [43:0] calc_op0_fp_50_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1846" *)
  reg [43:0] calc_op0_fp_51_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1847" *)
  reg [43:0] calc_op0_fp_52_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1848" *)
  reg [43:0] calc_op0_fp_53_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1849" *)
  reg [43:0] calc_op0_fp_54_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1850" *)
  reg [43:0] calc_op0_fp_55_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1851" *)
  reg [43:0] calc_op0_fp_56_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1852" *)
  reg [43:0] calc_op0_fp_57_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1853" *)
  reg [43:0] calc_op0_fp_58_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1854" *)
  reg [43:0] calc_op0_fp_59_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1855" *)
  reg [43:0] calc_op0_fp_5_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1856" *)
  reg [43:0] calc_op0_fp_60_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1857" *)
  reg [43:0] calc_op0_fp_61_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1858" *)
  reg [43:0] calc_op0_fp_62_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1859" *)
  reg [43:0] calc_op0_fp_63_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1860" *)
  reg [43:0] calc_op0_fp_6_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1861" *)
  reg [43:0] calc_op0_fp_7_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1862" *)
  reg [43:0] calc_op0_fp_8_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1863" *)
  reg [43:0] calc_op0_fp_9_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1864" *)
  reg [37:0] calc_op0_int_0_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1865" *)
  reg [21:0] calc_op0_int_100_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1866" *)
  reg [21:0] calc_op0_int_101_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1867" *)
  reg [21:0] calc_op0_int_102_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1868" *)
  reg [21:0] calc_op0_int_103_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1869" *)
  reg [21:0] calc_op0_int_104_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1870" *)
  reg [21:0] calc_op0_int_105_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1871" *)
  reg [21:0] calc_op0_int_106_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1872" *)
  reg [21:0] calc_op0_int_107_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1873" *)
  reg [21:0] calc_op0_int_108_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1874" *)
  reg [21:0] calc_op0_int_109_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1875" *)
  reg [37:0] calc_op0_int_10_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1876" *)
  reg [21:0] calc_op0_int_110_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1877" *)
  reg [21:0] calc_op0_int_111_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1878" *)
  reg [21:0] calc_op0_int_112_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1879" *)
  reg [21:0] calc_op0_int_113_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1880" *)
  reg [21:0] calc_op0_int_114_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1881" *)
  reg [21:0] calc_op0_int_115_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1882" *)
  reg [21:0] calc_op0_int_116_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1883" *)
  reg [21:0] calc_op0_int_117_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1884" *)
  reg [21:0] calc_op0_int_118_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1885" *)
  reg [21:0] calc_op0_int_119_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1886" *)
  reg [37:0] calc_op0_int_11_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1887" *)
  reg [21:0] calc_op0_int_120_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1888" *)
  reg [21:0] calc_op0_int_121_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1889" *)
  reg [21:0] calc_op0_int_122_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1890" *)
  reg [21:0] calc_op0_int_123_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1891" *)
  reg [21:0] calc_op0_int_124_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1892" *)
  reg [21:0] calc_op0_int_125_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1893" *)
  reg [21:0] calc_op0_int_126_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1894" *)
  reg [21:0] calc_op0_int_127_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1895" *)
  reg [37:0] calc_op0_int_12_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1896" *)
  reg [37:0] calc_op0_int_13_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1897" *)
  reg [37:0] calc_op0_int_14_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1898" *)
  reg [37:0] calc_op0_int_15_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1899" *)
  reg [37:0] calc_op0_int_16_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1900" *)
  reg [37:0] calc_op0_int_17_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1901" *)
  reg [37:0] calc_op0_int_18_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1902" *)
  reg [37:0] calc_op0_int_19_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1903" *)
  reg [37:0] calc_op0_int_1_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1904" *)
  reg [37:0] calc_op0_int_20_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1905" *)
  reg [37:0] calc_op0_int_21_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1906" *)
  reg [37:0] calc_op0_int_22_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1907" *)
  reg [37:0] calc_op0_int_23_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1908" *)
  reg [37:0] calc_op0_int_24_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1909" *)
  reg [37:0] calc_op0_int_25_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1910" *)
  reg [37:0] calc_op0_int_26_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1911" *)
  reg [37:0] calc_op0_int_27_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1912" *)
  reg [37:0] calc_op0_int_28_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1913" *)
  reg [37:0] calc_op0_int_29_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1914" *)
  reg [37:0] calc_op0_int_2_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1915" *)
  reg [37:0] calc_op0_int_30_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1916" *)
  reg [37:0] calc_op0_int_31_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1917" *)
  reg [37:0] calc_op0_int_32_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1918" *)
  reg [37:0] calc_op0_int_33_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1919" *)
  reg [37:0] calc_op0_int_34_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1920" *)
  reg [37:0] calc_op0_int_35_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1921" *)
  reg [37:0] calc_op0_int_36_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1922" *)
  reg [37:0] calc_op0_int_37_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1923" *)
  reg [37:0] calc_op0_int_38_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1924" *)
  reg [37:0] calc_op0_int_39_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1925" *)
  reg [37:0] calc_op0_int_3_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1926" *)
  reg [37:0] calc_op0_int_40_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1927" *)
  reg [37:0] calc_op0_int_41_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1928" *)
  reg [37:0] calc_op0_int_42_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1929" *)
  reg [37:0] calc_op0_int_43_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1930" *)
  reg [37:0] calc_op0_int_44_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1931" *)
  reg [37:0] calc_op0_int_45_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1932" *)
  reg [37:0] calc_op0_int_46_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1933" *)
  reg [37:0] calc_op0_int_47_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1934" *)
  reg [37:0] calc_op0_int_48_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1935" *)
  reg [37:0] calc_op0_int_49_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1936" *)
  reg [37:0] calc_op0_int_4_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1937" *)
  reg [37:0] calc_op0_int_50_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1938" *)
  reg [37:0] calc_op0_int_51_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1939" *)
  reg [37:0] calc_op0_int_52_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1940" *)
  reg [37:0] calc_op0_int_53_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1941" *)
  reg [37:0] calc_op0_int_54_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1942" *)
  reg [37:0] calc_op0_int_55_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1943" *)
  reg [37:0] calc_op0_int_56_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1944" *)
  reg [37:0] calc_op0_int_57_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1945" *)
  reg [37:0] calc_op0_int_58_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1946" *)
  reg [37:0] calc_op0_int_59_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1947" *)
  reg [37:0] calc_op0_int_5_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1948" *)
  reg [37:0] calc_op0_int_60_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1949" *)
  reg [37:0] calc_op0_int_61_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1950" *)
  reg [37:0] calc_op0_int_62_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1951" *)
  reg [37:0] calc_op0_int_63_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1952" *)
  reg [21:0] calc_op0_int_64_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1953" *)
  reg [21:0] calc_op0_int_65_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1954" *)
  reg [21:0] calc_op0_int_66_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1955" *)
  reg [21:0] calc_op0_int_67_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1956" *)
  reg [21:0] calc_op0_int_68_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1957" *)
  reg [21:0] calc_op0_int_69_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1958" *)
  reg [37:0] calc_op0_int_6_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1959" *)
  reg [21:0] calc_op0_int_70_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1960" *)
  reg [21:0] calc_op0_int_71_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1961" *)
  reg [21:0] calc_op0_int_72_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1962" *)
  reg [21:0] calc_op0_int_73_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1963" *)
  reg [21:0] calc_op0_int_74_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1964" *)
  reg [21:0] calc_op0_int_75_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1965" *)
  reg [21:0] calc_op0_int_76_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1966" *)
  reg [21:0] calc_op0_int_77_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1967" *)
  reg [21:0] calc_op0_int_78_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1968" *)
  reg [21:0] calc_op0_int_79_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1969" *)
  reg [37:0] calc_op0_int_7_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1970" *)
  reg [21:0] calc_op0_int_80_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1971" *)
  reg [21:0] calc_op0_int_81_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1972" *)
  reg [21:0] calc_op0_int_82_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1973" *)
  reg [21:0] calc_op0_int_83_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1974" *)
  reg [21:0] calc_op0_int_84_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1975" *)
  reg [21:0] calc_op0_int_85_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1976" *)
  reg [21:0] calc_op0_int_86_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1977" *)
  reg [21:0] calc_op0_int_87_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1978" *)
  reg [21:0] calc_op0_int_88_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1979" *)
  reg [21:0] calc_op0_int_89_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1980" *)
  reg [37:0] calc_op0_int_8_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1981" *)
  reg [21:0] calc_op0_int_90_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1982" *)
  reg [21:0] calc_op0_int_91_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1983" *)
  reg [21:0] calc_op0_int_92_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1984" *)
  reg [21:0] calc_op0_int_93_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1985" *)
  reg [21:0] calc_op0_int_94_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1986" *)
  reg [21:0] calc_op0_int_95_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1987" *)
  reg [21:0] calc_op0_int_96_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1988" *)
  reg [21:0] calc_op0_int_97_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1989" *)
  reg [21:0] calc_op0_int_98_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1990" *)
  reg [21:0] calc_op0_int_99_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1991" *)
  reg [37:0] calc_op0_int_9_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1992" *)
  reg [47:0] calc_op1_fp_0_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1993" *)
  reg [47:0] calc_op1_fp_10_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1994" *)
  reg [47:0] calc_op1_fp_11_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1995" *)
  reg [47:0] calc_op1_fp_12_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1996" *)
  reg [47:0] calc_op1_fp_13_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1997" *)
  reg [47:0] calc_op1_fp_14_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1998" *)
  reg [47:0] calc_op1_fp_15_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1999" *)
  reg [47:0] calc_op1_fp_16_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2000" *)
  reg [47:0] calc_op1_fp_17_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2001" *)
  reg [47:0] calc_op1_fp_18_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2002" *)
  reg [47:0] calc_op1_fp_19_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2003" *)
  reg [47:0] calc_op1_fp_1_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2004" *)
  reg [47:0] calc_op1_fp_20_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2005" *)
  reg [47:0] calc_op1_fp_21_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2006" *)
  reg [47:0] calc_op1_fp_22_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2007" *)
  reg [47:0] calc_op1_fp_23_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2008" *)
  reg [47:0] calc_op1_fp_24_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2009" *)
  reg [47:0] calc_op1_fp_25_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2010" *)
  reg [47:0] calc_op1_fp_26_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2011" *)
  reg [47:0] calc_op1_fp_27_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2012" *)
  reg [47:0] calc_op1_fp_28_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2013" *)
  reg [47:0] calc_op1_fp_29_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2014" *)
  reg [47:0] calc_op1_fp_2_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2015" *)
  reg [47:0] calc_op1_fp_30_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2016" *)
  reg [47:0] calc_op1_fp_31_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2017" *)
  reg [47:0] calc_op1_fp_32_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2018" *)
  reg [47:0] calc_op1_fp_33_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2019" *)
  reg [47:0] calc_op1_fp_34_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2020" *)
  reg [47:0] calc_op1_fp_35_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2021" *)
  reg [47:0] calc_op1_fp_36_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2022" *)
  reg [47:0] calc_op1_fp_37_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2023" *)
  reg [47:0] calc_op1_fp_38_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2024" *)
  reg [47:0] calc_op1_fp_39_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2025" *)
  reg [47:0] calc_op1_fp_3_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2026" *)
  reg [47:0] calc_op1_fp_40_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2027" *)
  reg [47:0] calc_op1_fp_41_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2028" *)
  reg [47:0] calc_op1_fp_42_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2029" *)
  reg [47:0] calc_op1_fp_43_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2030" *)
  reg [47:0] calc_op1_fp_44_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2031" *)
  reg [47:0] calc_op1_fp_45_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2032" *)
  reg [47:0] calc_op1_fp_46_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2033" *)
  reg [47:0] calc_op1_fp_47_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2034" *)
  reg [47:0] calc_op1_fp_48_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2035" *)
  reg [47:0] calc_op1_fp_49_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2036" *)
  reg [47:0] calc_op1_fp_4_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2037" *)
  reg [47:0] calc_op1_fp_50_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2038" *)
  reg [47:0] calc_op1_fp_51_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2039" *)
  reg [47:0] calc_op1_fp_52_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2040" *)
  reg [47:0] calc_op1_fp_53_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2041" *)
  reg [47:0] calc_op1_fp_54_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2042" *)
  reg [47:0] calc_op1_fp_55_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2043" *)
  reg [47:0] calc_op1_fp_56_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2044" *)
  reg [47:0] calc_op1_fp_57_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2045" *)
  reg [47:0] calc_op1_fp_58_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2046" *)
  reg [47:0] calc_op1_fp_59_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2047" *)
  reg [47:0] calc_op1_fp_5_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2048" *)
  reg [47:0] calc_op1_fp_60_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2049" *)
  reg [47:0] calc_op1_fp_61_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2050" *)
  reg [47:0] calc_op1_fp_62_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2051" *)
  reg [47:0] calc_op1_fp_63_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2052" *)
  reg [47:0] calc_op1_fp_6_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2053" *)
  reg [47:0] calc_op1_fp_7_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2054" *)
  reg [47:0] calc_op1_fp_8_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2055" *)
  reg [47:0] calc_op1_fp_9_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2056" *)
  reg [47:0] calc_op1_int_0_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2057" *)
  reg [33:0] calc_op1_int_100_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2058" *)
  reg [33:0] calc_op1_int_101_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2059" *)
  reg [33:0] calc_op1_int_102_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2060" *)
  reg [33:0] calc_op1_int_103_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2061" *)
  reg [33:0] calc_op1_int_104_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2062" *)
  reg [33:0] calc_op1_int_105_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2063" *)
  reg [33:0] calc_op1_int_106_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2064" *)
  reg [33:0] calc_op1_int_107_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2065" *)
  reg [33:0] calc_op1_int_108_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2066" *)
  reg [33:0] calc_op1_int_109_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2067" *)
  reg [47:0] calc_op1_int_10_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2068" *)
  reg [33:0] calc_op1_int_110_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2069" *)
  reg [33:0] calc_op1_int_111_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2070" *)
  reg [33:0] calc_op1_int_112_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2071" *)
  reg [33:0] calc_op1_int_113_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2072" *)
  reg [33:0] calc_op1_int_114_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2073" *)
  reg [33:0] calc_op1_int_115_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2074" *)
  reg [33:0] calc_op1_int_116_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2075" *)
  reg [33:0] calc_op1_int_117_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2076" *)
  reg [33:0] calc_op1_int_118_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2077" *)
  reg [33:0] calc_op1_int_119_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2078" *)
  reg [47:0] calc_op1_int_11_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2079" *)
  reg [33:0] calc_op1_int_120_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2080" *)
  reg [33:0] calc_op1_int_121_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2081" *)
  reg [33:0] calc_op1_int_122_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2082" *)
  reg [33:0] calc_op1_int_123_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2083" *)
  reg [33:0] calc_op1_int_124_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2084" *)
  reg [33:0] calc_op1_int_125_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2085" *)
  reg [33:0] calc_op1_int_126_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2086" *)
  reg [33:0] calc_op1_int_127_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2087" *)
  reg [47:0] calc_op1_int_12_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2088" *)
  reg [47:0] calc_op1_int_13_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2089" *)
  reg [47:0] calc_op1_int_14_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2090" *)
  reg [47:0] calc_op1_int_15_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2091" *)
  reg [47:0] calc_op1_int_16_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2092" *)
  reg [47:0] calc_op1_int_17_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2093" *)
  reg [47:0] calc_op1_int_18_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2094" *)
  reg [47:0] calc_op1_int_19_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2095" *)
  reg [47:0] calc_op1_int_1_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2096" *)
  reg [47:0] calc_op1_int_20_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2097" *)
  reg [47:0] calc_op1_int_21_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2098" *)
  reg [47:0] calc_op1_int_22_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2099" *)
  reg [47:0] calc_op1_int_23_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2100" *)
  reg [47:0] calc_op1_int_24_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2101" *)
  reg [47:0] calc_op1_int_25_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2102" *)
  reg [47:0] calc_op1_int_26_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2103" *)
  reg [47:0] calc_op1_int_27_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2104" *)
  reg [47:0] calc_op1_int_28_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2105" *)
  reg [47:0] calc_op1_int_29_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2106" *)
  reg [47:0] calc_op1_int_2_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2107" *)
  reg [47:0] calc_op1_int_30_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2108" *)
  reg [47:0] calc_op1_int_31_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2109" *)
  reg [47:0] calc_op1_int_32_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2110" *)
  reg [47:0] calc_op1_int_33_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2111" *)
  reg [47:0] calc_op1_int_34_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2112" *)
  reg [47:0] calc_op1_int_35_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2113" *)
  reg [47:0] calc_op1_int_36_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2114" *)
  reg [47:0] calc_op1_int_37_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2115" *)
  reg [47:0] calc_op1_int_38_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2116" *)
  reg [47:0] calc_op1_int_39_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2117" *)
  reg [47:0] calc_op1_int_3_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2118" *)
  reg [47:0] calc_op1_int_40_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2119" *)
  reg [47:0] calc_op1_int_41_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2120" *)
  reg [47:0] calc_op1_int_42_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2121" *)
  reg [47:0] calc_op1_int_43_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2122" *)
  reg [47:0] calc_op1_int_44_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2123" *)
  reg [47:0] calc_op1_int_45_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2124" *)
  reg [47:0] calc_op1_int_46_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2125" *)
  reg [47:0] calc_op1_int_47_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2126" *)
  reg [47:0] calc_op1_int_48_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2127" *)
  reg [47:0] calc_op1_int_49_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2128" *)
  reg [47:0] calc_op1_int_4_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2129" *)
  reg [47:0] calc_op1_int_50_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2130" *)
  reg [47:0] calc_op1_int_51_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2131" *)
  reg [47:0] calc_op1_int_52_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2132" *)
  reg [47:0] calc_op1_int_53_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2133" *)
  reg [47:0] calc_op1_int_54_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2134" *)
  reg [47:0] calc_op1_int_55_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2135" *)
  reg [47:0] calc_op1_int_56_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2136" *)
  reg [47:0] calc_op1_int_57_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2137" *)
  reg [47:0] calc_op1_int_58_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2138" *)
  reg [47:0] calc_op1_int_59_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2139" *)
  reg [47:0] calc_op1_int_5_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2140" *)
  reg [47:0] calc_op1_int_60_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2141" *)
  reg [47:0] calc_op1_int_61_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2142" *)
  reg [47:0] calc_op1_int_62_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2143" *)
  reg [47:0] calc_op1_int_63_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2144" *)
  reg [33:0] calc_op1_int_64_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2145" *)
  reg [33:0] calc_op1_int_65_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2146" *)
  reg [33:0] calc_op1_int_66_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2147" *)
  reg [33:0] calc_op1_int_67_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2148" *)
  reg [33:0] calc_op1_int_68_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2149" *)
  reg [33:0] calc_op1_int_69_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2150" *)
  reg [47:0] calc_op1_int_6_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2151" *)
  reg [33:0] calc_op1_int_70_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2152" *)
  reg [33:0] calc_op1_int_71_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2153" *)
  reg [33:0] calc_op1_int_72_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2154" *)
  reg [33:0] calc_op1_int_73_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2155" *)
  reg [33:0] calc_op1_int_74_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2156" *)
  reg [33:0] calc_op1_int_75_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2157" *)
  reg [33:0] calc_op1_int_76_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2158" *)
  reg [33:0] calc_op1_int_77_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2159" *)
  reg [33:0] calc_op1_int_78_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2160" *)
  reg [33:0] calc_op1_int_79_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2161" *)
  reg [47:0] calc_op1_int_7_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2162" *)
  reg [33:0] calc_op1_int_80_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2163" *)
  reg [33:0] calc_op1_int_81_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2164" *)
  reg [33:0] calc_op1_int_82_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2165" *)
  reg [33:0] calc_op1_int_83_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2166" *)
  reg [33:0] calc_op1_int_84_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2167" *)
  reg [33:0] calc_op1_int_85_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2168" *)
  reg [33:0] calc_op1_int_86_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2169" *)
  reg [33:0] calc_op1_int_87_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2170" *)
  reg [33:0] calc_op1_int_88_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2171" *)
  reg [33:0] calc_op1_int_89_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2172" *)
  reg [47:0] calc_op1_int_8_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2173" *)
  reg [33:0] calc_op1_int_90_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2174" *)
  reg [33:0] calc_op1_int_91_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2175" *)
  reg [33:0] calc_op1_int_92_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2176" *)
  reg [33:0] calc_op1_int_93_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2177" *)
  reg [33:0] calc_op1_int_94_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2178" *)
  reg [33:0] calc_op1_int_95_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2179" *)
  reg [33:0] calc_op1_int_96_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2180" *)
  reg [33:0] calc_op1_int_97_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2181" *)
  reg [33:0] calc_op1_int_98_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2182" *)
  reg [33:0] calc_op1_int_99_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2183" *)
  reg [47:0] calc_op1_int_9_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1059" *)
  wire [63:0] calc_op1_vld_fp;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2184" *)
  reg [63:0] calc_op1_vld_fp_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1060" *)
  wire [127:0] calc_op1_vld_int;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2185" *)
  reg [127:0] calc_op1_vld_int_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1061" *)
  wire [63:0] calc_op_en_fp;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2186" *)
  reg [63:0] calc_op_en_fp_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1062" *)
  wire [127:0] calc_op_en_int;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2187" *)
  reg [127:0] calc_op_en_int_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1063" *)
  wire [47:0] calc_pout_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1064" *)
  wire [47:0] calc_pout_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1065" *)
  wire [47:0] calc_pout_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1066" *)
  wire [33:0] calc_pout_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1067" *)
  wire [33:0] calc_pout_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1068" *)
  wire [33:0] calc_pout_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1069" *)
  wire [33:0] calc_pout_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1070" *)
  wire [33:0] calc_pout_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1071" *)
  wire [33:0] calc_pout_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1072" *)
  wire [33:0] calc_pout_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1073" *)
  wire [33:0] calc_pout_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1074" *)
  wire [33:0] calc_pout_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1075" *)
  wire [33:0] calc_pout_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1076" *)
  wire [47:0] calc_pout_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1077" *)
  wire [33:0] calc_pout_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1078" *)
  wire [33:0] calc_pout_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1079" *)
  wire [33:0] calc_pout_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1080" *)
  wire [33:0] calc_pout_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1081" *)
  wire [33:0] calc_pout_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1082" *)
  wire [33:0] calc_pout_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1083" *)
  wire [33:0] calc_pout_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1084" *)
  wire [33:0] calc_pout_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1085" *)
  wire [33:0] calc_pout_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1086" *)
  wire [33:0] calc_pout_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1087" *)
  wire [47:0] calc_pout_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1088" *)
  wire [33:0] calc_pout_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1089" *)
  wire [33:0] calc_pout_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1090" *)
  wire [33:0] calc_pout_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1091" *)
  wire [33:0] calc_pout_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1092" *)
  wire [33:0] calc_pout_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1093" *)
  wire [33:0] calc_pout_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1094" *)
  wire [33:0] calc_pout_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1095" *)
  wire [33:0] calc_pout_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1096" *)
  wire [47:0] calc_pout_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1097" *)
  wire [47:0] calc_pout_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1098" *)
  wire [47:0] calc_pout_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1099" *)
  wire [47:0] calc_pout_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1100" *)
  wire [47:0] calc_pout_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1101" *)
  wire [47:0] calc_pout_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1102" *)
  wire [47:0] calc_pout_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1103" *)
  wire [47:0] calc_pout_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1104" *)
  wire [47:0] calc_pout_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1105" *)
  wire [47:0] calc_pout_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1106" *)
  wire [47:0] calc_pout_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1107" *)
  wire [47:0] calc_pout_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1108" *)
  wire [47:0] calc_pout_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1109" *)
  wire [47:0] calc_pout_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1110" *)
  wire [47:0] calc_pout_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1111" *)
  wire [47:0] calc_pout_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1112" *)
  wire [47:0] calc_pout_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1113" *)
  wire [47:0] calc_pout_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1114" *)
  wire [47:0] calc_pout_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1115" *)
  wire [47:0] calc_pout_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1116" *)
  wire [47:0] calc_pout_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1117" *)
  wire [47:0] calc_pout_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1118" *)
  wire [47:0] calc_pout_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1119" *)
  wire [47:0] calc_pout_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1120" *)
  wire [47:0] calc_pout_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1121" *)
  wire [47:0] calc_pout_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1122" *)
  wire [47:0] calc_pout_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1123" *)
  wire [47:0] calc_pout_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1124" *)
  wire [47:0] calc_pout_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1125" *)
  wire [47:0] calc_pout_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1126" *)
  wire [47:0] calc_pout_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1127" *)
  wire [47:0] calc_pout_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1128" *)
  wire [47:0] calc_pout_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1129" *)
  wire [47:0] calc_pout_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1130" *)
  wire [47:0] calc_pout_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1131" *)
  wire [47:0] calc_pout_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1132" *)
  wire [47:0] calc_pout_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1133" *)
  wire [47:0] calc_pout_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1134" *)
  wire [47:0] calc_pout_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1135" *)
  wire [47:0] calc_pout_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1136" *)
  wire [47:0] calc_pout_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1137" *)
  wire [47:0] calc_pout_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1138" *)
  wire [47:0] calc_pout_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1139" *)
  wire [47:0] calc_pout_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1140" *)
  wire [47:0] calc_pout_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1141" *)
  wire [47:0] calc_pout_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1142" *)
  wire [47:0] calc_pout_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1143" *)
  wire [47:0] calc_pout_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1144" *)
  wire [47:0] calc_pout_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1145" *)
  wire [47:0] calc_pout_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1146" *)
  wire [47:0] calc_pout_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1147" *)
  wire [47:0] calc_pout_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1148" *)
  wire [47:0] calc_pout_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1149" *)
  wire [47:0] calc_pout_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1150" *)
  wire [47:0] calc_pout_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1151" *)
  wire [47:0] calc_pout_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1152" *)
  wire [33:0] calc_pout_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1153" *)
  wire [33:0] calc_pout_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1154" *)
  wire [33:0] calc_pout_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1155" *)
  wire [33:0] calc_pout_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1156" *)
  wire [33:0] calc_pout_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1157" *)
  wire [33:0] calc_pout_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1158" *)
  wire [47:0] calc_pout_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1159" *)
  wire [33:0] calc_pout_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1160" *)
  wire [33:0] calc_pout_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1161" *)
  wire [33:0] calc_pout_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1162" *)
  wire [33:0] calc_pout_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1163" *)
  wire [33:0] calc_pout_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1164" *)
  wire [33:0] calc_pout_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1165" *)
  wire [33:0] calc_pout_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1166" *)
  wire [33:0] calc_pout_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1167" *)
  wire [33:0] calc_pout_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1168" *)
  wire [33:0] calc_pout_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1169" *)
  wire [47:0] calc_pout_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1170" *)
  wire [33:0] calc_pout_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1171" *)
  wire [33:0] calc_pout_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1172" *)
  wire [33:0] calc_pout_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1173" *)
  wire [33:0] calc_pout_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1174" *)
  wire [33:0] calc_pout_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1175" *)
  wire [33:0] calc_pout_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1176" *)
  wire [33:0] calc_pout_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1177" *)
  wire [33:0] calc_pout_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1178" *)
  wire [33:0] calc_pout_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1179" *)
  wire [33:0] calc_pout_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1180" *)
  wire [47:0] calc_pout_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1181" *)
  wire [33:0] calc_pout_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1182" *)
  wire [33:0] calc_pout_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1183" *)
  wire [33:0] calc_pout_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1184" *)
  wire [33:0] calc_pout_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1185" *)
  wire [33:0] calc_pout_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1186" *)
  wire [33:0] calc_pout_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1187" *)
  wire [33:0] calc_pout_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1188" *)
  wire [33:0] calc_pout_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1189" *)
  wire [33:0] calc_pout_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1190" *)
  wire [33:0] calc_pout_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1191" *)
  wire [47:0] calc_pout_fp_0_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1192" *)
  wire [47:0] calc_pout_fp_0_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1193" *)
  wire [47:0] calc_pout_fp_10_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1194" *)
  wire [47:0] calc_pout_fp_10_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1195" *)
  wire [47:0] calc_pout_fp_11_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1196" *)
  wire [47:0] calc_pout_fp_11_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1197" *)
  wire [47:0] calc_pout_fp_12_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1198" *)
  wire [47:0] calc_pout_fp_12_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1199" *)
  wire [47:0] calc_pout_fp_13_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1200" *)
  wire [47:0] calc_pout_fp_13_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1201" *)
  wire [47:0] calc_pout_fp_14_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1202" *)
  wire [47:0] calc_pout_fp_14_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1203" *)
  wire [47:0] calc_pout_fp_15_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1204" *)
  wire [47:0] calc_pout_fp_15_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1205" *)
  wire [47:0] calc_pout_fp_16_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1206" *)
  wire [47:0] calc_pout_fp_16_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1207" *)
  wire [47:0] calc_pout_fp_17_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1208" *)
  wire [47:0] calc_pout_fp_17_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1209" *)
  wire [47:0] calc_pout_fp_18_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1210" *)
  wire [47:0] calc_pout_fp_18_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1211" *)
  wire [47:0] calc_pout_fp_19_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1212" *)
  wire [47:0] calc_pout_fp_19_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1213" *)
  wire [47:0] calc_pout_fp_1_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1214" *)
  wire [47:0] calc_pout_fp_1_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1215" *)
  wire [47:0] calc_pout_fp_20_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1216" *)
  wire [47:0] calc_pout_fp_20_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1217" *)
  wire [47:0] calc_pout_fp_21_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1218" *)
  wire [47:0] calc_pout_fp_21_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1219" *)
  wire [47:0] calc_pout_fp_22_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1220" *)
  wire [47:0] calc_pout_fp_22_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1221" *)
  wire [47:0] calc_pout_fp_23_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1222" *)
  wire [47:0] calc_pout_fp_23_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1223" *)
  wire [47:0] calc_pout_fp_24_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1224" *)
  wire [47:0] calc_pout_fp_24_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1225" *)
  wire [47:0] calc_pout_fp_25_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1226" *)
  wire [47:0] calc_pout_fp_25_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1227" *)
  wire [47:0] calc_pout_fp_26_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1228" *)
  wire [47:0] calc_pout_fp_26_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1229" *)
  wire [47:0] calc_pout_fp_27_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1230" *)
  wire [47:0] calc_pout_fp_27_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1231" *)
  wire [47:0] calc_pout_fp_28_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1232" *)
  wire [47:0] calc_pout_fp_28_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1233" *)
  wire [47:0] calc_pout_fp_29_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1234" *)
  wire [47:0] calc_pout_fp_29_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1235" *)
  wire [47:0] calc_pout_fp_2_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1236" *)
  wire [47:0] calc_pout_fp_2_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1237" *)
  wire [47:0] calc_pout_fp_30_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1238" *)
  wire [47:0] calc_pout_fp_30_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1239" *)
  wire [47:0] calc_pout_fp_31_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1240" *)
  wire [47:0] calc_pout_fp_31_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1241" *)
  wire [47:0] calc_pout_fp_32_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1242" *)
  wire [47:0] calc_pout_fp_32_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1243" *)
  wire [47:0] calc_pout_fp_33_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1244" *)
  wire [47:0] calc_pout_fp_33_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1245" *)
  wire [47:0] calc_pout_fp_34_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1246" *)
  wire [47:0] calc_pout_fp_34_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1247" *)
  wire [47:0] calc_pout_fp_35_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1248" *)
  wire [47:0] calc_pout_fp_35_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1249" *)
  wire [47:0] calc_pout_fp_36_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1250" *)
  wire [47:0] calc_pout_fp_36_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1251" *)
  wire [47:0] calc_pout_fp_37_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1252" *)
  wire [47:0] calc_pout_fp_37_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1253" *)
  wire [47:0] calc_pout_fp_38_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1254" *)
  wire [47:0] calc_pout_fp_38_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1255" *)
  wire [47:0] calc_pout_fp_39_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1256" *)
  wire [47:0] calc_pout_fp_39_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1257" *)
  wire [47:0] calc_pout_fp_3_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1258" *)
  wire [47:0] calc_pout_fp_3_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1259" *)
  wire [47:0] calc_pout_fp_40_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1260" *)
  wire [47:0] calc_pout_fp_40_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1261" *)
  wire [47:0] calc_pout_fp_41_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1262" *)
  wire [47:0] calc_pout_fp_41_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1263" *)
  wire [47:0] calc_pout_fp_42_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1264" *)
  wire [47:0] calc_pout_fp_42_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1265" *)
  wire [47:0] calc_pout_fp_43_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1266" *)
  wire [47:0] calc_pout_fp_43_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1267" *)
  wire [47:0] calc_pout_fp_44_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1268" *)
  wire [47:0] calc_pout_fp_44_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1269" *)
  wire [47:0] calc_pout_fp_45_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1270" *)
  wire [47:0] calc_pout_fp_45_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1271" *)
  wire [47:0] calc_pout_fp_46_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1272" *)
  wire [47:0] calc_pout_fp_46_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1273" *)
  wire [47:0] calc_pout_fp_47_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1274" *)
  wire [47:0] calc_pout_fp_47_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1275" *)
  wire [47:0] calc_pout_fp_48_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1276" *)
  wire [47:0] calc_pout_fp_48_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1277" *)
  wire [47:0] calc_pout_fp_49_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1278" *)
  wire [47:0] calc_pout_fp_49_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1279" *)
  wire [47:0] calc_pout_fp_4_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1280" *)
  wire [47:0] calc_pout_fp_4_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1281" *)
  wire [47:0] calc_pout_fp_50_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1282" *)
  wire [47:0] calc_pout_fp_50_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1283" *)
  wire [47:0] calc_pout_fp_51_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1284" *)
  wire [47:0] calc_pout_fp_51_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1285" *)
  wire [47:0] calc_pout_fp_52_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1286" *)
  wire [47:0] calc_pout_fp_52_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1287" *)
  wire [47:0] calc_pout_fp_53_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1288" *)
  wire [47:0] calc_pout_fp_53_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1289" *)
  wire [47:0] calc_pout_fp_54_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1290" *)
  wire [47:0] calc_pout_fp_54_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1291" *)
  wire [47:0] calc_pout_fp_55_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1292" *)
  wire [47:0] calc_pout_fp_55_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1293" *)
  wire [47:0] calc_pout_fp_56_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1294" *)
  wire [47:0] calc_pout_fp_56_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1295" *)
  wire [47:0] calc_pout_fp_57_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1296" *)
  wire [47:0] calc_pout_fp_57_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1297" *)
  wire [47:0] calc_pout_fp_58_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1298" *)
  wire [47:0] calc_pout_fp_58_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1299" *)
  wire [47:0] calc_pout_fp_59_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1300" *)
  wire [47:0] calc_pout_fp_59_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1301" *)
  wire [47:0] calc_pout_fp_5_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1302" *)
  wire [47:0] calc_pout_fp_5_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1303" *)
  wire [47:0] calc_pout_fp_60_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1304" *)
  wire [47:0] calc_pout_fp_60_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1305" *)
  wire [47:0] calc_pout_fp_61_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1306" *)
  wire [47:0] calc_pout_fp_61_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1307" *)
  wire [47:0] calc_pout_fp_62_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1308" *)
  wire [47:0] calc_pout_fp_62_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1309" *)
  wire [47:0] calc_pout_fp_63_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1310" *)
  wire [47:0] calc_pout_fp_63_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1311" *)
  wire [47:0] calc_pout_fp_6_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1312" *)
  wire [47:0] calc_pout_fp_6_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1313" *)
  wire [47:0] calc_pout_fp_7_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1314" *)
  wire [47:0] calc_pout_fp_7_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1315" *)
  wire [47:0] calc_pout_fp_8_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1316" *)
  wire [47:0] calc_pout_fp_8_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1317" *)
  wire [47:0] calc_pout_fp_9_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1318" *)
  wire [47:0] calc_pout_fp_9_sum_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1319" *)
  wire [63:0] calc_pout_fp_vld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1320" *)
  wire [47:0] calc_pout_int_0_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1321" *)
  wire [33:0] calc_pout_int_100_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1322" *)
  wire [33:0] calc_pout_int_101_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1323" *)
  wire [33:0] calc_pout_int_102_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1324" *)
  wire [33:0] calc_pout_int_103_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1325" *)
  wire [33:0] calc_pout_int_104_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1326" *)
  wire [33:0] calc_pout_int_105_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1327" *)
  wire [33:0] calc_pout_int_106_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1328" *)
  wire [33:0] calc_pout_int_107_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1329" *)
  wire [33:0] calc_pout_int_108_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1330" *)
  wire [33:0] calc_pout_int_109_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1331" *)
  wire [47:0] calc_pout_int_10_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1332" *)
  wire [33:0] calc_pout_int_110_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1333" *)
  wire [33:0] calc_pout_int_111_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1334" *)
  wire [33:0] calc_pout_int_112_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1335" *)
  wire [33:0] calc_pout_int_113_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1336" *)
  wire [33:0] calc_pout_int_114_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1337" *)
  wire [33:0] calc_pout_int_115_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1338" *)
  wire [33:0] calc_pout_int_116_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1339" *)
  wire [33:0] calc_pout_int_117_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1340" *)
  wire [33:0] calc_pout_int_118_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1341" *)
  wire [33:0] calc_pout_int_119_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1342" *)
  wire [47:0] calc_pout_int_11_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1343" *)
  wire [33:0] calc_pout_int_120_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1344" *)
  wire [33:0] calc_pout_int_121_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1345" *)
  wire [33:0] calc_pout_int_122_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1346" *)
  wire [33:0] calc_pout_int_123_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1347" *)
  wire [33:0] calc_pout_int_124_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1348" *)
  wire [33:0] calc_pout_int_125_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1349" *)
  wire [33:0] calc_pout_int_126_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1350" *)
  wire [33:0] calc_pout_int_127_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1351" *)
  wire [47:0] calc_pout_int_12_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1352" *)
  wire [47:0] calc_pout_int_13_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1353" *)
  wire [47:0] calc_pout_int_14_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1354" *)
  wire [47:0] calc_pout_int_15_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1355" *)
  wire [47:0] calc_pout_int_16_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1356" *)
  wire [47:0] calc_pout_int_17_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1357" *)
  wire [47:0] calc_pout_int_18_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1358" *)
  wire [47:0] calc_pout_int_19_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1359" *)
  wire [47:0] calc_pout_int_1_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1360" *)
  wire [47:0] calc_pout_int_20_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1361" *)
  wire [47:0] calc_pout_int_21_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1362" *)
  wire [47:0] calc_pout_int_22_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1363" *)
  wire [47:0] calc_pout_int_23_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1364" *)
  wire [47:0] calc_pout_int_24_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1365" *)
  wire [47:0] calc_pout_int_25_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1366" *)
  wire [47:0] calc_pout_int_26_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1367" *)
  wire [47:0] calc_pout_int_27_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1368" *)
  wire [47:0] calc_pout_int_28_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1369" *)
  wire [47:0] calc_pout_int_29_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1370" *)
  wire [47:0] calc_pout_int_2_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1371" *)
  wire [47:0] calc_pout_int_30_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1372" *)
  wire [47:0] calc_pout_int_31_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1373" *)
  wire [47:0] calc_pout_int_32_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1374" *)
  wire [47:0] calc_pout_int_33_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1375" *)
  wire [47:0] calc_pout_int_34_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1376" *)
  wire [47:0] calc_pout_int_35_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1377" *)
  wire [47:0] calc_pout_int_36_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1378" *)
  wire [47:0] calc_pout_int_37_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1379" *)
  wire [47:0] calc_pout_int_38_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1380" *)
  wire [47:0] calc_pout_int_39_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1381" *)
  wire [47:0] calc_pout_int_3_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1382" *)
  wire [47:0] calc_pout_int_40_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1383" *)
  wire [47:0] calc_pout_int_41_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1384" *)
  wire [47:0] calc_pout_int_42_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1385" *)
  wire [47:0] calc_pout_int_43_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1386" *)
  wire [47:0] calc_pout_int_44_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1387" *)
  wire [47:0] calc_pout_int_45_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1388" *)
  wire [47:0] calc_pout_int_46_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1389" *)
  wire [47:0] calc_pout_int_47_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1390" *)
  wire [47:0] calc_pout_int_48_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1391" *)
  wire [47:0] calc_pout_int_49_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1392" *)
  wire [47:0] calc_pout_int_4_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1393" *)
  wire [47:0] calc_pout_int_50_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1394" *)
  wire [47:0] calc_pout_int_51_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1395" *)
  wire [47:0] calc_pout_int_52_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1396" *)
  wire [47:0] calc_pout_int_53_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1397" *)
  wire [47:0] calc_pout_int_54_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1398" *)
  wire [47:0] calc_pout_int_55_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1399" *)
  wire [47:0] calc_pout_int_56_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1400" *)
  wire [47:0] calc_pout_int_57_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1401" *)
  wire [47:0] calc_pout_int_58_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1402" *)
  wire [47:0] calc_pout_int_59_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1403" *)
  wire [47:0] calc_pout_int_5_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1404" *)
  wire [47:0] calc_pout_int_60_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1405" *)
  wire [47:0] calc_pout_int_61_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1406" *)
  wire [47:0] calc_pout_int_62_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1407" *)
  wire [47:0] calc_pout_int_63_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1408" *)
  wire [33:0] calc_pout_int_64_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1409" *)
  wire [33:0] calc_pout_int_65_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1410" *)
  wire [33:0] calc_pout_int_66_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1411" *)
  wire [33:0] calc_pout_int_67_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1412" *)
  wire [33:0] calc_pout_int_68_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1413" *)
  wire [33:0] calc_pout_int_69_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1414" *)
  wire [47:0] calc_pout_int_6_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1415" *)
  wire [33:0] calc_pout_int_70_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1416" *)
  wire [33:0] calc_pout_int_71_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1417" *)
  wire [33:0] calc_pout_int_72_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1418" *)
  wire [33:0] calc_pout_int_73_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1419" *)
  wire [33:0] calc_pout_int_74_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1420" *)
  wire [33:0] calc_pout_int_75_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1421" *)
  wire [33:0] calc_pout_int_76_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1422" *)
  wire [33:0] calc_pout_int_77_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1423" *)
  wire [33:0] calc_pout_int_78_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1424" *)
  wire [33:0] calc_pout_int_79_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1425" *)
  wire [47:0] calc_pout_int_7_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1426" *)
  wire [33:0] calc_pout_int_80_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1427" *)
  wire [33:0] calc_pout_int_81_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1428" *)
  wire [33:0] calc_pout_int_82_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1429" *)
  wire [33:0] calc_pout_int_83_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1430" *)
  wire [33:0] calc_pout_int_84_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1431" *)
  wire [33:0] calc_pout_int_85_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1432" *)
  wire [33:0] calc_pout_int_86_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1433" *)
  wire [33:0] calc_pout_int_87_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1434" *)
  wire [33:0] calc_pout_int_88_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1435" *)
  wire [33:0] calc_pout_int_89_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1436" *)
  wire [47:0] calc_pout_int_8_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1437" *)
  wire [33:0] calc_pout_int_90_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1438" *)
  wire [33:0] calc_pout_int_91_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1439" *)
  wire [33:0] calc_pout_int_92_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1440" *)
  wire [33:0] calc_pout_int_93_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1441" *)
  wire [33:0] calc_pout_int_94_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1442" *)
  wire [33:0] calc_pout_int_95_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1443" *)
  wire [33:0] calc_pout_int_96_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1444" *)
  wire [33:0] calc_pout_int_97_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1445" *)
  wire [33:0] calc_pout_int_98_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1446" *)
  wire [33:0] calc_pout_int_99_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1447" *)
  wire [47:0] calc_pout_int_9_sum;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1448" *)
  wire [127:0] calc_pout_int_vld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1449" *)
  wire [15:0] calc_ram_sel_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1450" *)
  wire [767:0] calc_ram_sel_0_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1451" *)
  wire [15:0] calc_ram_sel_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1452" *)
  wire [767:0] calc_ram_sel_1_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1453" *)
  wire [15:0] calc_ram_sel_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1454" *)
  wire [767:0] calc_ram_sel_2_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1455" *)
  wire [15:0] calc_ram_sel_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1456" *)
  wire [767:0] calc_ram_sel_3_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1457" *)
  wire [15:0] calc_ram_sel_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1458" *)
  wire [543:0] calc_ram_sel_4_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1459" *)
  wire [15:0] calc_ram_sel_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1460" *)
  wire [543:0] calc_ram_sel_5_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1461" *)
  wire [15:0] calc_ram_sel_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1462" *)
  wire [543:0] calc_ram_sel_6_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1463" *)
  wire [15:0] calc_ram_sel_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1464" *)
  wire [543:0] calc_ram_sel_7_ext;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1465" *)
  wire [7:0] calc_rd_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1466" *)
  wire calc_stripe_end;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2188" *)
  reg calc_stripe_end_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2189" *)
  reg calc_stripe_end_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2190" *)
  reg calc_stripe_end_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2191" *)
  reg calc_stripe_end_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2192" *)
  reg calc_stripe_end_d5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1467" *)
  wire calc_stripe_end_out;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2193" *)
  reg calc_valid;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1468" *)
  wire calc_valid_d0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2194" *)
  reg calc_valid_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2195" *)
  reg calc_valid_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2196" *)
  reg calc_valid_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2197" *)
  reg calc_valid_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1469" *)
  wire calc_valid_fw_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2198" *)
  reg calc_valid_fw_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2199" *)
  reg calc_valid_fw_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2200" *)
  reg calc_valid_fw_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1471" *)
  wire calc_valid_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2201" *)
  wire [7:0] calc_wr_en;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2202" *)
  reg [7:0] calc_wr_en_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2203" *)
  reg [7:0] calc_wr_en_d2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2204" *)
  reg [7:0] calc_wr_en_d3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2205" *)
  reg [7:0] calc_wr_en_d4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1472" *)
  wire [7:0] calc_wr_en_out;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:95" *)
  input [191:0] cfg_in_en_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:96" *)
  input [24:0] cfg_is_fp;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:97" *)
  input [24:0] cfg_is_int;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:98" *)
  input [126:0] cfg_is_int8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:99" *)
  input [95:0] cfg_is_wg;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:100" *)
  input [639:0] cfg_truncate;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1473" *)
  wire [4:0] cfg_truncate_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1474" *)
  wire [4:0] cfg_truncate_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1475" *)
  wire [4:0] cfg_truncate_10;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1476" *)
  wire [4:0] cfg_truncate_100;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1477" *)
  wire [4:0] cfg_truncate_101;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1478" *)
  wire [4:0] cfg_truncate_102;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1479" *)
  wire [4:0] cfg_truncate_103;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1480" *)
  wire [4:0] cfg_truncate_104;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1481" *)
  wire [4:0] cfg_truncate_105;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1482" *)
  wire [4:0] cfg_truncate_106;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1483" *)
  wire [4:0] cfg_truncate_107;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1484" *)
  wire [4:0] cfg_truncate_108;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1485" *)
  wire [4:0] cfg_truncate_109;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1486" *)
  wire [4:0] cfg_truncate_11;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1487" *)
  wire [4:0] cfg_truncate_110;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1488" *)
  wire [4:0] cfg_truncate_111;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1489" *)
  wire [4:0] cfg_truncate_112;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1490" *)
  wire [4:0] cfg_truncate_113;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1491" *)
  wire [4:0] cfg_truncate_114;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1492" *)
  wire [4:0] cfg_truncate_115;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1493" *)
  wire [4:0] cfg_truncate_116;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1494" *)
  wire [4:0] cfg_truncate_117;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1495" *)
  wire [4:0] cfg_truncate_118;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1496" *)
  wire [4:0] cfg_truncate_119;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1497" *)
  wire [4:0] cfg_truncate_12;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1498" *)
  wire [4:0] cfg_truncate_120;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1499" *)
  wire [4:0] cfg_truncate_121;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1500" *)
  wire [4:0] cfg_truncate_122;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1501" *)
  wire [4:0] cfg_truncate_123;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1502" *)
  wire [4:0] cfg_truncate_124;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1503" *)
  wire [4:0] cfg_truncate_125;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1504" *)
  wire [4:0] cfg_truncate_126;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1505" *)
  wire [4:0] cfg_truncate_127;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1506" *)
  wire [4:0] cfg_truncate_13;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1507" *)
  wire [4:0] cfg_truncate_14;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1508" *)
  wire [4:0] cfg_truncate_15;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1509" *)
  wire [4:0] cfg_truncate_16;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1510" *)
  wire [4:0] cfg_truncate_17;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1511" *)
  wire [4:0] cfg_truncate_18;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1512" *)
  wire [4:0] cfg_truncate_19;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1513" *)
  wire [4:0] cfg_truncate_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1514" *)
  wire [4:0] cfg_truncate_20;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1515" *)
  wire [4:0] cfg_truncate_21;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1516" *)
  wire [4:0] cfg_truncate_22;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1517" *)
  wire [4:0] cfg_truncate_23;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1518" *)
  wire [4:0] cfg_truncate_24;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1519" *)
  wire [4:0] cfg_truncate_25;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1520" *)
  wire [4:0] cfg_truncate_26;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1521" *)
  wire [4:0] cfg_truncate_27;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1522" *)
  wire [4:0] cfg_truncate_28;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1523" *)
  wire [4:0] cfg_truncate_29;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1524" *)
  wire [4:0] cfg_truncate_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1525" *)
  wire [4:0] cfg_truncate_30;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1526" *)
  wire [4:0] cfg_truncate_31;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1527" *)
  wire [4:0] cfg_truncate_32;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1528" *)
  wire [4:0] cfg_truncate_33;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1529" *)
  wire [4:0] cfg_truncate_34;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1530" *)
  wire [4:0] cfg_truncate_35;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1531" *)
  wire [4:0] cfg_truncate_36;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1532" *)
  wire [4:0] cfg_truncate_37;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1533" *)
  wire [4:0] cfg_truncate_38;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1534" *)
  wire [4:0] cfg_truncate_39;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1535" *)
  wire [4:0] cfg_truncate_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1536" *)
  wire [4:0] cfg_truncate_40;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1537" *)
  wire [4:0] cfg_truncate_41;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1538" *)
  wire [4:0] cfg_truncate_42;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1539" *)
  wire [4:0] cfg_truncate_43;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1540" *)
  wire [4:0] cfg_truncate_44;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1541" *)
  wire [4:0] cfg_truncate_45;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1542" *)
  wire [4:0] cfg_truncate_46;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1543" *)
  wire [4:0] cfg_truncate_47;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1544" *)
  wire [4:0] cfg_truncate_48;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1545" *)
  wire [4:0] cfg_truncate_49;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1546" *)
  wire [4:0] cfg_truncate_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1547" *)
  wire [4:0] cfg_truncate_50;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1548" *)
  wire [4:0] cfg_truncate_51;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1549" *)
  wire [4:0] cfg_truncate_52;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1550" *)
  wire [4:0] cfg_truncate_53;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1551" *)
  wire [4:0] cfg_truncate_54;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1552" *)
  wire [4:0] cfg_truncate_55;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1553" *)
  wire [4:0] cfg_truncate_56;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1554" *)
  wire [4:0] cfg_truncate_57;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1555" *)
  wire [4:0] cfg_truncate_58;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1556" *)
  wire [4:0] cfg_truncate_59;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1557" *)
  wire [4:0] cfg_truncate_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1558" *)
  wire [4:0] cfg_truncate_60;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1559" *)
  wire [4:0] cfg_truncate_61;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1560" *)
  wire [4:0] cfg_truncate_62;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1561" *)
  wire [4:0] cfg_truncate_63;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1562" *)
  wire [4:0] cfg_truncate_64;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1563" *)
  wire [4:0] cfg_truncate_65;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1564" *)
  wire [4:0] cfg_truncate_66;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1565" *)
  wire [4:0] cfg_truncate_67;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1566" *)
  wire [4:0] cfg_truncate_68;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1567" *)
  wire [4:0] cfg_truncate_69;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1568" *)
  wire [4:0] cfg_truncate_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1569" *)
  wire [4:0] cfg_truncate_70;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1570" *)
  wire [4:0] cfg_truncate_71;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1571" *)
  wire [4:0] cfg_truncate_72;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1572" *)
  wire [4:0] cfg_truncate_73;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1573" *)
  wire [4:0] cfg_truncate_74;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1574" *)
  wire [4:0] cfg_truncate_75;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1575" *)
  wire [4:0] cfg_truncate_76;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1576" *)
  wire [4:0] cfg_truncate_77;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1577" *)
  wire [4:0] cfg_truncate_78;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1578" *)
  wire [4:0] cfg_truncate_79;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1579" *)
  wire [4:0] cfg_truncate_8;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1580" *)
  wire [4:0] cfg_truncate_80;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1581" *)
  wire [4:0] cfg_truncate_81;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1582" *)
  wire [4:0] cfg_truncate_82;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1583" *)
  wire [4:0] cfg_truncate_83;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1584" *)
  wire [4:0] cfg_truncate_84;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1585" *)
  wire [4:0] cfg_truncate_85;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1586" *)
  wire [4:0] cfg_truncate_86;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1587" *)
  wire [4:0] cfg_truncate_87;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1588" *)
  wire [4:0] cfg_truncate_88;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1589" *)
  wire [4:0] cfg_truncate_89;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1590" *)
  wire [4:0] cfg_truncate_9;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1591" *)
  wire [4:0] cfg_truncate_90;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1592" *)
  wire [4:0] cfg_truncate_91;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1593" *)
  wire [4:0] cfg_truncate_92;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1594" *)
  wire [4:0] cfg_truncate_93;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1595" *)
  wire [4:0] cfg_truncate_94;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1596" *)
  wire [4:0] cfg_truncate_95;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1597" *)
  wire [4:0] cfg_truncate_96;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1598" *)
  wire [4:0] cfg_truncate_97;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1599" *)
  wire [4:0] cfg_truncate_98;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1600" *)
  wire [4:0] cfg_truncate_99;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:133" *)
  output [511:0] dlv_data_0;
  reg [511:0] dlv_data_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2207" *)
  wire [511:0] dlv_data_0_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:134" *)
  output [511:0] dlv_data_1;
  reg [511:0] dlv_data_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2209" *)
  wire [511:0] dlv_data_1_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:135" *)
  output [511:0] dlv_data_2;
  reg [511:0] dlv_data_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2211" *)
  wire [511:0] dlv_data_2_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:136" *)
  output [511:0] dlv_data_3;
  reg [511:0] dlv_data_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2213" *)
  wire [511:0] dlv_data_3_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:137" *)
  output [511:0] dlv_data_4;
  reg [511:0] dlv_data_4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2215" *)
  wire [511:0] dlv_data_4_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:138" *)
  output [511:0] dlv_data_5;
  reg [511:0] dlv_data_5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2217" *)
  wire [511:0] dlv_data_5_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:139" *)
  output [511:0] dlv_data_6;
  reg [511:0] dlv_data_6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2219" *)
  wire [511:0] dlv_data_6_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:140" *)
  output [511:0] dlv_data_7;
  reg [511:0] dlv_data_7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2221" *)
  wire [511:0] dlv_data_7_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2222" *)
  reg dlv_layer_end;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:141" *)
  output [7:0] dlv_mask;
  reg [7:0] dlv_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:142" *)
  output [1:0] dlv_pd;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1601" *)
  wire [127:0] dlv_sat_bit;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2224" *)
  reg [127:0] dlv_sat_bit_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1602" *)
  wire dlv_sat_clr;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2225" *)
  reg dlv_sat_clr_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1603" *)
  wire dlv_sat_end;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2226" *)
  reg dlv_sat_end_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2227" *)
  reg dlv_sat_vld_d1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2228" *)
  reg dlv_stripe_end;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:143" *)
  output dlv_valid;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:144" *)
  output [31:0] dp2reg_sat_count;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:101" *)
  input [175:0] mac_a2accu_data0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:102" *)
  input [175:0] mac_a2accu_data1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:103" *)
  input [175:0] mac_a2accu_data2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:104" *)
  input [175:0] mac_a2accu_data3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:105" *)
  input [175:0] mac_a2accu_data4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:106" *)
  input [175:0] mac_a2accu_data5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:107" *)
  input [175:0] mac_a2accu_data6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:108" *)
  input [175:0] mac_a2accu_data7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:109" *)
  input [7:0] mac_a2accu_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:110" *)
  input [7:0] mac_a2accu_mode;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:111" *)
  input mac_a2accu_pvld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:112" *)
  input [175:0] mac_b2accu_data0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:113" *)
  input [175:0] mac_b2accu_data1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:114" *)
  input [175:0] mac_b2accu_data2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:115" *)
  input [175:0] mac_b2accu_data3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:116" *)
  input [175:0] mac_b2accu_data4;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:117" *)
  input [175:0] mac_b2accu_data5;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:118" *)
  input [175:0] mac_b2accu_data6;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:119" *)
  input [175:0] mac_b2accu_data7;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:120" *)
  input [7:0] mac_b2accu_mask;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:121" *)
  input [7:0] mac_b2accu_mode;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:122" *)
  input mac_b2accu_pvld;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:78" *)
  input nvdla_cell_clk_0;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:79" *)
  input nvdla_cell_clk_1;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:80" *)
  input nvdla_cell_clk_2;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:81" *)
  input nvdla_cell_clk_3;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:82" *)
  input nvdla_core_clk;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:83" *)
  input nvdla_core_rstn;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2230" *)
  wire sat_carry;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2231" *)
  reg [31:0] sat_count;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2232" *)
  wire [31:0] sat_count_inc;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1604" *)
  wire [31:0] sat_count_w;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:1605" *)
  wire sat_reg_en;
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2233" *)
  wire [7:0] sat_sum;
  assign _0469_ = dlv_sat_bit_d1[127] + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[126];
  assign _0470_ = _0469_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[125];
  assign _0471_ = _0470_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[124];
  assign _0472_ = _0471_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[123];
  assign _0473_ = _0472_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[122];
  assign _0474_ = _0473_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[121];
  assign _0475_ = _0474_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[120];
  assign _0476_ = _0475_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[119];
  assign _0477_ = _0476_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[118];
  assign _0478_ = _0477_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[117];
  assign _0479_ = _0478_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[116];
  assign _0480_ = _0479_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[115];
  assign _0481_ = _0480_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[114];
  assign _0482_ = _0481_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[113];
  assign _0483_ = _0482_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[112];
  assign _0484_ = _0483_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[111];
  assign _0485_ = _0484_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[110];
  assign _0486_ = _0485_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[109];
  assign _0487_ = _0486_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[108];
  assign _0488_ = _0487_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[107];
  assign _0489_ = _0488_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[106];
  assign _0490_ = _0489_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[105];
  assign _0491_ = _0490_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[104];
  assign _0492_ = _0491_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[103];
  assign _0493_ = _0492_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[102];
  assign _0494_ = _0493_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[101];
  assign _0495_ = _0494_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[100];
  assign _0496_ = _0495_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[99];
  assign _0497_ = _0496_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[98];
  assign _0498_ = _0497_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[97];
  assign _0499_ = _0498_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[96];
  assign _0500_ = _0499_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[95];
  assign _0501_ = _0500_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[94];
  assign _0502_ = _0501_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[93];
  assign _0503_ = _0502_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[92];
  assign _0504_ = _0503_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[91];
  assign _0505_ = _0504_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[90];
  assign _0506_ = _0505_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[89];
  assign _0507_ = _0506_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[88];
  assign _0508_ = _0507_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[87];
  assign _0509_ = _0508_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[86];
  assign _0510_ = _0509_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[85];
  assign _0511_ = _0510_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[84];
  assign _0512_ = _0511_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[83];
  assign _0513_ = _0512_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[82];
  assign _0514_ = _0513_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[81];
  assign _0515_ = _0514_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[80];
  assign _0516_ = _0515_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[79];
  assign _0517_ = _0516_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[78];
  assign _0518_ = _0517_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[77];
  assign _0519_ = _0518_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[76];
  assign _0520_ = _0519_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[75];
  assign _0521_ = _0520_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[74];
  assign _0522_ = _0521_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[73];
  assign _0523_ = _0522_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[72];
  assign _0524_ = _0523_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[71];
  assign _0525_ = _0524_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[70];
  assign _0526_ = _0525_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[69];
  assign _0527_ = _0526_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[68];
  assign _0528_ = _0527_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[67];
  assign _0529_ = _0528_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[66];
  assign _0530_ = _0529_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[65];
  assign _0531_ = _0530_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[64];
  assign _0532_ = _0531_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[63];
  assign _0533_ = _0532_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[62];
  assign _0534_ = _0533_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[61];
  assign _0535_ = _0534_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[60];
  assign _0536_ = _0535_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[59];
  assign _0537_ = _0536_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[58];
  assign _0538_ = _0537_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[57];
  assign _0539_ = _0538_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[56];
  assign _0540_ = _0539_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[55];
  assign _0541_ = _0540_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[54];
  assign _0542_ = _0541_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[53];
  assign _0543_ = _0542_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[52];
  assign _0544_ = _0543_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[51];
  assign _0545_ = _0544_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[50];
  assign _0546_ = _0545_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[49];
  assign _0547_ = _0546_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[48];
  assign _0548_ = _0547_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[47];
  assign _0549_ = _0548_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[46];
  assign _0550_ = _0549_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[45];
  assign _0551_ = _0550_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[44];
  assign _0552_ = _0551_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[43];
  assign _0553_ = _0552_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[42];
  assign _0554_ = _0553_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[41];
  assign _0555_ = _0554_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[40];
  assign _0556_ = _0555_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[39];
  assign _0557_ = _0556_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[38];
  assign _0558_ = _0557_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[37];
  assign _0559_ = _0558_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[36];
  assign _0560_ = _0559_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[35];
  assign _0561_ = _0560_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[34];
  assign _0562_ = _0561_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[33];
  assign _0563_ = _0562_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[32];
  assign _0564_ = _0563_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[31];
  assign _0565_ = _0564_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[30];
  assign _0566_ = _0565_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[29];
  assign _0567_ = _0566_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[28];
  assign _0568_ = _0567_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[27];
  assign _0569_ = _0568_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[26];
  assign _0570_ = _0569_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[25];
  assign _0571_ = _0570_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[24];
  assign _0572_ = _0571_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[23];
  assign _0573_ = _0572_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[22];
  assign _0574_ = _0573_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[21];
  assign _0575_ = _0574_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[20];
  assign _0576_ = _0575_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[19];
  assign _0577_ = _0576_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[18];
  assign _0578_ = _0577_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[17];
  assign _0579_ = _0578_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[16];
  assign _0580_ = _0579_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[15];
  assign _0581_ = _0580_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[14];
  assign _0582_ = _0581_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[13];
  assign _0583_ = _0582_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[12];
  assign _0584_ = _0583_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[11];
  assign _0585_ = _0584_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[10];
  assign _0586_ = _0585_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[9];
  assign _0587_ = _0586_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[8];
  assign _0588_ = _0587_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[7];
  assign _0589_ = _0588_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[6];
  assign _0590_ = _0589_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[5];
  assign _0591_ = _0590_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[4];
  assign _0592_ = _0591_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[3];
  assign _0593_ = _0592_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[2];
  assign _0594_ = _0593_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[1];
  assign sat_sum = _0594_ + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13408" *) dlv_sat_bit_d1[0];
  assign { sat_carry, sat_count_inc } = sat_count + (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13415" *) sat_sum;
  assign _0595_ = calc_wr_en_d3 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10902" *) cfg_is_int[8:1];
  assign _0596_ = calc_wr_en_d4 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10903" *) cfg_is_fp[8:1];
  assign _0597_ = calc_addr_d3 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10904" *) cfg_is_int[13:9];
  assign _0598_ = calc_addr_d4 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10905" *) cfg_is_fp[13:9];
  assign _0599_ = calc_dlv_valid_d3 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11666" *) cfg_is_int[14];
  assign _0600_ = calc_dlv_valid_d5 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11667" *) cfg_is_fp[14];
  assign _0601_ = calc_dlv_en_d3 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11668" *) cfg_is_int[22:15];
  assign _0602_ = calc_dlv_en_d5 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11669" *) cfg_is_fp[22:15];
  assign _0603_ = calc_stripe_end_d3 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11670" *) cfg_is_int[23];
  assign _0604_ = calc_stripe_end_d5 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11671" *) cfg_is_fp[23];
  assign _0605_ = calc_layer_end_d3 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11672" *) cfg_is_int[24];
  assign _0606_ = calc_layer_end_d5 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11673" *) cfg_is_fp[24];
  assign _0607_ = { calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0], calc_pout_int_vld[0] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11741" *) calc_pout_int_0_sum;
  assign _0608_ = { calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0], calc_pout_fp_vld[0] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11742" *) calc_pout_fp_0_sum;
  assign _0609_ = { calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1], calc_pout_int_vld[1] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11743" *) calc_pout_int_1_sum;
  assign _0610_ = { calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1], calc_pout_fp_vld[1] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11744" *) calc_pout_fp_1_sum;
  assign _0611_ = { calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2], calc_pout_int_vld[2] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11745" *) calc_pout_int_2_sum;
  assign _0612_ = { calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2], calc_pout_fp_vld[2] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11746" *) calc_pout_fp_2_sum;
  assign _0613_ = { calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3], calc_pout_int_vld[3] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11747" *) calc_pout_int_3_sum;
  assign _0614_ = { calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3], calc_pout_fp_vld[3] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11748" *) calc_pout_fp_3_sum;
  assign _0615_ = { calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4], calc_pout_int_vld[4] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11749" *) calc_pout_int_4_sum;
  assign _0616_ = { calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4], calc_pout_fp_vld[4] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11750" *) calc_pout_fp_4_sum;
  assign _0617_ = { calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5], calc_pout_int_vld[5] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11751" *) calc_pout_int_5_sum;
  assign _0618_ = { calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5], calc_pout_fp_vld[5] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11752" *) calc_pout_fp_5_sum;
  assign _0619_ = { calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6], calc_pout_int_vld[6] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11753" *) calc_pout_int_6_sum;
  assign _0620_ = { calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6], calc_pout_fp_vld[6] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11754" *) calc_pout_fp_6_sum;
  assign _0621_ = { calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7], calc_pout_int_vld[7] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11755" *) calc_pout_int_7_sum;
  assign _0622_ = { calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7], calc_pout_fp_vld[7] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11756" *) calc_pout_fp_7_sum;
  assign _0623_ = { calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8], calc_pout_int_vld[8] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11757" *) calc_pout_int_8_sum;
  assign _0624_ = { calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8], calc_pout_fp_vld[8] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11758" *) calc_pout_fp_8_sum;
  assign _0625_ = { calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9], calc_pout_int_vld[9] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11759" *) calc_pout_int_9_sum;
  assign _0626_ = { calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9], calc_pout_fp_vld[9] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11760" *) calc_pout_fp_9_sum;
  assign _0627_ = { calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10], calc_pout_int_vld[10] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11761" *) calc_pout_int_10_sum;
  assign _0628_ = { calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10], calc_pout_fp_vld[10] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11762" *) calc_pout_fp_10_sum;
  assign _0629_ = { calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11], calc_pout_int_vld[11] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11763" *) calc_pout_int_11_sum;
  assign _0630_ = { calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11], calc_pout_fp_vld[11] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11764" *) calc_pout_fp_11_sum;
  assign _0631_ = { calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12], calc_pout_int_vld[12] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11765" *) calc_pout_int_12_sum;
  assign _0632_ = { calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12], calc_pout_fp_vld[12] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11766" *) calc_pout_fp_12_sum;
  assign _0633_ = { calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13], calc_pout_int_vld[13] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11767" *) calc_pout_int_13_sum;
  assign _0634_ = { calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13], calc_pout_fp_vld[13] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11768" *) calc_pout_fp_13_sum;
  assign _0635_ = { calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14], calc_pout_int_vld[14] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11769" *) calc_pout_int_14_sum;
  assign _0636_ = { calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14], calc_pout_fp_vld[14] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11770" *) calc_pout_fp_14_sum;
  assign _0637_ = { calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15], calc_pout_int_vld[15] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11771" *) calc_pout_int_15_sum;
  assign _0638_ = { calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15], calc_pout_fp_vld[15] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11772" *) calc_pout_fp_15_sum;
  assign _0639_ = { calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16], calc_pout_int_vld[16] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11773" *) calc_pout_int_16_sum;
  assign _0640_ = { calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16], calc_pout_fp_vld[16] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11774" *) calc_pout_fp_16_sum;
  assign _0641_ = { calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17], calc_pout_int_vld[17] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11775" *) calc_pout_int_17_sum;
  assign _0642_ = { calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17], calc_pout_fp_vld[17] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11776" *) calc_pout_fp_17_sum;
  assign _0643_ = { calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18], calc_pout_int_vld[18] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11777" *) calc_pout_int_18_sum;
  assign _0644_ = { calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18], calc_pout_fp_vld[18] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11778" *) calc_pout_fp_18_sum;
  assign _0645_ = { calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19], calc_pout_int_vld[19] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11779" *) calc_pout_int_19_sum;
  assign _0646_ = { calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19], calc_pout_fp_vld[19] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11780" *) calc_pout_fp_19_sum;
  assign _0647_ = { calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20], calc_pout_int_vld[20] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11781" *) calc_pout_int_20_sum;
  assign _0648_ = { calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20], calc_pout_fp_vld[20] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11782" *) calc_pout_fp_20_sum;
  assign _0649_ = { calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21], calc_pout_int_vld[21] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11783" *) calc_pout_int_21_sum;
  assign _0650_ = { calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21], calc_pout_fp_vld[21] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11784" *) calc_pout_fp_21_sum;
  assign _0651_ = { calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22], calc_pout_int_vld[22] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11785" *) calc_pout_int_22_sum;
  assign _0652_ = { calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22], calc_pout_fp_vld[22] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11786" *) calc_pout_fp_22_sum;
  assign _0653_ = { calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23], calc_pout_int_vld[23] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11787" *) calc_pout_int_23_sum;
  assign _0654_ = { calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23], calc_pout_fp_vld[23] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11788" *) calc_pout_fp_23_sum;
  assign _0655_ = { calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24], calc_pout_int_vld[24] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11789" *) calc_pout_int_24_sum;
  assign _0656_ = { calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24], calc_pout_fp_vld[24] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11790" *) calc_pout_fp_24_sum;
  assign _0657_ = { calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25], calc_pout_int_vld[25] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11791" *) calc_pout_int_25_sum;
  assign _0658_ = { calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25], calc_pout_fp_vld[25] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11792" *) calc_pout_fp_25_sum;
  assign _0659_ = { calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26], calc_pout_int_vld[26] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11793" *) calc_pout_int_26_sum;
  assign _0660_ = { calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26], calc_pout_fp_vld[26] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11794" *) calc_pout_fp_26_sum;
  assign _0661_ = { calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27], calc_pout_int_vld[27] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11795" *) calc_pout_int_27_sum;
  assign _0662_ = { calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27], calc_pout_fp_vld[27] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11796" *) calc_pout_fp_27_sum;
  assign _0663_ = { calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28], calc_pout_int_vld[28] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11797" *) calc_pout_int_28_sum;
  assign _0664_ = { calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28], calc_pout_fp_vld[28] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11798" *) calc_pout_fp_28_sum;
  assign _0665_ = { calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29], calc_pout_int_vld[29] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11799" *) calc_pout_int_29_sum;
  assign _0666_ = { calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29], calc_pout_fp_vld[29] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11800" *) calc_pout_fp_29_sum;
  assign _0667_ = { calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30], calc_pout_int_vld[30] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11801" *) calc_pout_int_30_sum;
  assign _0668_ = { calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30], calc_pout_fp_vld[30] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11802" *) calc_pout_fp_30_sum;
  assign _0669_ = { calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31], calc_pout_int_vld[31] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11803" *) calc_pout_int_31_sum;
  assign _0670_ = { calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31], calc_pout_fp_vld[31] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11804" *) calc_pout_fp_31_sum;
  assign _0671_ = { calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32], calc_pout_int_vld[32] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11805" *) calc_pout_int_32_sum;
  assign _0672_ = { calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32], calc_pout_fp_vld[32] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11806" *) calc_pout_fp_32_sum;
  assign _0673_ = { calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33], calc_pout_int_vld[33] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11807" *) calc_pout_int_33_sum;
  assign _0674_ = { calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33], calc_pout_fp_vld[33] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11808" *) calc_pout_fp_33_sum;
  assign _0675_ = { calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34], calc_pout_int_vld[34] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11809" *) calc_pout_int_34_sum;
  assign _0676_ = { calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34], calc_pout_fp_vld[34] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11810" *) calc_pout_fp_34_sum;
  assign _0677_ = { calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35], calc_pout_int_vld[35] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11811" *) calc_pout_int_35_sum;
  assign _0678_ = { calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35], calc_pout_fp_vld[35] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11812" *) calc_pout_fp_35_sum;
  assign _0679_ = { calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36], calc_pout_int_vld[36] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11813" *) calc_pout_int_36_sum;
  assign _0680_ = { calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36], calc_pout_fp_vld[36] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11814" *) calc_pout_fp_36_sum;
  assign _0681_ = { calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37], calc_pout_int_vld[37] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11815" *) calc_pout_int_37_sum;
  assign _0682_ = { calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37], calc_pout_fp_vld[37] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11816" *) calc_pout_fp_37_sum;
  assign _0683_ = { calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38], calc_pout_int_vld[38] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11817" *) calc_pout_int_38_sum;
  assign _0684_ = { calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38], calc_pout_fp_vld[38] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11818" *) calc_pout_fp_38_sum;
  assign _0685_ = { calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39], calc_pout_int_vld[39] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11819" *) calc_pout_int_39_sum;
  assign _0686_ = { calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39], calc_pout_fp_vld[39] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11820" *) calc_pout_fp_39_sum;
  assign _0687_ = { calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40], calc_pout_int_vld[40] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11821" *) calc_pout_int_40_sum;
  assign _0688_ = { calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40], calc_pout_fp_vld[40] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11822" *) calc_pout_fp_40_sum;
  assign _0689_ = { calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41], calc_pout_int_vld[41] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11823" *) calc_pout_int_41_sum;
  assign _0690_ = { calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41], calc_pout_fp_vld[41] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11824" *) calc_pout_fp_41_sum;
  assign _0691_ = { calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42], calc_pout_int_vld[42] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11825" *) calc_pout_int_42_sum;
  assign _0692_ = { calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42], calc_pout_fp_vld[42] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11826" *) calc_pout_fp_42_sum;
  assign _0693_ = { calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43], calc_pout_int_vld[43] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11827" *) calc_pout_int_43_sum;
  assign _0694_ = { calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43], calc_pout_fp_vld[43] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11828" *) calc_pout_fp_43_sum;
  assign _0695_ = { calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44], calc_pout_int_vld[44] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11829" *) calc_pout_int_44_sum;
  assign _0696_ = { calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44], calc_pout_fp_vld[44] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11830" *) calc_pout_fp_44_sum;
  assign _0697_ = { calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45], calc_pout_int_vld[45] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11831" *) calc_pout_int_45_sum;
  assign _0698_ = { calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45], calc_pout_fp_vld[45] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11832" *) calc_pout_fp_45_sum;
  assign _0699_ = { calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46], calc_pout_int_vld[46] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11833" *) calc_pout_int_46_sum;
  assign _0700_ = { calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46], calc_pout_fp_vld[46] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11834" *) calc_pout_fp_46_sum;
  assign _0701_ = { calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47], calc_pout_int_vld[47] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11835" *) calc_pout_int_47_sum;
  assign _0702_ = { calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47], calc_pout_fp_vld[47] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11836" *) calc_pout_fp_47_sum;
  assign _0703_ = { calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48], calc_pout_int_vld[48] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11837" *) calc_pout_int_48_sum;
  assign _0704_ = { calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48], calc_pout_fp_vld[48] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11838" *) calc_pout_fp_48_sum;
  assign _0705_ = { calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49], calc_pout_int_vld[49] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11839" *) calc_pout_int_49_sum;
  assign _0706_ = { calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49], calc_pout_fp_vld[49] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11840" *) calc_pout_fp_49_sum;
  assign _0707_ = { calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50], calc_pout_int_vld[50] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11841" *) calc_pout_int_50_sum;
  assign _0708_ = { calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50], calc_pout_fp_vld[50] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11842" *) calc_pout_fp_50_sum;
  assign _0709_ = { calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51], calc_pout_int_vld[51] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11843" *) calc_pout_int_51_sum;
  assign _0710_ = { calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51], calc_pout_fp_vld[51] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11844" *) calc_pout_fp_51_sum;
  assign _0711_ = { calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52], calc_pout_int_vld[52] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11845" *) calc_pout_int_52_sum;
  assign _0712_ = { calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52], calc_pout_fp_vld[52] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11846" *) calc_pout_fp_52_sum;
  assign _0713_ = { calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53], calc_pout_int_vld[53] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11847" *) calc_pout_int_53_sum;
  assign _0714_ = { calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53], calc_pout_fp_vld[53] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11848" *) calc_pout_fp_53_sum;
  assign _0715_ = { calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54], calc_pout_int_vld[54] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11849" *) calc_pout_int_54_sum;
  assign _0716_ = { calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54], calc_pout_fp_vld[54] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11850" *) calc_pout_fp_54_sum;
  assign _0717_ = { calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55], calc_pout_int_vld[55] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11851" *) calc_pout_int_55_sum;
  assign _0718_ = { calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55], calc_pout_fp_vld[55] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11852" *) calc_pout_fp_55_sum;
  assign _0719_ = { calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56], calc_pout_int_vld[56] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11853" *) calc_pout_int_56_sum;
  assign _0720_ = { calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56], calc_pout_fp_vld[56] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11854" *) calc_pout_fp_56_sum;
  assign _0721_ = { calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57], calc_pout_int_vld[57] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11855" *) calc_pout_int_57_sum;
  assign _0722_ = { calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57], calc_pout_fp_vld[57] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11856" *) calc_pout_fp_57_sum;
  assign _0723_ = { calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58], calc_pout_int_vld[58] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11857" *) calc_pout_int_58_sum;
  assign _0724_ = { calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58], calc_pout_fp_vld[58] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11858" *) calc_pout_fp_58_sum;
  assign _0725_ = { calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59], calc_pout_int_vld[59] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11859" *) calc_pout_int_59_sum;
  assign _0726_ = { calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59], calc_pout_fp_vld[59] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11860" *) calc_pout_fp_59_sum;
  assign _0727_ = { calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60], calc_pout_int_vld[60] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11861" *) calc_pout_int_60_sum;
  assign _0728_ = { calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60], calc_pout_fp_vld[60] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11862" *) calc_pout_fp_60_sum;
  assign _0729_ = { calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61], calc_pout_int_vld[61] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11863" *) calc_pout_int_61_sum;
  assign _0730_ = { calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61], calc_pout_fp_vld[61] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11864" *) calc_pout_fp_61_sum;
  assign _0731_ = { calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62], calc_pout_int_vld[62] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11865" *) calc_pout_int_62_sum;
  assign _0732_ = { calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62], calc_pout_fp_vld[62] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11866" *) calc_pout_fp_62_sum;
  assign _0733_ = { calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63], calc_pout_int_vld[63] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11867" *) calc_pout_int_63_sum;
  assign _0734_ = { calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63], calc_pout_fp_vld[63] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11868" *) calc_pout_fp_63_sum;
  assign calc_pout_64 = { calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64], calc_pout_int_vld[64] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11869" *) calc_pout_int_64_sum;
  assign calc_pout_65 = { calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65], calc_pout_int_vld[65] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11870" *) calc_pout_int_65_sum;
  assign calc_pout_66 = { calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66], calc_pout_int_vld[66] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11871" *) calc_pout_int_66_sum;
  assign calc_pout_67 = { calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67], calc_pout_int_vld[67] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11872" *) calc_pout_int_67_sum;
  assign calc_pout_68 = { calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68], calc_pout_int_vld[68] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11873" *) calc_pout_int_68_sum;
  assign calc_pout_69 = { calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69], calc_pout_int_vld[69] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11874" *) calc_pout_int_69_sum;
  assign calc_pout_70 = { calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70], calc_pout_int_vld[70] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11875" *) calc_pout_int_70_sum;
  assign calc_pout_71 = { calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71], calc_pout_int_vld[71] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11876" *) calc_pout_int_71_sum;
  assign calc_pout_72 = { calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72], calc_pout_int_vld[72] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11877" *) calc_pout_int_72_sum;
  assign calc_pout_73 = { calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73], calc_pout_int_vld[73] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11878" *) calc_pout_int_73_sum;
  assign calc_pout_74 = { calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74], calc_pout_int_vld[74] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11879" *) calc_pout_int_74_sum;
  assign calc_pout_75 = { calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75], calc_pout_int_vld[75] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11880" *) calc_pout_int_75_sum;
  assign calc_pout_76 = { calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76], calc_pout_int_vld[76] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11881" *) calc_pout_int_76_sum;
  assign calc_pout_77 = { calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77], calc_pout_int_vld[77] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11882" *) calc_pout_int_77_sum;
  assign calc_pout_78 = { calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78], calc_pout_int_vld[78] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11883" *) calc_pout_int_78_sum;
  assign calc_pout_79 = { calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79], calc_pout_int_vld[79] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11884" *) calc_pout_int_79_sum;
  assign calc_pout_80 = { calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80], calc_pout_int_vld[80] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11885" *) calc_pout_int_80_sum;
  assign calc_pout_81 = { calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81], calc_pout_int_vld[81] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11886" *) calc_pout_int_81_sum;
  assign calc_pout_82 = { calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82], calc_pout_int_vld[82] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11887" *) calc_pout_int_82_sum;
  assign calc_pout_83 = { calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83], calc_pout_int_vld[83] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11888" *) calc_pout_int_83_sum;
  assign calc_pout_84 = { calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84], calc_pout_int_vld[84] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11889" *) calc_pout_int_84_sum;
  assign calc_pout_85 = { calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85], calc_pout_int_vld[85] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11890" *) calc_pout_int_85_sum;
  assign calc_pout_86 = { calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86], calc_pout_int_vld[86] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11891" *) calc_pout_int_86_sum;
  assign calc_pout_87 = { calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87], calc_pout_int_vld[87] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11892" *) calc_pout_int_87_sum;
  assign calc_pout_88 = { calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88], calc_pout_int_vld[88] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11893" *) calc_pout_int_88_sum;
  assign calc_pout_89 = { calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89], calc_pout_int_vld[89] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11894" *) calc_pout_int_89_sum;
  assign calc_pout_90 = { calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90], calc_pout_int_vld[90] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11895" *) calc_pout_int_90_sum;
  assign calc_pout_91 = { calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91], calc_pout_int_vld[91] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11896" *) calc_pout_int_91_sum;
  assign calc_pout_92 = { calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92], calc_pout_int_vld[92] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11897" *) calc_pout_int_92_sum;
  assign calc_pout_93 = { calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93], calc_pout_int_vld[93] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11898" *) calc_pout_int_93_sum;
  assign calc_pout_94 = { calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94], calc_pout_int_vld[94] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11899" *) calc_pout_int_94_sum;
  assign calc_pout_95 = { calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95], calc_pout_int_vld[95] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11900" *) calc_pout_int_95_sum;
  assign calc_pout_96 = { calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96], calc_pout_int_vld[96] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11901" *) calc_pout_int_96_sum;
  assign calc_pout_97 = { calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97], calc_pout_int_vld[97] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11902" *) calc_pout_int_97_sum;
  assign calc_pout_98 = { calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98], calc_pout_int_vld[98] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11903" *) calc_pout_int_98_sum;
  assign calc_pout_99 = { calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99], calc_pout_int_vld[99] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11904" *) calc_pout_int_99_sum;
  assign calc_pout_100 = { calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100], calc_pout_int_vld[100] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11905" *) calc_pout_int_100_sum;
  assign calc_pout_101 = { calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101], calc_pout_int_vld[101] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11906" *) calc_pout_int_101_sum;
  assign calc_pout_102 = { calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102], calc_pout_int_vld[102] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11907" *) calc_pout_int_102_sum;
  assign calc_pout_103 = { calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103], calc_pout_int_vld[103] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11908" *) calc_pout_int_103_sum;
  assign calc_pout_104 = { calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104], calc_pout_int_vld[104] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11909" *) calc_pout_int_104_sum;
  assign calc_pout_105 = { calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105], calc_pout_int_vld[105] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11910" *) calc_pout_int_105_sum;
  assign calc_pout_106 = { calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106], calc_pout_int_vld[106] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11911" *) calc_pout_int_106_sum;
  assign calc_pout_107 = { calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107], calc_pout_int_vld[107] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11912" *) calc_pout_int_107_sum;
  assign calc_pout_108 = { calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108], calc_pout_int_vld[108] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11913" *) calc_pout_int_108_sum;
  assign calc_pout_109 = { calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109], calc_pout_int_vld[109] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11914" *) calc_pout_int_109_sum;
  assign calc_pout_110 = { calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110], calc_pout_int_vld[110] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11915" *) calc_pout_int_110_sum;
  assign calc_pout_111 = { calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111], calc_pout_int_vld[111] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11916" *) calc_pout_int_111_sum;
  assign calc_pout_112 = { calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112], calc_pout_int_vld[112] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11917" *) calc_pout_int_112_sum;
  assign calc_pout_113 = { calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113], calc_pout_int_vld[113] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11918" *) calc_pout_int_113_sum;
  assign calc_pout_114 = { calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114], calc_pout_int_vld[114] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11919" *) calc_pout_int_114_sum;
  assign calc_pout_115 = { calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115], calc_pout_int_vld[115] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11920" *) calc_pout_int_115_sum;
  assign calc_pout_116 = { calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116], calc_pout_int_vld[116] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11921" *) calc_pout_int_116_sum;
  assign calc_pout_117 = { calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117], calc_pout_int_vld[117] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11922" *) calc_pout_int_117_sum;
  assign calc_pout_118 = { calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118], calc_pout_int_vld[118] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11923" *) calc_pout_int_118_sum;
  assign calc_pout_119 = { calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119], calc_pout_int_vld[119] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11924" *) calc_pout_int_119_sum;
  assign calc_pout_120 = { calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120], calc_pout_int_vld[120] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11925" *) calc_pout_int_120_sum;
  assign calc_pout_121 = { calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121], calc_pout_int_vld[121] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11926" *) calc_pout_int_121_sum;
  assign calc_pout_122 = { calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122], calc_pout_int_vld[122] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11927" *) calc_pout_int_122_sum;
  assign calc_pout_123 = { calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123], calc_pout_int_vld[123] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11928" *) calc_pout_int_123_sum;
  assign calc_pout_124 = { calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124], calc_pout_int_vld[124] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11929" *) calc_pout_int_124_sum;
  assign calc_pout_125 = { calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125], calc_pout_int_vld[125] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11930" *) calc_pout_int_125_sum;
  assign calc_pout_126 = { calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126], calc_pout_int_vld[126] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11931" *) calc_pout_int_126_sum;
  assign calc_pout_127 = { calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127], calc_pout_int_vld[127] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11932" *) calc_pout_int_127_sum;
  assign _0735_ = { calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0], calc_fout_int_vld[0] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11933" *) calc_fout_int_0_sum;
  assign _0736_ = { calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0], calc_fout_fp_vld[0] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11934" *) calc_fout_fp_0_sum;
  assign _0737_ = { calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1], calc_fout_int_vld[1] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11935" *) calc_fout_int_1_sum;
  assign _0738_ = { calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1], calc_fout_fp_vld[1] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11936" *) calc_fout_fp_1_sum;
  assign _0739_ = { calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2], calc_fout_int_vld[2] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11937" *) calc_fout_int_2_sum;
  assign _0740_ = { calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2], calc_fout_fp_vld[2] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11938" *) calc_fout_fp_2_sum;
  assign _0741_ = { calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3], calc_fout_int_vld[3] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11939" *) calc_fout_int_3_sum;
  assign _0742_ = { calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3], calc_fout_fp_vld[3] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11940" *) calc_fout_fp_3_sum;
  assign _0743_ = { calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4], calc_fout_int_vld[4] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11941" *) calc_fout_int_4_sum;
  assign _0744_ = { calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4], calc_fout_fp_vld[4] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11942" *) calc_fout_fp_4_sum;
  assign _0745_ = { calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5], calc_fout_int_vld[5] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11943" *) calc_fout_int_5_sum;
  assign _0746_ = { calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5], calc_fout_fp_vld[5] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11944" *) calc_fout_fp_5_sum;
  assign _0747_ = { calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6], calc_fout_int_vld[6] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11945" *) calc_fout_int_6_sum;
  assign _0748_ = { calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6], calc_fout_fp_vld[6] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11946" *) calc_fout_fp_6_sum;
  assign _0749_ = { calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7], calc_fout_int_vld[7] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11947" *) calc_fout_int_7_sum;
  assign _0750_ = { calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7], calc_fout_fp_vld[7] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11948" *) calc_fout_fp_7_sum;
  assign _0751_ = { calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8], calc_fout_int_vld[8] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11949" *) calc_fout_int_8_sum;
  assign _0752_ = { calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8], calc_fout_fp_vld[8] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11950" *) calc_fout_fp_8_sum;
  assign _0753_ = { calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9], calc_fout_int_vld[9] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11951" *) calc_fout_int_9_sum;
  assign _0754_ = { calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9], calc_fout_fp_vld[9] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11952" *) calc_fout_fp_9_sum;
  assign _0755_ = { calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10], calc_fout_int_vld[10] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11953" *) calc_fout_int_10_sum;
  assign _0756_ = { calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10], calc_fout_fp_vld[10] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11954" *) calc_fout_fp_10_sum;
  assign _0757_ = { calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11], calc_fout_int_vld[11] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11955" *) calc_fout_int_11_sum;
  assign _0758_ = { calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11], calc_fout_fp_vld[11] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11956" *) calc_fout_fp_11_sum;
  assign _0759_ = { calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12], calc_fout_int_vld[12] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11957" *) calc_fout_int_12_sum;
  assign _0760_ = { calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12], calc_fout_fp_vld[12] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11958" *) calc_fout_fp_12_sum;
  assign _0761_ = { calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13], calc_fout_int_vld[13] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11959" *) calc_fout_int_13_sum;
  assign _0762_ = { calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13], calc_fout_fp_vld[13] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11960" *) calc_fout_fp_13_sum;
  assign _0763_ = { calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14], calc_fout_int_vld[14] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11961" *) calc_fout_int_14_sum;
  assign _0764_ = { calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14], calc_fout_fp_vld[14] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11962" *) calc_fout_fp_14_sum;
  assign _0765_ = { calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15], calc_fout_int_vld[15] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11963" *) calc_fout_int_15_sum;
  assign _0766_ = { calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15], calc_fout_fp_vld[15] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11964" *) calc_fout_fp_15_sum;
  assign _0767_ = { calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16], calc_fout_int_vld[16] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11965" *) calc_fout_int_16_sum;
  assign _0768_ = { calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16], calc_fout_fp_vld[16] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11966" *) calc_fout_fp_16_sum;
  assign _0769_ = { calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17], calc_fout_int_vld[17] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11967" *) calc_fout_int_17_sum;
  assign _0770_ = { calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17], calc_fout_fp_vld[17] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11968" *) calc_fout_fp_17_sum;
  assign _0771_ = { calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18], calc_fout_int_vld[18] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11969" *) calc_fout_int_18_sum;
  assign _0772_ = { calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18], calc_fout_fp_vld[18] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11970" *) calc_fout_fp_18_sum;
  assign _0773_ = { calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19], calc_fout_int_vld[19] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11971" *) calc_fout_int_19_sum;
  assign _0774_ = { calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19], calc_fout_fp_vld[19] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11972" *) calc_fout_fp_19_sum;
  assign _0775_ = { calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20], calc_fout_int_vld[20] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11973" *) calc_fout_int_20_sum;
  assign _0776_ = { calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20], calc_fout_fp_vld[20] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11974" *) calc_fout_fp_20_sum;
  assign _0777_ = { calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21], calc_fout_int_vld[21] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11975" *) calc_fout_int_21_sum;
  assign _0778_ = { calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21], calc_fout_fp_vld[21] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11976" *) calc_fout_fp_21_sum;
  assign _0779_ = { calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22], calc_fout_int_vld[22] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11977" *) calc_fout_int_22_sum;
  assign _0780_ = { calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22], calc_fout_fp_vld[22] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11978" *) calc_fout_fp_22_sum;
  assign _0781_ = { calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23], calc_fout_int_vld[23] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11979" *) calc_fout_int_23_sum;
  assign _0782_ = { calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23], calc_fout_fp_vld[23] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11980" *) calc_fout_fp_23_sum;
  assign _0783_ = { calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24], calc_fout_int_vld[24] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11981" *) calc_fout_int_24_sum;
  assign _0784_ = { calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24], calc_fout_fp_vld[24] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11982" *) calc_fout_fp_24_sum;
  assign _0785_ = { calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25], calc_fout_int_vld[25] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11983" *) calc_fout_int_25_sum;
  assign _0786_ = { calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25], calc_fout_fp_vld[25] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11984" *) calc_fout_fp_25_sum;
  assign _0787_ = { calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26], calc_fout_int_vld[26] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11985" *) calc_fout_int_26_sum;
  assign _0788_ = { calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26], calc_fout_fp_vld[26] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11986" *) calc_fout_fp_26_sum;
  assign _0789_ = { calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27], calc_fout_int_vld[27] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11987" *) calc_fout_int_27_sum;
  assign _0790_ = { calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27], calc_fout_fp_vld[27] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11988" *) calc_fout_fp_27_sum;
  assign _0791_ = { calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28], calc_fout_int_vld[28] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11989" *) calc_fout_int_28_sum;
  assign _0792_ = { calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28], calc_fout_fp_vld[28] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11990" *) calc_fout_fp_28_sum;
  assign _0793_ = { calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29], calc_fout_int_vld[29] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11991" *) calc_fout_int_29_sum;
  assign _0794_ = { calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29], calc_fout_fp_vld[29] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11992" *) calc_fout_fp_29_sum;
  assign _0795_ = { calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30], calc_fout_int_vld[30] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11993" *) calc_fout_int_30_sum;
  assign _0796_ = { calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30], calc_fout_fp_vld[30] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11994" *) calc_fout_fp_30_sum;
  assign _0797_ = { calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31], calc_fout_int_vld[31] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11995" *) calc_fout_int_31_sum;
  assign _0798_ = { calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31], calc_fout_fp_vld[31] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11996" *) calc_fout_fp_31_sum;
  assign _0799_ = { calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32], calc_fout_int_vld[32] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11997" *) calc_fout_int_32_sum;
  assign _0800_ = { calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32], calc_fout_fp_vld[32] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11998" *) calc_fout_fp_32_sum;
  assign _0801_ = { calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33], calc_fout_int_vld[33] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11999" *) calc_fout_int_33_sum;
  assign _0802_ = { calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33], calc_fout_fp_vld[33] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12000" *) calc_fout_fp_33_sum;
  assign _0803_ = { calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34], calc_fout_int_vld[34] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12001" *) calc_fout_int_34_sum;
  assign _0804_ = { calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34], calc_fout_fp_vld[34] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12002" *) calc_fout_fp_34_sum;
  assign _0805_ = { calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35], calc_fout_int_vld[35] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12003" *) calc_fout_int_35_sum;
  assign _0806_ = { calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35], calc_fout_fp_vld[35] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12004" *) calc_fout_fp_35_sum;
  assign _0807_ = { calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36], calc_fout_int_vld[36] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12005" *) calc_fout_int_36_sum;
  assign _0808_ = { calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36], calc_fout_fp_vld[36] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12006" *) calc_fout_fp_36_sum;
  assign _0809_ = { calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37], calc_fout_int_vld[37] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12007" *) calc_fout_int_37_sum;
  assign _0810_ = { calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37], calc_fout_fp_vld[37] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12008" *) calc_fout_fp_37_sum;
  assign _0811_ = { calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38], calc_fout_int_vld[38] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12009" *) calc_fout_int_38_sum;
  assign _0812_ = { calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38], calc_fout_fp_vld[38] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12010" *) calc_fout_fp_38_sum;
  assign _0813_ = { calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39], calc_fout_int_vld[39] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12011" *) calc_fout_int_39_sum;
  assign _0814_ = { calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39], calc_fout_fp_vld[39] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12012" *) calc_fout_fp_39_sum;
  assign _0815_ = { calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40], calc_fout_int_vld[40] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12013" *) calc_fout_int_40_sum;
  assign _0816_ = { calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40], calc_fout_fp_vld[40] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12014" *) calc_fout_fp_40_sum;
  assign _0817_ = { calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41], calc_fout_int_vld[41] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12015" *) calc_fout_int_41_sum;
  assign _0818_ = { calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41], calc_fout_fp_vld[41] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12016" *) calc_fout_fp_41_sum;
  assign _0819_ = { calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42], calc_fout_int_vld[42] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12017" *) calc_fout_int_42_sum;
  assign _0820_ = { calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42], calc_fout_fp_vld[42] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12018" *) calc_fout_fp_42_sum;
  assign _0821_ = { calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43], calc_fout_int_vld[43] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12019" *) calc_fout_int_43_sum;
  assign _0822_ = { calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43], calc_fout_fp_vld[43] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12020" *) calc_fout_fp_43_sum;
  assign _0823_ = { calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44], calc_fout_int_vld[44] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12021" *) calc_fout_int_44_sum;
  assign _0824_ = { calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44], calc_fout_fp_vld[44] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12022" *) calc_fout_fp_44_sum;
  assign _0825_ = { calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45], calc_fout_int_vld[45] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12023" *) calc_fout_int_45_sum;
  assign _0826_ = { calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45], calc_fout_fp_vld[45] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12024" *) calc_fout_fp_45_sum;
  assign _0827_ = { calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46], calc_fout_int_vld[46] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12025" *) calc_fout_int_46_sum;
  assign _0828_ = { calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46], calc_fout_fp_vld[46] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12026" *) calc_fout_fp_46_sum;
  assign _0829_ = { calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47], calc_fout_int_vld[47] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12027" *) calc_fout_int_47_sum;
  assign _0830_ = { calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47], calc_fout_fp_vld[47] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12028" *) calc_fout_fp_47_sum;
  assign _0831_ = { calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48], calc_fout_int_vld[48] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12029" *) calc_fout_int_48_sum;
  assign _0832_ = { calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48], calc_fout_fp_vld[48] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12030" *) calc_fout_fp_48_sum;
  assign _0833_ = { calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49], calc_fout_int_vld[49] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12031" *) calc_fout_int_49_sum;
  assign _0834_ = { calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49], calc_fout_fp_vld[49] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12032" *) calc_fout_fp_49_sum;
  assign _0835_ = { calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50], calc_fout_int_vld[50] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12033" *) calc_fout_int_50_sum;
  assign _0836_ = { calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50], calc_fout_fp_vld[50] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12034" *) calc_fout_fp_50_sum;
  assign _0837_ = { calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51], calc_fout_int_vld[51] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12035" *) calc_fout_int_51_sum;
  assign _0838_ = { calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51], calc_fout_fp_vld[51] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12036" *) calc_fout_fp_51_sum;
  assign _0839_ = { calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52], calc_fout_int_vld[52] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12037" *) calc_fout_int_52_sum;
  assign _0840_ = { calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52], calc_fout_fp_vld[52] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12038" *) calc_fout_fp_52_sum;
  assign _0841_ = { calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53], calc_fout_int_vld[53] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12039" *) calc_fout_int_53_sum;
  assign _0842_ = { calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53], calc_fout_fp_vld[53] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12040" *) calc_fout_fp_53_sum;
  assign _0843_ = { calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54], calc_fout_int_vld[54] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12041" *) calc_fout_int_54_sum;
  assign _0844_ = { calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54], calc_fout_fp_vld[54] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12042" *) calc_fout_fp_54_sum;
  assign _0845_ = { calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55], calc_fout_int_vld[55] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12043" *) calc_fout_int_55_sum;
  assign _0846_ = { calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55], calc_fout_fp_vld[55] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12044" *) calc_fout_fp_55_sum;
  assign _0847_ = { calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56], calc_fout_int_vld[56] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12045" *) calc_fout_int_56_sum;
  assign _0848_ = { calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56], calc_fout_fp_vld[56] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12046" *) calc_fout_fp_56_sum;
  assign _0849_ = { calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57], calc_fout_int_vld[57] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12047" *) calc_fout_int_57_sum;
  assign _0850_ = { calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57], calc_fout_fp_vld[57] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12048" *) calc_fout_fp_57_sum;
  assign _0851_ = { calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58], calc_fout_int_vld[58] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12049" *) calc_fout_int_58_sum;
  assign _0852_ = { calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58], calc_fout_fp_vld[58] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12050" *) calc_fout_fp_58_sum;
  assign _0853_ = { calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59], calc_fout_int_vld[59] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12051" *) calc_fout_int_59_sum;
  assign _0854_ = { calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59], calc_fout_fp_vld[59] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12052" *) calc_fout_fp_59_sum;
  assign _0855_ = { calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60], calc_fout_int_vld[60] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12053" *) calc_fout_int_60_sum;
  assign _0856_ = { calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60], calc_fout_fp_vld[60] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12054" *) calc_fout_fp_60_sum;
  assign _0857_ = { calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61], calc_fout_int_vld[61] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12055" *) calc_fout_int_61_sum;
  assign _0858_ = { calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61], calc_fout_fp_vld[61] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12056" *) calc_fout_fp_61_sum;
  assign _0859_ = { calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62], calc_fout_int_vld[62] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12057" *) calc_fout_int_62_sum;
  assign _0860_ = { calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62], calc_fout_fp_vld[62] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12058" *) calc_fout_fp_62_sum;
  assign _0861_ = { calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63], calc_fout_int_vld[63] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12059" *) calc_fout_int_63_sum;
  assign _0862_ = { calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63], calc_fout_fp_vld[63] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12060" *) calc_fout_fp_63_sum;
  assign calc_fout_64 = { calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64], calc_fout_int_vld[64] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12061" *) calc_fout_int_64_sum;
  assign calc_fout_65 = { calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65], calc_fout_int_vld[65] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12062" *) calc_fout_int_65_sum;
  assign calc_fout_66 = { calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66], calc_fout_int_vld[66] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12063" *) calc_fout_int_66_sum;
  assign calc_fout_67 = { calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67], calc_fout_int_vld[67] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12064" *) calc_fout_int_67_sum;
  assign calc_fout_68 = { calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68], calc_fout_int_vld[68] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12065" *) calc_fout_int_68_sum;
  assign calc_fout_69 = { calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69], calc_fout_int_vld[69] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12066" *) calc_fout_int_69_sum;
  assign calc_fout_70 = { calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70], calc_fout_int_vld[70] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12067" *) calc_fout_int_70_sum;
  assign calc_fout_71 = { calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71], calc_fout_int_vld[71] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12068" *) calc_fout_int_71_sum;
  assign calc_fout_72 = { calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72], calc_fout_int_vld[72] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12069" *) calc_fout_int_72_sum;
  assign calc_fout_73 = { calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73], calc_fout_int_vld[73] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12070" *) calc_fout_int_73_sum;
  assign calc_fout_74 = { calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74], calc_fout_int_vld[74] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12071" *) calc_fout_int_74_sum;
  assign calc_fout_75 = { calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75], calc_fout_int_vld[75] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12072" *) calc_fout_int_75_sum;
  assign calc_fout_76 = { calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76], calc_fout_int_vld[76] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12073" *) calc_fout_int_76_sum;
  assign calc_fout_77 = { calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77], calc_fout_int_vld[77] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12074" *) calc_fout_int_77_sum;
  assign calc_fout_78 = { calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78], calc_fout_int_vld[78] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12075" *) calc_fout_int_78_sum;
  assign calc_fout_79 = { calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79], calc_fout_int_vld[79] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12076" *) calc_fout_int_79_sum;
  assign calc_fout_80 = { calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80], calc_fout_int_vld[80] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12077" *) calc_fout_int_80_sum;
  assign calc_fout_81 = { calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81], calc_fout_int_vld[81] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12078" *) calc_fout_int_81_sum;
  assign calc_fout_82 = { calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82], calc_fout_int_vld[82] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12079" *) calc_fout_int_82_sum;
  assign calc_fout_83 = { calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83], calc_fout_int_vld[83] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12080" *) calc_fout_int_83_sum;
  assign calc_fout_84 = { calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84], calc_fout_int_vld[84] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12081" *) calc_fout_int_84_sum;
  assign calc_fout_85 = { calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85], calc_fout_int_vld[85] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12082" *) calc_fout_int_85_sum;
  assign calc_fout_86 = { calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86], calc_fout_int_vld[86] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12083" *) calc_fout_int_86_sum;
  assign calc_fout_87 = { calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87], calc_fout_int_vld[87] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12084" *) calc_fout_int_87_sum;
  assign calc_fout_88 = { calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88], calc_fout_int_vld[88] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12085" *) calc_fout_int_88_sum;
  assign calc_fout_89 = { calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89], calc_fout_int_vld[89] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12086" *) calc_fout_int_89_sum;
  assign calc_fout_90 = { calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90], calc_fout_int_vld[90] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12087" *) calc_fout_int_90_sum;
  assign calc_fout_91 = { calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91], calc_fout_int_vld[91] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12088" *) calc_fout_int_91_sum;
  assign calc_fout_92 = { calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92], calc_fout_int_vld[92] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12089" *) calc_fout_int_92_sum;
  assign calc_fout_93 = { calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93], calc_fout_int_vld[93] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12090" *) calc_fout_int_93_sum;
  assign calc_fout_94 = { calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94], calc_fout_int_vld[94] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12091" *) calc_fout_int_94_sum;
  assign calc_fout_95 = { calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95], calc_fout_int_vld[95] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12092" *) calc_fout_int_95_sum;
  assign calc_dlv_elem_65 = { calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96], calc_fout_int_vld[96] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12093" *) calc_fout_int_96_sum;
  assign calc_dlv_elem_67 = { calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97], calc_fout_int_vld[97] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12094" *) calc_fout_int_97_sum;
  assign calc_dlv_elem_69 = { calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98], calc_fout_int_vld[98] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12095" *) calc_fout_int_98_sum;
  assign calc_dlv_elem_71 = { calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99], calc_fout_int_vld[99] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12096" *) calc_fout_int_99_sum;
  assign calc_dlv_elem_73 = { calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100], calc_fout_int_vld[100] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12097" *) calc_fout_int_100_sum;
  assign calc_dlv_elem_75 = { calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101], calc_fout_int_vld[101] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12098" *) calc_fout_int_101_sum;
  assign calc_dlv_elem_77 = { calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102], calc_fout_int_vld[102] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12099" *) calc_fout_int_102_sum;
  assign calc_dlv_elem_79 = { calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103], calc_fout_int_vld[103] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12100" *) calc_fout_int_103_sum;
  assign calc_dlv_elem_81 = { calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104], calc_fout_int_vld[104] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12101" *) calc_fout_int_104_sum;
  assign calc_dlv_elem_83 = { calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105], calc_fout_int_vld[105] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12102" *) calc_fout_int_105_sum;
  assign calc_dlv_elem_85 = { calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106], calc_fout_int_vld[106] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12103" *) calc_fout_int_106_sum;
  assign calc_dlv_elem_87 = { calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107], calc_fout_int_vld[107] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12104" *) calc_fout_int_107_sum;
  assign calc_dlv_elem_89 = { calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108], calc_fout_int_vld[108] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12105" *) calc_fout_int_108_sum;
  assign calc_dlv_elem_91 = { calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109], calc_fout_int_vld[109] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12106" *) calc_fout_int_109_sum;
  assign calc_dlv_elem_93 = { calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110], calc_fout_int_vld[110] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12107" *) calc_fout_int_110_sum;
  assign calc_dlv_elem_95 = { calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111], calc_fout_int_vld[111] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12108" *) calc_fout_int_111_sum;
  assign calc_dlv_elem_97 = { calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112], calc_fout_int_vld[112] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12109" *) calc_fout_int_112_sum;
  assign calc_dlv_elem_99 = { calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113], calc_fout_int_vld[113] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12110" *) calc_fout_int_113_sum;
  assign calc_dlv_elem_101 = { calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114], calc_fout_int_vld[114] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12111" *) calc_fout_int_114_sum;
  assign calc_dlv_elem_103 = { calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115], calc_fout_int_vld[115] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12112" *) calc_fout_int_115_sum;
  assign calc_dlv_elem_105 = { calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116], calc_fout_int_vld[116] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12113" *) calc_fout_int_116_sum;
  assign calc_dlv_elem_107 = { calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117], calc_fout_int_vld[117] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12114" *) calc_fout_int_117_sum;
  assign calc_dlv_elem_109 = { calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118], calc_fout_int_vld[118] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12115" *) calc_fout_int_118_sum;
  assign calc_dlv_elem_111 = { calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119], calc_fout_int_vld[119] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12116" *) calc_fout_int_119_sum;
  assign calc_dlv_elem_113 = { calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120], calc_fout_int_vld[120] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12117" *) calc_fout_int_120_sum;
  assign calc_dlv_elem_115 = { calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121], calc_fout_int_vld[121] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12118" *) calc_fout_int_121_sum;
  assign calc_dlv_elem_117 = { calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122], calc_fout_int_vld[122] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12119" *) calc_fout_int_122_sum;
  assign calc_dlv_elem_119 = { calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123], calc_fout_int_vld[123] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12120" *) calc_fout_int_123_sum;
  assign calc_dlv_elem_121 = { calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124], calc_fout_int_vld[124] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12121" *) calc_fout_int_124_sum;
  assign calc_dlv_elem_123 = { calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125], calc_fout_int_vld[125] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12122" *) calc_fout_int_125_sum;
  assign calc_dlv_elem_125 = { calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126], calc_fout_int_vld[126] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12123" *) calc_fout_int_126_sum;
  assign calc_dlv_elem_127 = { calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127], calc_fout_int_vld[127] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12124" *) calc_fout_int_127_sum;
  assign dlv_sat_end = calc_layer_end_out & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13266" *) calc_stripe_end_out;
  assign _0863_ = calc_dlv_valid_out & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13267" *) _0898_;
  assign dlv_sat_clr = _0863_ & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13267" *) dlv_sat_end_d1;
  assign sat_reg_en = dlv_sat_vld_d1 & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13420" *) _0902_;
  assign _0864_ = mac_a2accu_mask[0] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2280" *) mac_a2accu_mode[0];
  assign _0865_ = mac_a2accu_mask[1] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2300" *) mac_a2accu_mode[1];
  assign _0866_ = mac_a2accu_mask[2] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2320" *) mac_a2accu_mode[2];
  assign _0867_ = mac_a2accu_mask[3] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2340" *) mac_a2accu_mode[3];
  assign _0868_ = mac_a2accu_mask[4] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2360" *) mac_a2accu_mode[4];
  assign _0869_ = mac_a2accu_mask[5] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2380" *) mac_a2accu_mode[5];
  assign _0870_ = mac_a2accu_mask[6] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2400" *) mac_a2accu_mode[6];
  assign _0871_ = mac_a2accu_mask[7] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2420" *) mac_a2accu_mode[7];
  assign _0872_ = mac_b2accu_mask[0] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2440" *) mac_b2accu_mode[0];
  assign _0873_ = mac_b2accu_mask[1] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2460" *) mac_b2accu_mode[1];
  assign _0874_ = mac_b2accu_mask[2] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2480" *) mac_b2accu_mode[2];
  assign _0875_ = mac_b2accu_mask[3] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2500" *) mac_b2accu_mode[3];
  assign _0876_ = mac_b2accu_mask[4] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2520" *) mac_b2accu_mode[4];
  assign _0877_ = mac_b2accu_mask[5] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2540" *) mac_b2accu_mode[5];
  assign _0878_ = mac_b2accu_mask[6] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2560" *) mac_b2accu_mode[6];
  assign _0879_ = mac_b2accu_mask[7] & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2580" *) mac_b2accu_mode[7];
  assign _0880_ = { accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35:34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34:33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33:32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32:31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31:30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30:29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29:28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28:27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27:26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26:25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25:24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24:23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23:22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22:21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21:20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3138" *) abuf_rd_data_0;
  assign _0881_ = { accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51:50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50:49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49:48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48:47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47:46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46:45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45:44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44:43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43:42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42:41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41:40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40:39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39:38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38:37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37:36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3139" *) abuf_rd_data_1;
  assign _0882_ = { accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67:66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66:65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65:64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64:63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63:62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62:61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61:60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60:59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59:58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58:57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57:56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56:55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55:54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54:53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53:52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3140" *) abuf_rd_data_2;
  assign _0883_ = { accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83:82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82:81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81:80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80:79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79:78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78:77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77:76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76:75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75:74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74:73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73:72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72:71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71:70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70:69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69:68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3141" *) abuf_rd_data_3;
  assign _0884_ = { accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99:98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98:97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97:96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96:95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95:94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94:93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93:92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92:91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91:90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90:89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89:88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88:87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87:86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86:85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85:84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3162" *) abuf_rd_data_4;
  assign _0885_ = { accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115:114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114:113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113:112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112:111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111:110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110:109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109:108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108:107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107:106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106:105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105:104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104:103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103:102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102:101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101:100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3163" *) abuf_rd_data_5;
  assign _0886_ = { accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131:130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130:129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129:128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128:127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127:126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126:125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125:124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124:123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123:122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122:121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121:120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120:119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119:118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118:117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117:116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3164" *) abuf_rd_data_6;
  assign _0887_ = { accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147:146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146:145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145:144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144:143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143:142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142:141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141:140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140:139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139:138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138:137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137:136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136:135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135:134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134:133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133:132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132] } & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3165" *) abuf_rd_data_7;
  assign calc_elem_en = calc_in_mask & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3191" *) cfg_in_en_mask;
  assign calc_elem_op1_vld = calc_elem_en & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3194" *) accu_ctrl_ram_valid;
  assign calc_dlv_elem_en = calc_elem_en & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3197" *) accu_ctrl_pd[339:148];
  assign calc_dlv_valid = accu_ctrl_valid & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3223" *) accu_ctrl_pd[18];
  assign calc_valid_d0 = accu_ctrl_valid & (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3225" *) calc_valid;
  assign _0898_ = ~ (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13267" *) dlv_sat_end;
  assign _0899_ = ~ (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3205" *) calc_valid;
  assign _0900_ = ~ (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3205" *) accu_ctrl_pd[18];
  assign _0901_ = ~ (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3216" *) accu_ctrl_valid;
  assign _0888_ = calc_valid_d1 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10524" *) calc_valid_d2;
  assign _0889_ = calc_valid_d2 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10653" *) calc_valid_d3;
  assign _0890_ = calc_valid_d3 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10782" *) calc_valid_d4;
  assign calc_wr_en_out = _0595_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10903" *) _0596_;
  assign calc_addr_out = _0597_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10905" *) _0598_;
  assign _0891_ = calc_dlv_valid_d1 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10917" *) calc_dlv_valid_d2;
  assign _0892_ = calc_dlv_valid_d2 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11107" *) calc_dlv_valid_d3;
  assign _0893_ = calc_dlv_valid_d3 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11297" *) calc_dlv_valid_d4;
  assign _0894_ = calc_dlv_valid_d4 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11487" *) calc_dlv_valid_d5;
  assign calc_dlv_valid_out = _0599_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11667" *) _0600_;
  assign calc_dlv_en_out = _0601_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11669" *) _0602_;
  assign calc_stripe_end_out = _0603_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11671" *) _0604_;
  assign calc_layer_end_out = _0605_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11673" *) _0606_;
  assign calc_pout_0 = _0607_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11742" *) _0608_;
  assign calc_pout_1 = _0609_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11744" *) _0610_;
  assign calc_pout_2 = _0611_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11746" *) _0612_;
  assign calc_pout_3 = _0613_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11748" *) _0614_;
  assign calc_pout_4 = _0615_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11750" *) _0616_;
  assign calc_pout_5 = _0617_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11752" *) _0618_;
  assign calc_pout_6 = _0619_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11754" *) _0620_;
  assign calc_pout_7 = _0621_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11756" *) _0622_;
  assign calc_pout_8 = _0623_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11758" *) _0624_;
  assign calc_pout_9 = _0625_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11760" *) _0626_;
  assign calc_pout_10 = _0627_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11762" *) _0628_;
  assign calc_pout_11 = _0629_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11764" *) _0630_;
  assign calc_pout_12 = _0631_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11766" *) _0632_;
  assign calc_pout_13 = _0633_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11768" *) _0634_;
  assign calc_pout_14 = _0635_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11770" *) _0636_;
  assign calc_pout_15 = _0637_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11772" *) _0638_;
  assign calc_pout_16 = _0639_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11774" *) _0640_;
  assign calc_pout_17 = _0641_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11776" *) _0642_;
  assign calc_pout_18 = _0643_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11778" *) _0644_;
  assign calc_pout_19 = _0645_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11780" *) _0646_;
  assign calc_pout_20 = _0647_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11782" *) _0648_;
  assign calc_pout_21 = _0649_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11784" *) _0650_;
  assign calc_pout_22 = _0651_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11786" *) _0652_;
  assign calc_pout_23 = _0653_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11788" *) _0654_;
  assign calc_pout_24 = _0655_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11790" *) _0656_;
  assign calc_pout_25 = _0657_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11792" *) _0658_;
  assign calc_pout_26 = _0659_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11794" *) _0660_;
  assign calc_pout_27 = _0661_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11796" *) _0662_;
  assign calc_pout_28 = _0663_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11798" *) _0664_;
  assign calc_pout_29 = _0665_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11800" *) _0666_;
  assign calc_pout_30 = _0667_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11802" *) _0668_;
  assign calc_pout_31 = _0669_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11804" *) _0670_;
  assign calc_pout_32 = _0671_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11806" *) _0672_;
  assign calc_pout_33 = _0673_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11808" *) _0674_;
  assign calc_pout_34 = _0675_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11810" *) _0676_;
  assign calc_pout_35 = _0677_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11812" *) _0678_;
  assign calc_pout_36 = _0679_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11814" *) _0680_;
  assign calc_pout_37 = _0681_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11816" *) _0682_;
  assign calc_pout_38 = _0683_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11818" *) _0684_;
  assign calc_pout_39 = _0685_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11820" *) _0686_;
  assign calc_pout_40 = _0687_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11822" *) _0688_;
  assign calc_pout_41 = _0689_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11824" *) _0690_;
  assign calc_pout_42 = _0691_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11826" *) _0692_;
  assign calc_pout_43 = _0693_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11828" *) _0694_;
  assign calc_pout_44 = _0695_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11830" *) _0696_;
  assign calc_pout_45 = _0697_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11832" *) _0698_;
  assign calc_pout_46 = _0699_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11834" *) _0700_;
  assign calc_pout_47 = _0701_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11836" *) _0702_;
  assign calc_pout_48 = _0703_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11838" *) _0704_;
  assign calc_pout_49 = _0705_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11840" *) _0706_;
  assign calc_pout_50 = _0707_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11842" *) _0708_;
  assign calc_pout_51 = _0709_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11844" *) _0710_;
  assign calc_pout_52 = _0711_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11846" *) _0712_;
  assign calc_pout_53 = _0713_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11848" *) _0714_;
  assign calc_pout_54 = _0715_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11850" *) _0716_;
  assign calc_pout_55 = _0717_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11852" *) _0718_;
  assign calc_pout_56 = _0719_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11854" *) _0720_;
  assign calc_pout_57 = _0721_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11856" *) _0722_;
  assign calc_pout_58 = _0723_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11858" *) _0724_;
  assign calc_pout_59 = _0725_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11860" *) _0726_;
  assign calc_pout_60 = _0727_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11862" *) _0728_;
  assign calc_pout_61 = _0729_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11864" *) _0730_;
  assign calc_pout_62 = _0731_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11866" *) _0732_;
  assign calc_pout_63 = _0733_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11868" *) _0734_;
  assign calc_dlv_elem_0 = _0735_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11934" *) _0736_;
  assign calc_fout_1 = _0737_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11936" *) _0738_;
  assign calc_fout_2 = _0739_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11938" *) _0740_;
  assign calc_fout_3 = _0741_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11940" *) _0742_;
  assign calc_fout_4 = _0743_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11942" *) _0744_;
  assign calc_fout_5 = _0745_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11944" *) _0746_;
  assign calc_fout_6 = _0747_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11946" *) _0748_;
  assign calc_fout_7 = _0749_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11948" *) _0750_;
  assign calc_fout_8 = _0751_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11950" *) _0752_;
  assign calc_fout_9 = _0753_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11952" *) _0754_;
  assign calc_fout_10 = _0755_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11954" *) _0756_;
  assign calc_fout_11 = _0757_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11956" *) _0758_;
  assign calc_fout_12 = _0759_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11958" *) _0760_;
  assign calc_fout_13 = _0761_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11960" *) _0762_;
  assign calc_fout_14 = _0763_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11962" *) _0764_;
  assign calc_fout_15 = _0765_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11964" *) _0766_;
  assign calc_fout_16 = _0767_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11966" *) _0768_;
  assign calc_fout_17 = _0769_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11968" *) _0770_;
  assign calc_fout_18 = _0771_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11970" *) _0772_;
  assign calc_fout_19 = _0773_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11972" *) _0774_;
  assign calc_fout_20 = _0775_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11974" *) _0776_;
  assign calc_fout_21 = _0777_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11976" *) _0778_;
  assign calc_fout_22 = _0779_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11978" *) _0780_;
  assign calc_fout_23 = _0781_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11980" *) _0782_;
  assign calc_fout_24 = _0783_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11982" *) _0784_;
  assign calc_fout_25 = _0785_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11984" *) _0786_;
  assign calc_fout_26 = _0787_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11986" *) _0788_;
  assign calc_fout_27 = _0789_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11988" *) _0790_;
  assign calc_fout_28 = _0791_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11990" *) _0792_;
  assign calc_fout_29 = _0793_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11992" *) _0794_;
  assign calc_fout_30 = _0795_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11994" *) _0796_;
  assign calc_fout_31 = _0797_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11996" *) _0798_;
  assign calc_fout_32 = _0799_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11998" *) _0800_;
  assign calc_fout_33 = _0801_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12000" *) _0802_;
  assign calc_fout_34 = _0803_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12002" *) _0804_;
  assign calc_fout_35 = _0805_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12004" *) _0806_;
  assign calc_fout_36 = _0807_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12006" *) _0808_;
  assign calc_fout_37 = _0809_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12008" *) _0810_;
  assign calc_fout_38 = _0811_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12010" *) _0812_;
  assign calc_fout_39 = _0813_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12012" *) _0814_;
  assign calc_fout_40 = _0815_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12014" *) _0816_;
  assign calc_fout_41 = _0817_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12016" *) _0818_;
  assign calc_fout_42 = _0819_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12018" *) _0820_;
  assign calc_fout_43 = _0821_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12020" *) _0822_;
  assign calc_fout_44 = _0823_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12022" *) _0824_;
  assign calc_fout_45 = _0825_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12024" *) _0826_;
  assign calc_fout_46 = _0827_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12026" *) _0828_;
  assign calc_fout_47 = _0829_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12028" *) _0830_;
  assign calc_fout_48 = _0831_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12030" *) _0832_;
  assign calc_fout_49 = _0833_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12032" *) _0834_;
  assign calc_fout_50 = _0835_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12034" *) _0836_;
  assign calc_fout_51 = _0837_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12036" *) _0838_;
  assign calc_fout_52 = _0839_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12038" *) _0840_;
  assign calc_fout_53 = _0841_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12040" *) _0842_;
  assign calc_fout_54 = _0843_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12042" *) _0844_;
  assign calc_fout_55 = _0845_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12044" *) _0846_;
  assign calc_fout_56 = _0847_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12046" *) _0848_;
  assign calc_fout_57 = _0849_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12048" *) _0850_;
  assign calc_fout_58 = _0851_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12050" *) _0852_;
  assign calc_fout_59 = _0853_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12052" *) _0854_;
  assign calc_fout_60 = _0855_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12054" *) _0856_;
  assign calc_fout_61 = _0857_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12056" *) _0858_;
  assign calc_fout_62 = _0859_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12058" *) _0860_;
  assign calc_fout_63 = _0861_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12060" *) _0862_;
  assign _0902_ = _0909_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13420" *) dlv_sat_clr_d1;
  assign calc_valid_fw_0 = mac_b2accu_pvld | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2589" *) mac_a2accu_pvld;
  assign _0896_ = calc_valid_fw_3 | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2616" *) calc_valid;
  assign _0903_ = _0880_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3139" *) _0881_;
  assign _0904_ = _0903_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3140" *) _0882_;
  assign abuf_rd_data_0_sft = _0904_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3141" *) _0883_;
  assign _0905_ = _0884_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3163" *) _0885_;
  assign _0906_ = _0905_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3164" *) _0886_;
  assign abuf_rd_data_4_sft = _0906_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3165" *) _0887_;
  assign _0907_ = _0899_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3205" *) _0900_;
  assign _0908_ = _0901_ | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3216" *) accu_ctrl_pd[18];
  assign _0897_ = accu_ctrl_valid | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7080" *) calc_valid_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      sat_count <= 32'd0;
    else
      sat_count <= _0468_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_sat_clr_d1 <= 1'b0;
    else
      dlv_sat_clr_d1 <= dlv_sat_clr;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_sat_bit_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      dlv_sat_bit_d1 <= _0465_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_sat_end_d1 <= 1'b1;
    else
      dlv_sat_end_d1 <= _0466_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_sat_vld_d1 <= 1'b0;
    else
      dlv_sat_vld_d1 <= calc_dlv_valid_out;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_layer_end <= 1'b0;
    else
      dlv_layer_end <= _0463_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_stripe_end <= 1'b0;
    else
      dlv_stripe_end <= _0467_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      dlv_mask <= 8'b00000000;
    else
      dlv_mask <= _0464_;
  always @(posedge nvdla_core_clk)
      dlv_data_7 <= _0462_;
  always @(posedge nvdla_core_clk)
      dlv_data_6 <= _0461_;
  always @(posedge nvdla_core_clk)
      dlv_data_5 <= _0460_;
  always @(posedge nvdla_core_clk)
      dlv_data_4 <= _0459_;
  always @(posedge nvdla_core_clk)
      dlv_data_3 <= _0458_;
  always @(posedge nvdla_core_clk)
      dlv_data_2 <= _0457_;
  always @(posedge nvdla_core_clk)
      dlv_data_1 <= _0456_;
  always @(posedge nvdla_core_clk)
      dlv_data_0 <= _0455_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_7 <= _0008_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_6 <= _0007_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_5 <= _0006_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_4 <= _0005_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_3 <= _0004_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_2 <= _0003_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_1 <= _0002_;
  always @(posedge nvdla_core_clk)
      abuf_wr_data_0 <= _0001_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      abuf_wr_addr <= 5'b00000;
    else
      abuf_wr_addr <= _0000_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      abuf_wr_en <= 8'b00000000;
    else
      abuf_wr_en <= calc_wr_en_out;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_layer_end_d5 <= 1'b0;
    else
      calc_layer_end_d5 <= _0057_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_stripe_end_d5 <= 1'b0;
    else
      calc_stripe_end_d5 <= _0450_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_d5 <= 8'b00000000;
    else
      calc_dlv_en_d5 <= _0049_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_valid_d5 <= 1'b0;
    else
      calc_dlv_valid_d5 <= calc_dlv_valid_d4;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_layer_end_d4 <= 1'b0;
    else
      calc_layer_end_d4 <= _0056_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_stripe_end_d4 <= 1'b0;
    else
      calc_stripe_end_d4 <= _0449_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_d4 <= 8'b00000000;
    else
      calc_dlv_en_d4 <= _0048_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_valid_d4 <= 1'b0;
    else
      calc_dlv_valid_d4 <= calc_dlv_valid_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_layer_end_d3 <= 1'b0;
    else
      calc_layer_end_d3 <= _0055_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_stripe_end_d3 <= 1'b0;
    else
      calc_stripe_end_d3 <= _0448_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_d3 <= 8'b00000000;
    else
      calc_dlv_en_d3 <= _0047_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_valid_d3 <= 1'b0;
    else
      calc_dlv_valid_d3 <= calc_dlv_valid_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_layer_end_d2 <= 1'b0;
    else
      calc_layer_end_d2 <= _0054_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_stripe_end_d2 <= 1'b0;
    else
      calc_stripe_end_d2 <= _0447_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_d2 <= 8'b00000000;
    else
      calc_dlv_en_d2 <= _0046_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_valid_d2 <= 1'b0;
    else
      calc_dlv_valid_d2 <= calc_dlv_valid_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_addr_d4 <= 5'b00000;
    else
      calc_addr_d4 <= _0012_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_wr_en_d4 <= 8'b00000000;
    else
      calc_wr_en_d4 <= _0454_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_d4 <= 1'b0;
    else
      calc_valid_d4 <= calc_valid_d3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_addr_d3 <= 5'b00000;
    else
      calc_addr_d3 <= _0011_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_wr_en_d3 <= 8'b00000000;
    else
      calc_wr_en_d3 <= _0453_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_d3 <= 1'b0;
    else
      calc_valid_d3 <= calc_valid_d2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_addr_d2 <= 5'b00000;
    else
      calc_addr_d2 <= _0010_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_wr_en_d2 <= 8'b00000000;
    else
      calc_wr_en_d2 <= _0452_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_d2 <= 1'b0;
    else
      calc_valid_d2 <= calc_valid_d1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_fp_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_dlv_en_fp_d1 <= _0050_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_int_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_dlv_en_int_d1 <= _0051_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_op1_vld_fp_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_op1_vld_fp_d1 <= _0442_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_op1_vld_int_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_op1_vld_int_d1 <= _0443_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_op_en_fp_d1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_op_en_fp_d1 <= _0444_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_op_en_int_d1 <= 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_op_en_int_d1 <= _0445_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_layer_end_d1 <= 1'b0;
    else
      calc_layer_end_d1 <= _0053_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_stripe_end_d1 <= 1'b0;
    else
      calc_stripe_end_d1 <= _0446_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_en_d1 <= 8'b00000000;
    else
      calc_dlv_en_d1 <= _0045_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_dlv_valid_d1 <= 1'b0;
    else
      calc_dlv_valid_d1 <= calc_dlv_valid;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_addr_d1 <= 5'b00000;
    else
      calc_addr_d1 <= _0009_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_wr_en_d1 <= 8'b00000000;
    else
      calc_wr_en_d1 <= _0451_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_d1 <= 1'b0;
    else
      calc_valid_d1 <= calc_valid_d0;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_63_d1 <= _0309_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_62_d1 <= _0308_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_61_d1 <= _0307_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_60_d1 <= _0306_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_59_d1 <= _0304_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_58_d1 <= _0303_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_57_d1 <= _0302_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_56_d1 <= _0301_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_55_d1 <= _0300_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_54_d1 <= _0299_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_53_d1 <= _0298_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_52_d1 <= _0297_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_51_d1 <= _0296_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_50_d1 <= _0295_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_49_d1 <= _0293_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_48_d1 <= _0292_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_47_d1 <= _0291_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_46_d1 <= _0290_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_45_d1 <= _0289_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_44_d1 <= _0288_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_43_d1 <= _0287_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_42_d1 <= _0286_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_41_d1 <= _0285_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_40_d1 <= _0284_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_39_d1 <= _0282_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_38_d1 <= _0281_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_37_d1 <= _0280_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_36_d1 <= _0279_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_35_d1 <= _0278_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_34_d1 <= _0277_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_33_d1 <= _0276_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_32_d1 <= _0275_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_31_d1 <= _0274_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_30_d1 <= _0273_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_29_d1 <= _0271_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_28_d1 <= _0270_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_27_d1 <= _0269_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_26_d1 <= _0268_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_25_d1 <= _0267_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_24_d1 <= _0266_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_23_d1 <= _0265_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_22_d1 <= _0264_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_21_d1 <= _0263_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_20_d1 <= _0262_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_19_d1 <= _0260_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_18_d1 <= _0259_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_17_d1 <= _0258_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_16_d1 <= _0257_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_15_d1 <= _0256_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_14_d1 <= _0255_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_13_d1 <= _0254_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_12_d1 <= _0253_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_11_d1 <= _0252_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_10_d1 <= _0251_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_9_d1 <= _0313_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_8_d1 <= _0312_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_7_d1 <= _0311_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_6_d1 <= _0310_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_5_d1 <= _0305_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_4_d1 <= _0294_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_3_d1 <= _0283_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_2_d1 <= _0272_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_1_d1 <= _0261_;
  always @(posedge nvdla_core_clk)
      calc_op1_fp_0_d1 <= _0250_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_127_d1 <= _0344_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_126_d1 <= _0343_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_125_d1 <= _0342_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_124_d1 <= _0341_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_123_d1 <= _0340_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_122_d1 <= _0339_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_121_d1 <= _0338_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_120_d1 <= _0337_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_119_d1 <= _0335_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_118_d1 <= _0334_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_117_d1 <= _0333_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_116_d1 <= _0332_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_115_d1 <= _0331_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_114_d1 <= _0330_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_113_d1 <= _0329_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_112_d1 <= _0328_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_111_d1 <= _0327_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_110_d1 <= _0326_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_109_d1 <= _0324_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_108_d1 <= _0323_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_107_d1 <= _0322_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_106_d1 <= _0321_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_105_d1 <= _0320_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_104_d1 <= _0319_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_103_d1 <= _0318_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_102_d1 <= _0317_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_101_d1 <= _0316_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_100_d1 <= _0315_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_99_d1 <= _0440_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_98_d1 <= _0439_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_97_d1 <= _0438_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_96_d1 <= _0437_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_95_d1 <= _0436_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_94_d1 <= _0435_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_93_d1 <= _0434_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_92_d1 <= _0433_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_91_d1 <= _0432_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_90_d1 <= _0431_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_89_d1 <= _0429_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_88_d1 <= _0428_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_87_d1 <= _0427_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_86_d1 <= _0426_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_85_d1 <= _0425_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_84_d1 <= _0424_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_83_d1 <= _0423_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_82_d1 <= _0422_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_81_d1 <= _0421_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_80_d1 <= _0420_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_79_d1 <= _0418_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_78_d1 <= _0417_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_77_d1 <= _0416_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_76_d1 <= _0415_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_75_d1 <= _0414_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_74_d1 <= _0413_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_73_d1 <= _0412_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_72_d1 <= _0411_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_71_d1 <= _0410_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_70_d1 <= _0409_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_69_d1 <= _0407_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_68_d1 <= _0406_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_67_d1 <= _0405_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_66_d1 <= _0404_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_65_d1 <= _0403_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_64_d1 <= _0402_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_63_d1 <= _0401_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_62_d1 <= _0400_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_61_d1 <= _0399_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_60_d1 <= _0398_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_59_d1 <= _0396_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_58_d1 <= _0395_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_57_d1 <= _0394_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_56_d1 <= _0393_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_55_d1 <= _0392_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_54_d1 <= _0391_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_53_d1 <= _0390_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_52_d1 <= _0389_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_51_d1 <= _0388_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_50_d1 <= _0387_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_49_d1 <= _0385_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_48_d1 <= _0384_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_47_d1 <= _0383_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_46_d1 <= _0382_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_45_d1 <= _0381_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_44_d1 <= _0380_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_43_d1 <= _0379_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_42_d1 <= _0378_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_41_d1 <= _0377_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_40_d1 <= _0376_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_39_d1 <= _0374_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_38_d1 <= _0373_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_37_d1 <= _0372_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_36_d1 <= _0371_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_35_d1 <= _0370_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_34_d1 <= _0369_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_33_d1 <= _0368_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_32_d1 <= _0367_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_31_d1 <= _0366_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_30_d1 <= _0365_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_29_d1 <= _0363_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_28_d1 <= _0362_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_27_d1 <= _0361_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_26_d1 <= _0360_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_25_d1 <= _0359_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_24_d1 <= _0358_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_23_d1 <= _0357_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_22_d1 <= _0356_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_21_d1 <= _0355_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_20_d1 <= _0354_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_19_d1 <= _0352_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_18_d1 <= _0351_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_17_d1 <= _0350_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_16_d1 <= _0349_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_15_d1 <= _0348_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_14_d1 <= _0347_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_13_d1 <= _0346_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_12_d1 <= _0345_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_11_d1 <= _0336_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_10_d1 <= _0325_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_9_d1 <= _0441_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_8_d1 <= _0430_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_7_d1 <= _0419_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_6_d1 <= _0408_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_5_d1 <= _0397_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_4_d1 <= _0386_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_3_d1 <= _0375_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_2_d1 <= _0364_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_1_d1 <= _0353_;
  always @(posedge nvdla_core_clk)
      calc_op1_int_0_d1 <= _0314_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_63_d1 <= _0117_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_62_d1 <= _0116_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_61_d1 <= _0115_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_60_d1 <= _0114_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_59_d1 <= _0112_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_58_d1 <= _0111_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_57_d1 <= _0110_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_56_d1 <= _0109_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_55_d1 <= _0108_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_54_d1 <= _0107_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_53_d1 <= _0106_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_52_d1 <= _0105_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_51_d1 <= _0104_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_50_d1 <= _0103_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_49_d1 <= _0101_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_48_d1 <= _0100_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_47_d1 <= _0099_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_46_d1 <= _0098_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_45_d1 <= _0097_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_44_d1 <= _0096_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_43_d1 <= _0095_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_42_d1 <= _0094_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_41_d1 <= _0093_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_40_d1 <= _0092_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_39_d1 <= _0090_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_38_d1 <= _0089_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_37_d1 <= _0088_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_36_d1 <= _0087_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_35_d1 <= _0086_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_34_d1 <= _0085_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_33_d1 <= _0084_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_32_d1 <= _0083_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_31_d1 <= _0082_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_30_d1 <= _0081_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_29_d1 <= _0079_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_28_d1 <= _0078_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_27_d1 <= _0077_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_26_d1 <= _0076_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_25_d1 <= _0075_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_24_d1 <= _0074_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_23_d1 <= _0073_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_22_d1 <= _0072_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_21_d1 <= _0071_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_20_d1 <= _0070_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_19_d1 <= _0068_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_18_d1 <= _0067_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_17_d1 <= _0066_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_16_d1 <= _0065_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_15_d1 <= _0064_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_14_d1 <= _0063_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_13_d1 <= _0062_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_12_d1 <= _0061_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_11_d1 <= _0060_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_10_d1 <= _0059_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_9_d1 <= _0121_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_8_d1 <= _0120_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_7_d1 <= _0119_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_6_d1 <= _0118_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_5_d1 <= _0113_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_4_d1 <= _0102_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_3_d1 <= _0091_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_2_d1 <= _0080_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_1_d1 <= _0069_;
  always @(posedge nvdla_core_clk)
      calc_op0_fp_0_d1 <= _0058_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_127_d1 <= _0152_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_126_d1 <= _0151_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_125_d1 <= _0150_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_124_d1 <= _0149_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_123_d1 <= _0148_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_122_d1 <= _0147_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_121_d1 <= _0146_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_120_d1 <= _0145_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_119_d1 <= _0143_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_118_d1 <= _0142_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_117_d1 <= _0141_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_116_d1 <= _0140_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_115_d1 <= _0139_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_114_d1 <= _0138_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_113_d1 <= _0137_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_112_d1 <= _0136_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_111_d1 <= _0135_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_110_d1 <= _0134_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_109_d1 <= _0132_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_108_d1 <= _0131_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_107_d1 <= _0130_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_106_d1 <= _0129_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_105_d1 <= _0128_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_104_d1 <= _0127_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_103_d1 <= _0126_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_102_d1 <= _0125_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_101_d1 <= _0124_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_100_d1 <= _0123_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_99_d1 <= _0248_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_98_d1 <= _0247_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_97_d1 <= _0246_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_96_d1 <= _0245_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_95_d1 <= _0244_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_94_d1 <= _0243_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_93_d1 <= _0242_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_92_d1 <= _0241_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_91_d1 <= _0240_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_90_d1 <= _0239_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_89_d1 <= _0237_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_88_d1 <= _0236_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_87_d1 <= _0235_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_86_d1 <= _0234_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_85_d1 <= _0233_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_84_d1 <= _0232_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_83_d1 <= _0231_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_82_d1 <= _0230_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_81_d1 <= _0229_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_80_d1 <= _0228_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_79_d1 <= _0226_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_78_d1 <= _0225_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_77_d1 <= _0224_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_76_d1 <= _0223_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_75_d1 <= _0222_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_74_d1 <= _0221_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_73_d1 <= _0220_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_72_d1 <= _0219_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_71_d1 <= _0218_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_70_d1 <= _0217_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_69_d1 <= _0215_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_68_d1 <= _0214_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_67_d1 <= _0213_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_66_d1 <= _0212_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_65_d1 <= _0211_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_64_d1 <= _0210_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_63_d1 <= _0209_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_62_d1 <= _0208_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_61_d1 <= _0207_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_60_d1 <= _0206_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_59_d1 <= _0204_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_58_d1 <= _0203_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_57_d1 <= _0202_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_56_d1 <= _0201_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_55_d1 <= _0200_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_54_d1 <= _0199_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_53_d1 <= _0198_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_52_d1 <= _0197_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_51_d1 <= _0196_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_50_d1 <= _0195_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_49_d1 <= _0193_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_48_d1 <= _0192_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_47_d1 <= _0191_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_46_d1 <= _0190_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_45_d1 <= _0189_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_44_d1 <= _0188_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_43_d1 <= _0187_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_42_d1 <= _0186_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_41_d1 <= _0185_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_40_d1 <= _0184_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_39_d1 <= _0182_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_38_d1 <= _0181_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_37_d1 <= _0180_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_36_d1 <= _0179_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_35_d1 <= _0178_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_34_d1 <= _0177_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_33_d1 <= _0176_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_32_d1 <= _0175_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_31_d1 <= _0174_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_30_d1 <= _0173_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_29_d1 <= _0171_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_28_d1 <= _0170_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_27_d1 <= _0169_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_26_d1 <= _0168_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_25_d1 <= _0167_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_24_d1 <= _0166_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_23_d1 <= _0165_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_22_d1 <= _0164_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_21_d1 <= _0163_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_20_d1 <= _0162_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_19_d1 <= _0160_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_18_d1 <= _0159_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_17_d1 <= _0158_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_16_d1 <= _0157_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_15_d1 <= _0156_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_14_d1 <= _0155_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_13_d1 <= _0154_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_12_d1 <= _0153_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_11_d1 <= _0144_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_10_d1 <= _0133_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_9_d1 <= _0249_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_8_d1 <= _0238_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_7_d1 <= _0227_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_6_d1 <= _0216_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_5_d1 <= _0205_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_4_d1 <= _0194_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_3_d1 <= _0183_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_2_d1 <= _0172_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_1_d1 <= _0161_;
  always @(posedge nvdla_core_clk)
      calc_op0_int_0_d1 <= _0122_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid <= 1'b0;
    else
      calc_valid <= calc_valid_fw_3;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_in_mask <= 192'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    else
      calc_in_mask <= _0052_;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_fw_3 <= 1'b0;
    else
      calc_valid_fw_3 <= calc_valid_fw_2;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_fw_2 <= 1'b0;
    else
      calc_valid_fw_2 <= calc_valid_fw_1;
  always @(posedge nvdla_core_clk or negedge nvdla_core_rstn)
    if (!nvdla_core_rstn)
      calc_valid_fw_1 <= 1'b0;
    else
      calc_valid_fw_1 <= calc_valid_fw_0;
  always @(posedge nvdla_core_clk)
      calc_data_15[175:44] <= _0025_;
  always @(posedge nvdla_core_clk)
      calc_data_15[43:0] <= _0026_;
  always @(posedge nvdla_core_clk)
      calc_data_14[175:44] <= _0023_;
  always @(posedge nvdla_core_clk)
      calc_data_14[43:0] <= _0024_;
  always @(posedge nvdla_core_clk)
      calc_data_13[175:44] <= _0021_;
  always @(posedge nvdla_core_clk)
      calc_data_13[43:0] <= _0022_;
  always @(posedge nvdla_core_clk)
      calc_data_12[175:44] <= _0019_;
  always @(posedge nvdla_core_clk)
      calc_data_12[43:0] <= _0020_;
  always @(posedge nvdla_core_clk)
      calc_data_11[175:44] <= _0017_;
  always @(posedge nvdla_core_clk)
      calc_data_11[43:0] <= _0018_;
  always @(posedge nvdla_core_clk)
      calc_data_10[175:44] <= _0015_;
  always @(posedge nvdla_core_clk)
      calc_data_10[43:0] <= _0016_;
  always @(posedge nvdla_core_clk)
      calc_data_9[175:44] <= _0043_;
  always @(posedge nvdla_core_clk)
      calc_data_9[43:0] <= _0044_;
  always @(posedge nvdla_core_clk)
      calc_data_8[175:44] <= _0041_;
  always @(posedge nvdla_core_clk)
      calc_data_8[43:0] <= _0042_;
  always @(posedge nvdla_core_clk)
      calc_data_7[175:44] <= _0039_;
  always @(posedge nvdla_core_clk)
      calc_data_7[43:0] <= _0040_;
  always @(posedge nvdla_core_clk)
      calc_data_6[175:44] <= _0037_;
  always @(posedge nvdla_core_clk)
      calc_data_6[43:0] <= _0038_;
  always @(posedge nvdla_core_clk)
      calc_data_5[175:44] <= _0035_;
  always @(posedge nvdla_core_clk)
      calc_data_5[43:0] <= _0036_;
  always @(posedge nvdla_core_clk)
      calc_data_4[175:44] <= _0033_;
  always @(posedge nvdla_core_clk)
      calc_data_4[43:0] <= _0034_;
  always @(posedge nvdla_core_clk)
      calc_data_3[175:44] <= _0031_;
  always @(posedge nvdla_core_clk)
      calc_data_3[43:0] <= _0032_;
  always @(posedge nvdla_core_clk)
      calc_data_2[175:44] <= _0029_;
  always @(posedge nvdla_core_clk)
      calc_data_2[43:0] <= _0030_;
  always @(posedge nvdla_core_clk)
      calc_data_1[175:44] <= _0027_;
  always @(posedge nvdla_core_clk)
      calc_data_1[43:0] <= _0028_;
  always @(posedge nvdla_core_clk)
      calc_data_0[175:44] <= _0013_;
  always @(posedge nvdla_core_clk)
      calc_data_0[43:0] <= _0014_;
  assign _0468_ = sat_reg_en ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13425" *) sat_count_w : sat_count;
  assign _0465_ = calc_dlv_valid_out ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13340" *) calc_fout_int_sat : dlv_sat_bit_d1;
  assign _0466_ = calc_dlv_valid_out ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13279" *) dlv_sat_end : dlv_sat_end_d1;
  assign _0463_ = calc_dlv_valid_out ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13202" *) calc_layer_end_out : dlv_layer_end;
  assign _0467_ = calc_dlv_valid_out ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13141" *) calc_stripe_end_out : dlv_stripe_end;
  assign _0464_ = calc_dlv_valid_out ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13080" *) calc_dlv_en_out : dlv_mask;
  assign _0462_ = calc_dlv_en_out[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13060" *) { calc_dlv_elem_127, calc_fout_63, calc_dlv_elem_125, calc_fout_62, calc_dlv_elem_123, calc_fout_61, calc_dlv_elem_121, calc_fout_60, calc_dlv_elem_119, calc_fout_59, calc_dlv_elem_117, calc_fout_58, calc_dlv_elem_115, calc_fout_57, calc_dlv_elem_113, calc_fout_56 } : dlv_data_7;
  assign _0461_ = calc_dlv_en_out[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13050" *) { calc_dlv_elem_111, calc_fout_55, calc_dlv_elem_109, calc_fout_54, calc_dlv_elem_107, calc_fout_53, calc_dlv_elem_105, calc_fout_52, calc_dlv_elem_103, calc_fout_51, calc_dlv_elem_101, calc_fout_50, calc_dlv_elem_99, calc_fout_49, calc_dlv_elem_97, calc_fout_48 } : dlv_data_6;
  assign _0460_ = calc_dlv_en_out[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13040" *) { calc_dlv_elem_95, calc_fout_47, calc_dlv_elem_93, calc_fout_46, calc_dlv_elem_91, calc_fout_45, calc_dlv_elem_89, calc_fout_44, calc_dlv_elem_87, calc_fout_43, calc_dlv_elem_85, calc_fout_42, calc_dlv_elem_83, calc_fout_41, calc_dlv_elem_81, calc_fout_40 } : dlv_data_5;
  assign _0459_ = calc_dlv_en_out[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13030" *) { calc_dlv_elem_79, calc_fout_39, calc_dlv_elem_77, calc_fout_38, calc_dlv_elem_75, calc_fout_37, calc_dlv_elem_73, calc_fout_36, calc_dlv_elem_71, calc_fout_35, calc_dlv_elem_69, calc_fout_34, calc_dlv_elem_67, calc_fout_33, calc_dlv_elem_65, calc_fout_32 } : dlv_data_4;
  assign _0458_ = calc_dlv_en_out[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13020" *) { calc_dlv_elem_63, calc_dlv_elem_62, calc_dlv_elem_61, calc_dlv_elem_60, calc_dlv_elem_59, calc_dlv_elem_58, calc_dlv_elem_57, calc_dlv_elem_56, calc_dlv_elem_55, calc_dlv_elem_54, calc_dlv_elem_53, calc_dlv_elem_52, calc_dlv_elem_51, calc_dlv_elem_50, calc_dlv_elem_49, calc_dlv_elem_48 } : dlv_data_3;
  assign _0457_ = calc_dlv_en_out[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13010" *) { calc_dlv_elem_47, calc_dlv_elem_46, calc_dlv_elem_45, calc_dlv_elem_44, calc_dlv_elem_43, calc_dlv_elem_42, calc_dlv_elem_41, calc_dlv_elem_40, calc_dlv_elem_39, calc_dlv_elem_38, calc_dlv_elem_37, calc_dlv_elem_36, calc_dlv_elem_35, calc_dlv_elem_34, calc_dlv_elem_33, calc_dlv_elem_32 } : dlv_data_2;
  assign _0456_ = calc_dlv_en_out[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13000" *) { calc_dlv_elem_31, calc_dlv_elem_30, calc_dlv_elem_29, calc_dlv_elem_28, calc_dlv_elem_27, calc_dlv_elem_26, calc_dlv_elem_25, calc_dlv_elem_24, calc_dlv_elem_23, calc_dlv_elem_22, calc_dlv_elem_21, calc_dlv_elem_20, calc_dlv_elem_19, calc_dlv_elem_18, calc_dlv_elem_17, calc_dlv_elem_16 } : dlv_data_1;
  assign _0455_ = calc_dlv_en_out[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12990" *) { calc_dlv_elem_15, calc_dlv_elem_14, calc_dlv_elem_13, calc_dlv_elem_12, calc_dlv_elem_11, calc_dlv_elem_10, calc_dlv_elem_9, calc_dlv_elem_8, calc_dlv_elem_7, calc_dlv_elem_6, calc_dlv_elem_5, calc_dlv_elem_4, calc_dlv_elem_3, calc_dlv_elem_2, calc_dlv_elem_1, calc_dlv_elem_0 } : dlv_data_0;
  assign _0008_ = calc_wr_en_out[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12716" *) { abuf_wr_elem_127, abuf_wr_elem_126, abuf_wr_elem_125, abuf_wr_elem_124, abuf_wr_elem_123, abuf_wr_elem_122, abuf_wr_elem_121, abuf_wr_elem_120, abuf_wr_elem_119, abuf_wr_elem_118, abuf_wr_elem_117, abuf_wr_elem_116, abuf_wr_elem_115, abuf_wr_elem_114, abuf_wr_elem_113, abuf_wr_elem_112 } : abuf_wr_data_7;
  assign _0007_ = calc_wr_en_out[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12706" *) { abuf_wr_elem_111, abuf_wr_elem_110, abuf_wr_elem_109, abuf_wr_elem_108, abuf_wr_elem_107, abuf_wr_elem_106, abuf_wr_elem_105, abuf_wr_elem_104, abuf_wr_elem_103, abuf_wr_elem_102, abuf_wr_elem_101, abuf_wr_elem_100, abuf_wr_elem_99, abuf_wr_elem_98, abuf_wr_elem_97, abuf_wr_elem_96 } : abuf_wr_data_6;
  assign _0006_ = calc_wr_en_out[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12696" *) { abuf_wr_elem_95, abuf_wr_elem_94, abuf_wr_elem_93, abuf_wr_elem_92, abuf_wr_elem_91, abuf_wr_elem_90, abuf_wr_elem_89, abuf_wr_elem_88, abuf_wr_elem_87, abuf_wr_elem_86, abuf_wr_elem_85, abuf_wr_elem_84, abuf_wr_elem_83, abuf_wr_elem_82, abuf_wr_elem_81, abuf_wr_elem_80 } : abuf_wr_data_5;
  assign _0005_ = calc_wr_en_out[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12686" *) { calc_pout_79, calc_pout_78, calc_pout_77, calc_pout_76, calc_pout_75, calc_pout_74, calc_pout_73, calc_pout_72, calc_pout_71, calc_pout_70, calc_pout_69, calc_pout_68, calc_pout_67, calc_pout_66, calc_pout_65, calc_pout_64 } : abuf_wr_data_4;
  assign _0004_ = calc_wr_en_out[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12676" *) { abuf_wr_elem_63, abuf_wr_elem_62, abuf_wr_elem_61, abuf_wr_elem_60, abuf_wr_elem_59, abuf_wr_elem_58, abuf_wr_elem_57, abuf_wr_elem_56, abuf_wr_elem_55, abuf_wr_elem_54, abuf_wr_elem_53, abuf_wr_elem_52, abuf_wr_elem_51, abuf_wr_elem_50, abuf_wr_elem_49, abuf_wr_elem_48 } : abuf_wr_data_3;
  assign _0003_ = calc_wr_en_out[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12666" *) { abuf_wr_elem_47, abuf_wr_elem_46, abuf_wr_elem_45, abuf_wr_elem_44, abuf_wr_elem_43, abuf_wr_elem_42, abuf_wr_elem_41, abuf_wr_elem_40, abuf_wr_elem_39, abuf_wr_elem_38, abuf_wr_elem_37, abuf_wr_elem_36, abuf_wr_elem_35, abuf_wr_elem_34, abuf_wr_elem_33, abuf_wr_elem_32 } : abuf_wr_data_2;
  assign _0002_ = calc_wr_en_out[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12656" *) { abuf_wr_elem_31, abuf_wr_elem_30, abuf_wr_elem_29, abuf_wr_elem_28, abuf_wr_elem_27, abuf_wr_elem_26, abuf_wr_elem_25, abuf_wr_elem_24, abuf_wr_elem_23, abuf_wr_elem_22, abuf_wr_elem_21, abuf_wr_elem_20, abuf_wr_elem_19, abuf_wr_elem_18, abuf_wr_elem_17, abuf_wr_elem_16 } : abuf_wr_data_1;
  assign _0001_ = calc_wr_en_out[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12646" *) { calc_pout_15, calc_pout_14, calc_pout_13, calc_pout_12, calc_pout_11, calc_pout_10, calc_pout_9, calc_pout_8, calc_pout_7, calc_pout_6, calc_pout_5, calc_pout_4, calc_pout_3, calc_pout_2, calc_pout_1, calc_pout_0 } : abuf_wr_data_0;
  assign _0000_ = _0895_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12588" *) calc_addr_out : abuf_wr_addr;
  assign _0057_ = calc_dlv_valid_d4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11609" *) calc_layer_end_d4 : calc_layer_end_d5;
  assign _0450_ = calc_dlv_valid_d4 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11548" *) calc_stripe_end_d4 : calc_stripe_end_d5;
  assign _0049_ = _0894_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11487" *) calc_dlv_en_d4 : calc_dlv_en_d5;
  assign _0056_ = calc_dlv_valid_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11419" *) calc_layer_end_d3 : calc_layer_end_d4;
  assign _0449_ = calc_dlv_valid_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11358" *) calc_stripe_end_d3 : calc_stripe_end_d4;
  assign _0048_ = _0893_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11297" *) calc_dlv_en_d3 : calc_dlv_en_d4;
  assign _0055_ = calc_dlv_valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11229" *) calc_layer_end_d2 : calc_layer_end_d3;
  assign _0448_ = calc_dlv_valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11168" *) calc_stripe_end_d2 : calc_stripe_end_d3;
  assign _0047_ = _0892_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11107" *) calc_dlv_en_d2 : calc_dlv_en_d3;
  assign _0054_ = calc_dlv_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:11039" *) calc_layer_end_d1 : calc_layer_end_d2;
  assign _0447_ = calc_dlv_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10978" *) calc_stripe_end_d1 : calc_stripe_end_d2;
  assign _0046_ = _0891_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10917" *) calc_dlv_en_d1 : calc_dlv_en_d2;
  assign _0012_ = calc_valid_d3 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10843" *) calc_addr_d3 : calc_addr_d4;
  assign _0454_ = _0890_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10782" *) calc_wr_en_d3 : calc_wr_en_d4;
  assign _0011_ = calc_valid_d2 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10714" *) calc_addr_d2 : calc_addr_d3;
  assign _0453_ = _0889_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10653" *) calc_wr_en_d2 : calc_wr_en_d3;
  assign _0010_ = calc_valid_d1 ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10585" *) calc_addr_d1 : calc_addr_d2;
  assign _0452_ = _0888_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10524" *) calc_wr_en_d1 : calc_wr_en_d2;
  assign _0050_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7697" *) calc_dlv_elem_en[191:128] : calc_dlv_en_fp_d1;
  assign _0051_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7636" *) calc_dlv_elem_en[127:0] : calc_dlv_en_int_d1;
  assign _0442_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7575" *) calc_elem_op1_vld[191:128] : calc_op1_vld_fp_d1;
  assign _0443_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7514" *) calc_elem_op1_vld[127:0] : calc_op1_vld_int_d1;
  assign _0444_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7453" *) calc_elem_en[191:128] : calc_op_en_fp_d1;
  assign _0445_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7392" *) calc_elem_en[127:0] : calc_op_en_int_d1;
  assign _0053_ = accu_ctrl_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7331" *) accu_ctrl_pd[19] : calc_layer_end_d1;
  assign _0446_ = accu_ctrl_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7270" *) accu_ctrl_pd[17] : calc_stripe_end_d1;
  assign _0045_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7209" *) calc_dlv_en : calc_dlv_en_d1;
  assign _0009_ = accu_ctrl_valid ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7141" *) accu_ctrl_pd[4:0] : calc_addr_d1;
  assign _0451_ = _0897_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7080" *) calc_wr_en : calc_wr_en_d1;
  assign _0309_ = calc_elem_en[191] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7060" *) abuf_rd_data_3[767:720] : calc_op1_fp_63_d1;
  assign _0308_ = calc_elem_en[190] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7050" *) abuf_rd_data_3[719:672] : calc_op1_fp_62_d1;
  assign _0307_ = calc_elem_en[189] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7040" *) abuf_rd_data_3[671:624] : calc_op1_fp_61_d1;
  assign _0306_ = calc_elem_en[188] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7030" *) abuf_rd_data_3[623:576] : calc_op1_fp_60_d1;
  assign _0304_ = calc_elem_en[187] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7020" *) abuf_rd_data_3[575:528] : calc_op1_fp_59_d1;
  assign _0303_ = calc_elem_en[186] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7010" *) abuf_rd_data_3[527:480] : calc_op1_fp_58_d1;
  assign _0302_ = calc_elem_en[185] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7000" *) abuf_rd_data_3[479:432] : calc_op1_fp_57_d1;
  assign _0301_ = calc_elem_en[184] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6990" *) abuf_rd_data_3[431:384] : calc_op1_fp_56_d1;
  assign _0300_ = calc_elem_en[183] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6980" *) abuf_rd_data_3[383:336] : calc_op1_fp_55_d1;
  assign _0299_ = calc_elem_en[182] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6970" *) abuf_rd_data_3[335:288] : calc_op1_fp_54_d1;
  assign _0298_ = calc_elem_en[181] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6960" *) abuf_rd_data_3[287:240] : calc_op1_fp_53_d1;
  assign _0297_ = calc_elem_en[180] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6950" *) abuf_rd_data_3[239:192] : calc_op1_fp_52_d1;
  assign _0296_ = calc_elem_en[179] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6940" *) abuf_rd_data_3[191:144] : calc_op1_fp_51_d1;
  assign _0295_ = calc_elem_en[178] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6930" *) abuf_rd_data_3[143:96] : calc_op1_fp_50_d1;
  assign _0293_ = calc_elem_en[177] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6920" *) abuf_rd_data_3[95:48] : calc_op1_fp_49_d1;
  assign _0292_ = calc_elem_en[176] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6910" *) abuf_rd_data_3[47:0] : calc_op1_fp_48_d1;
  assign _0291_ = calc_elem_en[175] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6900" *) abuf_rd_data_2[767:720] : calc_op1_fp_47_d1;
  assign _0290_ = calc_elem_en[174] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6890" *) abuf_rd_data_2[719:672] : calc_op1_fp_46_d1;
  assign _0289_ = calc_elem_en[173] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6880" *) abuf_rd_data_2[671:624] : calc_op1_fp_45_d1;
  assign _0288_ = calc_elem_en[172] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6870" *) abuf_rd_data_2[623:576] : calc_op1_fp_44_d1;
  assign _0287_ = calc_elem_en[171] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6860" *) abuf_rd_data_2[575:528] : calc_op1_fp_43_d1;
  assign _0286_ = calc_elem_en[170] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6850" *) abuf_rd_data_2[527:480] : calc_op1_fp_42_d1;
  assign _0285_ = calc_elem_en[169] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6840" *) abuf_rd_data_2[479:432] : calc_op1_fp_41_d1;
  assign _0284_ = calc_elem_en[168] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6830" *) abuf_rd_data_2[431:384] : calc_op1_fp_40_d1;
  assign _0282_ = calc_elem_en[167] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6820" *) abuf_rd_data_2[383:336] : calc_op1_fp_39_d1;
  assign _0281_ = calc_elem_en[166] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6810" *) abuf_rd_data_2[335:288] : calc_op1_fp_38_d1;
  assign _0280_ = calc_elem_en[165] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6800" *) abuf_rd_data_2[287:240] : calc_op1_fp_37_d1;
  assign _0279_ = calc_elem_en[164] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6790" *) abuf_rd_data_2[239:192] : calc_op1_fp_36_d1;
  assign _0278_ = calc_elem_en[163] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6780" *) abuf_rd_data_2[191:144] : calc_op1_fp_35_d1;
  assign _0277_ = calc_elem_en[162] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6770" *) abuf_rd_data_2[143:96] : calc_op1_fp_34_d1;
  assign _0276_ = calc_elem_en[161] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6760" *) abuf_rd_data_2[95:48] : calc_op1_fp_33_d1;
  assign _0275_ = calc_elem_en[160] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6750" *) abuf_rd_data_2[47:0] : calc_op1_fp_32_d1;
  assign _0274_ = calc_elem_en[159] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6740" *) abuf_rd_data_1[767:720] : calc_op1_fp_31_d1;
  assign _0273_ = calc_elem_en[158] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6730" *) abuf_rd_data_1[719:672] : calc_op1_fp_30_d1;
  assign _0271_ = calc_elem_en[157] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6720" *) abuf_rd_data_1[671:624] : calc_op1_fp_29_d1;
  assign _0270_ = calc_elem_en[156] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6710" *) abuf_rd_data_1[623:576] : calc_op1_fp_28_d1;
  assign _0269_ = calc_elem_en[155] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6700" *) abuf_rd_data_1[575:528] : calc_op1_fp_27_d1;
  assign _0268_ = calc_elem_en[154] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6690" *) abuf_rd_data_1[527:480] : calc_op1_fp_26_d1;
  assign _0267_ = calc_elem_en[153] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6680" *) abuf_rd_data_1[479:432] : calc_op1_fp_25_d1;
  assign _0266_ = calc_elem_en[152] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6670" *) abuf_rd_data_1[431:384] : calc_op1_fp_24_d1;
  assign _0265_ = calc_elem_en[151] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6660" *) abuf_rd_data_1[383:336] : calc_op1_fp_23_d1;
  assign _0264_ = calc_elem_en[150] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6650" *) abuf_rd_data_1[335:288] : calc_op1_fp_22_d1;
  assign _0263_ = calc_elem_en[149] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6640" *) abuf_rd_data_1[287:240] : calc_op1_fp_21_d1;
  assign _0262_ = calc_elem_en[148] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6630" *) abuf_rd_data_1[239:192] : calc_op1_fp_20_d1;
  assign _0260_ = calc_elem_en[147] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6620" *) abuf_rd_data_1[191:144] : calc_op1_fp_19_d1;
  assign _0259_ = calc_elem_en[146] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6610" *) abuf_rd_data_1[143:96] : calc_op1_fp_18_d1;
  assign _0258_ = calc_elem_en[145] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6600" *) abuf_rd_data_1[95:48] : calc_op1_fp_17_d1;
  assign _0257_ = calc_elem_en[144] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6590" *) abuf_rd_data_1[47:0] : calc_op1_fp_16_d1;
  assign _0256_ = calc_elem_en[143] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6580" *) abuf_rd_data_0_sft[767:720] : calc_op1_fp_15_d1;
  assign _0255_ = calc_elem_en[142] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6570" *) abuf_rd_data_0_sft[719:672] : calc_op1_fp_14_d1;
  assign _0254_ = calc_elem_en[141] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6560" *) abuf_rd_data_0_sft[671:624] : calc_op1_fp_13_d1;
  assign _0253_ = calc_elem_en[140] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6550" *) abuf_rd_data_0_sft[623:576] : calc_op1_fp_12_d1;
  assign _0252_ = calc_elem_en[139] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6540" *) abuf_rd_data_0_sft[575:528] : calc_op1_fp_11_d1;
  assign _0251_ = calc_elem_en[138] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6530" *) abuf_rd_data_0_sft[527:480] : calc_op1_fp_10_d1;
  assign _0313_ = calc_elem_en[137] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6520" *) abuf_rd_data_0_sft[479:432] : calc_op1_fp_9_d1;
  assign _0312_ = calc_elem_en[136] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6510" *) abuf_rd_data_0_sft[431:384] : calc_op1_fp_8_d1;
  assign _0311_ = calc_elem_en[135] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6500" *) abuf_rd_data_0_sft[383:336] : calc_op1_fp_7_d1;
  assign _0310_ = calc_elem_en[134] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6490" *) abuf_rd_data_0_sft[335:288] : calc_op1_fp_6_d1;
  assign _0305_ = calc_elem_en[133] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6480" *) abuf_rd_data_0_sft[287:240] : calc_op1_fp_5_d1;
  assign _0294_ = calc_elem_en[132] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6470" *) abuf_rd_data_0_sft[239:192] : calc_op1_fp_4_d1;
  assign _0283_ = calc_elem_en[131] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6460" *) abuf_rd_data_0_sft[191:144] : calc_op1_fp_3_d1;
  assign _0272_ = calc_elem_en[130] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6450" *) abuf_rd_data_0_sft[143:96] : calc_op1_fp_2_d1;
  assign _0261_ = calc_elem_en[129] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6440" *) abuf_rd_data_0_sft[95:48] : calc_op1_fp_1_d1;
  assign _0250_ = calc_elem_en[128] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6430" *) abuf_rd_data_0_sft[47:0] : calc_op1_fp_0_d1;
  assign _0344_ = calc_elem_en[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6420" *) abuf_rd_data_7[543:510] : calc_op1_int_127_d1;
  assign _0343_ = calc_elem_en[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6410" *) abuf_rd_data_7[509:476] : calc_op1_int_126_d1;
  assign _0342_ = calc_elem_en[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6400" *) abuf_rd_data_7[475:442] : calc_op1_int_125_d1;
  assign _0341_ = calc_elem_en[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6390" *) abuf_rd_data_7[441:408] : calc_op1_int_124_d1;
  assign _0340_ = calc_elem_en[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6380" *) abuf_rd_data_7[407:374] : calc_op1_int_123_d1;
  assign _0339_ = calc_elem_en[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6370" *) abuf_rd_data_7[373:340] : calc_op1_int_122_d1;
  assign _0338_ = calc_elem_en[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6360" *) abuf_rd_data_7[339:306] : calc_op1_int_121_d1;
  assign _0337_ = calc_elem_en[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6350" *) abuf_rd_data_7[305:272] : calc_op1_int_120_d1;
  assign _0335_ = calc_elem_en[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6340" *) abuf_rd_data_7[271:238] : calc_op1_int_119_d1;
  assign _0334_ = calc_elem_en[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6330" *) abuf_rd_data_7[237:204] : calc_op1_int_118_d1;
  assign _0333_ = calc_elem_en[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6320" *) abuf_rd_data_7[203:170] : calc_op1_int_117_d1;
  assign _0332_ = calc_elem_en[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6310" *) abuf_rd_data_7[169:136] : calc_op1_int_116_d1;
  assign _0331_ = calc_elem_en[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6300" *) abuf_rd_data_7[135:102] : calc_op1_int_115_d1;
  assign _0330_ = calc_elem_en[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6290" *) abuf_rd_data_7[101:68] : calc_op1_int_114_d1;
  assign _0329_ = calc_elem_en[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6280" *) abuf_rd_data_7[67:34] : calc_op1_int_113_d1;
  assign _0328_ = calc_elem_en[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6270" *) abuf_rd_data_7[33:0] : calc_op1_int_112_d1;
  assign _0327_ = calc_elem_en[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6260" *) abuf_rd_data_6[543:510] : calc_op1_int_111_d1;
  assign _0326_ = calc_elem_en[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6250" *) abuf_rd_data_6[509:476] : calc_op1_int_110_d1;
  assign _0324_ = calc_elem_en[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6240" *) abuf_rd_data_6[475:442] : calc_op1_int_109_d1;
  assign _0323_ = calc_elem_en[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6230" *) abuf_rd_data_6[441:408] : calc_op1_int_108_d1;
  assign _0322_ = calc_elem_en[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6220" *) abuf_rd_data_6[407:374] : calc_op1_int_107_d1;
  assign _0321_ = calc_elem_en[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6210" *) abuf_rd_data_6[373:340] : calc_op1_int_106_d1;
  assign _0320_ = calc_elem_en[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6200" *) abuf_rd_data_6[339:306] : calc_op1_int_105_d1;
  assign _0319_ = calc_elem_en[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6190" *) abuf_rd_data_6[305:272] : calc_op1_int_104_d1;
  assign _0318_ = calc_elem_en[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6180" *) abuf_rd_data_6[271:238] : calc_op1_int_103_d1;
  assign _0317_ = calc_elem_en[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6170" *) abuf_rd_data_6[237:204] : calc_op1_int_102_d1;
  assign _0316_ = calc_elem_en[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6160" *) abuf_rd_data_6[203:170] : calc_op1_int_101_d1;
  assign _0315_ = calc_elem_en[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6150" *) abuf_rd_data_6[169:136] : calc_op1_int_100_d1;
  assign _0440_ = calc_elem_en[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6140" *) abuf_rd_data_6[135:102] : calc_op1_int_99_d1;
  assign _0439_ = calc_elem_en[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6130" *) abuf_rd_data_6[101:68] : calc_op1_int_98_d1;
  assign _0438_ = calc_elem_en[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6120" *) abuf_rd_data_6[67:34] : calc_op1_int_97_d1;
  assign _0437_ = calc_elem_en[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6110" *) abuf_rd_data_6[33:0] : calc_op1_int_96_d1;
  assign _0436_ = calc_elem_en[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6100" *) abuf_rd_data_5[543:510] : calc_op1_int_95_d1;
  assign _0435_ = calc_elem_en[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6090" *) abuf_rd_data_5[509:476] : calc_op1_int_94_d1;
  assign _0434_ = calc_elem_en[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6080" *) abuf_rd_data_5[475:442] : calc_op1_int_93_d1;
  assign _0433_ = calc_elem_en[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6070" *) abuf_rd_data_5[441:408] : calc_op1_int_92_d1;
  assign _0432_ = calc_elem_en[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6060" *) abuf_rd_data_5[407:374] : calc_op1_int_91_d1;
  assign _0431_ = calc_elem_en[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6050" *) abuf_rd_data_5[373:340] : calc_op1_int_90_d1;
  assign _0429_ = calc_elem_en[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6040" *) abuf_rd_data_5[339:306] : calc_op1_int_89_d1;
  assign _0428_ = calc_elem_en[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6030" *) abuf_rd_data_5[305:272] : calc_op1_int_88_d1;
  assign _0427_ = calc_elem_en[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6020" *) abuf_rd_data_5[271:238] : calc_op1_int_87_d1;
  assign _0426_ = calc_elem_en[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6010" *) abuf_rd_data_5[237:204] : calc_op1_int_86_d1;
  assign _0425_ = calc_elem_en[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:6000" *) abuf_rd_data_5[203:170] : calc_op1_int_85_d1;
  assign _0424_ = calc_elem_en[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5990" *) abuf_rd_data_5[169:136] : calc_op1_int_84_d1;
  assign _0423_ = calc_elem_en[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5980" *) abuf_rd_data_5[135:102] : calc_op1_int_83_d1;
  assign _0422_ = calc_elem_en[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5970" *) abuf_rd_data_5[101:68] : calc_op1_int_82_d1;
  assign _0421_ = calc_elem_en[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5960" *) abuf_rd_data_5[67:34] : calc_op1_int_81_d1;
  assign _0420_ = calc_elem_en[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5950" *) abuf_rd_data_5[33:0] : calc_op1_int_80_d1;
  assign _0418_ = calc_elem_en[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5940" *) abuf_rd_data_4_sft[543:510] : calc_op1_int_79_d1;
  assign _0417_ = calc_elem_en[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5930" *) abuf_rd_data_4_sft[509:476] : calc_op1_int_78_d1;
  assign _0416_ = calc_elem_en[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5920" *) abuf_rd_data_4_sft[475:442] : calc_op1_int_77_d1;
  assign _0415_ = calc_elem_en[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5910" *) abuf_rd_data_4_sft[441:408] : calc_op1_int_76_d1;
  assign _0414_ = calc_elem_en[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5900" *) abuf_rd_data_4_sft[407:374] : calc_op1_int_75_d1;
  assign _0413_ = calc_elem_en[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5890" *) abuf_rd_data_4_sft[373:340] : calc_op1_int_74_d1;
  assign _0412_ = calc_elem_en[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5880" *) abuf_rd_data_4_sft[339:306] : calc_op1_int_73_d1;
  assign _0411_ = calc_elem_en[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5870" *) abuf_rd_data_4_sft[305:272] : calc_op1_int_72_d1;
  assign _0410_ = calc_elem_en[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5860" *) abuf_rd_data_4_sft[271:238] : calc_op1_int_71_d1;
  assign _0409_ = calc_elem_en[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5850" *) abuf_rd_data_4_sft[237:204] : calc_op1_int_70_d1;
  assign _0407_ = calc_elem_en[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5840" *) abuf_rd_data_4_sft[203:170] : calc_op1_int_69_d1;
  assign _0406_ = calc_elem_en[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5830" *) abuf_rd_data_4_sft[169:136] : calc_op1_int_68_d1;
  assign _0405_ = calc_elem_en[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5820" *) abuf_rd_data_4_sft[135:102] : calc_op1_int_67_d1;
  assign _0404_ = calc_elem_en[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5810" *) abuf_rd_data_4_sft[101:68] : calc_op1_int_66_d1;
  assign _0403_ = calc_elem_en[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5800" *) abuf_rd_data_4_sft[67:34] : calc_op1_int_65_d1;
  assign _0402_ = calc_elem_en[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5790" *) abuf_rd_data_4_sft[33:0] : calc_op1_int_64_d1;
  assign _0401_ = calc_elem_en[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5780" *) abuf_rd_data_3[767:720] : calc_op1_int_63_d1;
  assign _0400_ = calc_elem_en[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5770" *) abuf_rd_data_3[719:672] : calc_op1_int_62_d1;
  assign _0399_ = calc_elem_en[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5760" *) abuf_rd_data_3[671:624] : calc_op1_int_61_d1;
  assign _0398_ = calc_elem_en[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5750" *) abuf_rd_data_3[623:576] : calc_op1_int_60_d1;
  assign _0396_ = calc_elem_en[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5740" *) abuf_rd_data_3[575:528] : calc_op1_int_59_d1;
  assign _0395_ = calc_elem_en[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5730" *) abuf_rd_data_3[527:480] : calc_op1_int_58_d1;
  assign _0394_ = calc_elem_en[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5720" *) abuf_rd_data_3[479:432] : calc_op1_int_57_d1;
  assign _0393_ = calc_elem_en[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5710" *) abuf_rd_data_3[431:384] : calc_op1_int_56_d1;
  assign _0392_ = calc_elem_en[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5700" *) abuf_rd_data_3[383:336] : calc_op1_int_55_d1;
  assign _0391_ = calc_elem_en[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5690" *) abuf_rd_data_3[335:288] : calc_op1_int_54_d1;
  assign _0390_ = calc_elem_en[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5680" *) abuf_rd_data_3[287:240] : calc_op1_int_53_d1;
  assign _0389_ = calc_elem_en[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5670" *) abuf_rd_data_3[239:192] : calc_op1_int_52_d1;
  assign _0388_ = calc_elem_en[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5660" *) abuf_rd_data_3[191:144] : calc_op1_int_51_d1;
  assign _0387_ = calc_elem_en[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5650" *) abuf_rd_data_3[143:96] : calc_op1_int_50_d1;
  assign _0385_ = calc_elem_en[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5640" *) abuf_rd_data_3[95:48] : calc_op1_int_49_d1;
  assign _0384_ = calc_elem_en[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5630" *) abuf_rd_data_3[47:0] : calc_op1_int_48_d1;
  assign _0383_ = calc_elem_en[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5620" *) abuf_rd_data_2[767:720] : calc_op1_int_47_d1;
  assign _0382_ = calc_elem_en[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5610" *) abuf_rd_data_2[719:672] : calc_op1_int_46_d1;
  assign _0381_ = calc_elem_en[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5600" *) abuf_rd_data_2[671:624] : calc_op1_int_45_d1;
  assign _0380_ = calc_elem_en[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5590" *) abuf_rd_data_2[623:576] : calc_op1_int_44_d1;
  assign _0379_ = calc_elem_en[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5580" *) abuf_rd_data_2[575:528] : calc_op1_int_43_d1;
  assign _0378_ = calc_elem_en[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5570" *) abuf_rd_data_2[527:480] : calc_op1_int_42_d1;
  assign _0377_ = calc_elem_en[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5560" *) abuf_rd_data_2[479:432] : calc_op1_int_41_d1;
  assign _0376_ = calc_elem_en[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5550" *) abuf_rd_data_2[431:384] : calc_op1_int_40_d1;
  assign _0374_ = calc_elem_en[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5540" *) abuf_rd_data_2[383:336] : calc_op1_int_39_d1;
  assign _0373_ = calc_elem_en[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5530" *) abuf_rd_data_2[335:288] : calc_op1_int_38_d1;
  assign _0372_ = calc_elem_en[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5520" *) abuf_rd_data_2[287:240] : calc_op1_int_37_d1;
  assign _0371_ = calc_elem_en[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5510" *) abuf_rd_data_2[239:192] : calc_op1_int_36_d1;
  assign _0370_ = calc_elem_en[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5500" *) abuf_rd_data_2[191:144] : calc_op1_int_35_d1;
  assign _0369_ = calc_elem_en[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5490" *) abuf_rd_data_2[143:96] : calc_op1_int_34_d1;
  assign _0368_ = calc_elem_en[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5480" *) abuf_rd_data_2[95:48] : calc_op1_int_33_d1;
  assign _0367_ = calc_elem_en[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5470" *) abuf_rd_data_2[47:0] : calc_op1_int_32_d1;
  assign _0366_ = calc_elem_en[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5460" *) abuf_rd_data_1[767:720] : calc_op1_int_31_d1;
  assign _0365_ = calc_elem_en[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5450" *) abuf_rd_data_1[719:672] : calc_op1_int_30_d1;
  assign _0363_ = calc_elem_en[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5440" *) abuf_rd_data_1[671:624] : calc_op1_int_29_d1;
  assign _0362_ = calc_elem_en[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5430" *) abuf_rd_data_1[623:576] : calc_op1_int_28_d1;
  assign _0361_ = calc_elem_en[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5420" *) abuf_rd_data_1[575:528] : calc_op1_int_27_d1;
  assign _0360_ = calc_elem_en[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5410" *) abuf_rd_data_1[527:480] : calc_op1_int_26_d1;
  assign _0359_ = calc_elem_en[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5400" *) abuf_rd_data_1[479:432] : calc_op1_int_25_d1;
  assign _0358_ = calc_elem_en[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5390" *) abuf_rd_data_1[431:384] : calc_op1_int_24_d1;
  assign _0357_ = calc_elem_en[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5380" *) abuf_rd_data_1[383:336] : calc_op1_int_23_d1;
  assign _0356_ = calc_elem_en[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5370" *) abuf_rd_data_1[335:288] : calc_op1_int_22_d1;
  assign _0355_ = calc_elem_en[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5360" *) abuf_rd_data_1[287:240] : calc_op1_int_21_d1;
  assign _0354_ = calc_elem_en[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5350" *) abuf_rd_data_1[239:192] : calc_op1_int_20_d1;
  assign _0352_ = calc_elem_en[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5340" *) abuf_rd_data_1[191:144] : calc_op1_int_19_d1;
  assign _0351_ = calc_elem_en[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5330" *) abuf_rd_data_1[143:96] : calc_op1_int_18_d1;
  assign _0350_ = calc_elem_en[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5320" *) abuf_rd_data_1[95:48] : calc_op1_int_17_d1;
  assign _0349_ = calc_elem_en[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5310" *) abuf_rd_data_1[47:0] : calc_op1_int_16_d1;
  assign _0348_ = calc_elem_en[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5300" *) abuf_rd_data_0_sft[767:720] : calc_op1_int_15_d1;
  assign _0347_ = calc_elem_en[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5290" *) abuf_rd_data_0_sft[719:672] : calc_op1_int_14_d1;
  assign _0346_ = calc_elem_en[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5280" *) abuf_rd_data_0_sft[671:624] : calc_op1_int_13_d1;
  assign _0345_ = calc_elem_en[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5270" *) abuf_rd_data_0_sft[623:576] : calc_op1_int_12_d1;
  assign _0336_ = calc_elem_en[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5260" *) abuf_rd_data_0_sft[575:528] : calc_op1_int_11_d1;
  assign _0325_ = calc_elem_en[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5250" *) abuf_rd_data_0_sft[527:480] : calc_op1_int_10_d1;
  assign _0441_ = calc_elem_en[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5240" *) abuf_rd_data_0_sft[479:432] : calc_op1_int_9_d1;
  assign _0430_ = calc_elem_en[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5230" *) abuf_rd_data_0_sft[431:384] : calc_op1_int_8_d1;
  assign _0419_ = calc_elem_en[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5220" *) abuf_rd_data_0_sft[383:336] : calc_op1_int_7_d1;
  assign _0408_ = calc_elem_en[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5210" *) abuf_rd_data_0_sft[335:288] : calc_op1_int_6_d1;
  assign _0397_ = calc_elem_en[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5200" *) abuf_rd_data_0_sft[287:240] : calc_op1_int_5_d1;
  assign _0386_ = calc_elem_en[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5190" *) abuf_rd_data_0_sft[239:192] : calc_op1_int_4_d1;
  assign _0375_ = calc_elem_en[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5180" *) abuf_rd_data_0_sft[191:144] : calc_op1_int_3_d1;
  assign _0364_ = calc_elem_en[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5170" *) abuf_rd_data_0_sft[143:96] : calc_op1_int_2_d1;
  assign _0353_ = calc_elem_en[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5160" *) abuf_rd_data_0_sft[95:48] : calc_op1_int_1_d1;
  assign _0314_ = calc_elem_en[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5150" *) abuf_rd_data_0_sft[47:0] : calc_op1_int_0_d1;
  assign _0117_ = calc_elem_en[191] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5140" *) calc_elem_63_w : calc_op0_fp_63_d1;
  assign _0116_ = calc_elem_en[190] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5130" *) calc_elem_62_w : calc_op0_fp_62_d1;
  assign _0115_ = calc_elem_en[189] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5120" *) calc_elem_61_w : calc_op0_fp_61_d1;
  assign _0114_ = calc_elem_en[188] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5110" *) calc_elem_60_w : calc_op0_fp_60_d1;
  assign _0112_ = calc_elem_en[187] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5100" *) calc_elem_59_w : calc_op0_fp_59_d1;
  assign _0111_ = calc_elem_en[186] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5090" *) calc_elem_58_w : calc_op0_fp_58_d1;
  assign _0110_ = calc_elem_en[185] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5080" *) calc_elem_57_w : calc_op0_fp_57_d1;
  assign _0109_ = calc_elem_en[184] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5070" *) calc_elem_56_w : calc_op0_fp_56_d1;
  assign _0108_ = calc_elem_en[183] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5060" *) calc_elem_55_w : calc_op0_fp_55_d1;
  assign _0107_ = calc_elem_en[182] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5050" *) calc_elem_54_w : calc_op0_fp_54_d1;
  assign _0106_ = calc_elem_en[181] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5040" *) calc_elem_53_w : calc_op0_fp_53_d1;
  assign _0105_ = calc_elem_en[180] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5030" *) calc_elem_52_w : calc_op0_fp_52_d1;
  assign _0104_ = calc_elem_en[179] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5020" *) calc_elem_51_w : calc_op0_fp_51_d1;
  assign _0103_ = calc_elem_en[178] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5010" *) calc_elem_50_w : calc_op0_fp_50_d1;
  assign _0101_ = calc_elem_en[177] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:5000" *) calc_elem_49_w : calc_op0_fp_49_d1;
  assign _0100_ = calc_elem_en[176] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4990" *) calc_elem_48_w : calc_op0_fp_48_d1;
  assign _0099_ = calc_elem_en[175] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4980" *) calc_elem_47_w : calc_op0_fp_47_d1;
  assign _0098_ = calc_elem_en[174] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4970" *) calc_elem_46_w : calc_op0_fp_46_d1;
  assign _0097_ = calc_elem_en[173] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4960" *) calc_elem_45_w : calc_op0_fp_45_d1;
  assign _0096_ = calc_elem_en[172] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4950" *) calc_elem_44_w : calc_op0_fp_44_d1;
  assign _0095_ = calc_elem_en[171] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4940" *) calc_elem_43_w : calc_op0_fp_43_d1;
  assign _0094_ = calc_elem_en[170] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4930" *) calc_elem_42_w : calc_op0_fp_42_d1;
  assign _0093_ = calc_elem_en[169] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4920" *) calc_elem_41_w : calc_op0_fp_41_d1;
  assign _0092_ = calc_elem_en[168] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4910" *) calc_elem_40_w : calc_op0_fp_40_d1;
  assign _0090_ = calc_elem_en[167] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4900" *) calc_elem_39_w : calc_op0_fp_39_d1;
  assign _0089_ = calc_elem_en[166] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4890" *) calc_elem_38_w : calc_op0_fp_38_d1;
  assign _0088_ = calc_elem_en[165] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4880" *) calc_elem_37_w : calc_op0_fp_37_d1;
  assign _0087_ = calc_elem_en[164] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4870" *) calc_elem_36_w : calc_op0_fp_36_d1;
  assign _0086_ = calc_elem_en[163] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4860" *) calc_elem_35_w : calc_op0_fp_35_d1;
  assign _0085_ = calc_elem_en[162] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4850" *) calc_elem_34_w : calc_op0_fp_34_d1;
  assign _0084_ = calc_elem_en[161] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4840" *) calc_elem_33_w : calc_op0_fp_33_d1;
  assign _0083_ = calc_elem_en[160] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4830" *) calc_elem_32_w : calc_op0_fp_32_d1;
  assign _0082_ = calc_elem_en[159] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4820" *) calc_elem_31_w : calc_op0_fp_31_d1;
  assign _0081_ = calc_elem_en[158] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4810" *) calc_elem_30_w : calc_op0_fp_30_d1;
  assign _0079_ = calc_elem_en[157] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4800" *) calc_elem_29_w : calc_op0_fp_29_d1;
  assign _0078_ = calc_elem_en[156] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4790" *) calc_elem_28_w : calc_op0_fp_28_d1;
  assign _0077_ = calc_elem_en[155] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4780" *) calc_elem_27_w : calc_op0_fp_27_d1;
  assign _0076_ = calc_elem_en[154] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4770" *) calc_elem_26_w : calc_op0_fp_26_d1;
  assign _0075_ = calc_elem_en[153] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4760" *) calc_elem_25_w : calc_op0_fp_25_d1;
  assign _0074_ = calc_elem_en[152] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4750" *) calc_elem_24_w : calc_op0_fp_24_d1;
  assign _0073_ = calc_elem_en[151] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4740" *) calc_elem_23_w : calc_op0_fp_23_d1;
  assign _0072_ = calc_elem_en[150] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4730" *) calc_elem_22_w : calc_op0_fp_22_d1;
  assign _0071_ = calc_elem_en[149] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4720" *) calc_elem_21_w : calc_op0_fp_21_d1;
  assign _0070_ = calc_elem_en[148] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4710" *) calc_elem_20_w : calc_op0_fp_20_d1;
  assign _0068_ = calc_elem_en[147] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4700" *) calc_elem_19_w : calc_op0_fp_19_d1;
  assign _0067_ = calc_elem_en[146] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4690" *) calc_elem_18_w : calc_op0_fp_18_d1;
  assign _0066_ = calc_elem_en[145] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4680" *) calc_elem_17_w : calc_op0_fp_17_d1;
  assign _0065_ = calc_elem_en[144] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4670" *) calc_elem_16_w : calc_op0_fp_16_d1;
  assign _0064_ = calc_elem_en[143] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4660" *) calc_elem_15_w : calc_op0_fp_15_d1;
  assign _0063_ = calc_elem_en[142] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4650" *) calc_elem_14_w : calc_op0_fp_14_d1;
  assign _0062_ = calc_elem_en[141] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4640" *) calc_elem_13_w : calc_op0_fp_13_d1;
  assign _0061_ = calc_elem_en[140] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4630" *) calc_elem_12_w : calc_op0_fp_12_d1;
  assign _0060_ = calc_elem_en[139] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4620" *) calc_elem_11_w : calc_op0_fp_11_d1;
  assign _0059_ = calc_elem_en[138] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4610" *) calc_elem_10_w : calc_op0_fp_10_d1;
  assign _0121_ = calc_elem_en[137] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4600" *) calc_elem_9_w : calc_op0_fp_9_d1;
  assign _0120_ = calc_elem_en[136] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4590" *) calc_elem_8_w : calc_op0_fp_8_d1;
  assign _0119_ = calc_elem_en[135] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4580" *) calc_elem_7_w : calc_op0_fp_7_d1;
  assign _0118_ = calc_elem_en[134] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4570" *) calc_elem_6_w : calc_op0_fp_6_d1;
  assign _0113_ = calc_elem_en[133] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4560" *) calc_elem_5_w : calc_op0_fp_5_d1;
  assign _0102_ = calc_elem_en[132] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4550" *) calc_elem_4_w : calc_op0_fp_4_d1;
  assign _0091_ = calc_elem_en[131] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4540" *) calc_elem_3_w : calc_op0_fp_3_d1;
  assign _0080_ = calc_elem_en[130] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4530" *) calc_elem_2_w : calc_op0_fp_2_d1;
  assign _0069_ = calc_elem_en[129] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4520" *) calc_elem_1_w : calc_op0_fp_1_d1;
  assign _0058_ = calc_elem_en[128] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4510" *) calc_elem_0_w : calc_op0_fp_0_d1;
  assign _0152_ = calc_elem_en[127] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4500" *) calc_data_15[175:154] : calc_op0_int_127_d1;
  assign _0151_ = calc_elem_en[126] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4490" *) calc_data_14[175:154] : calc_op0_int_126_d1;
  assign _0150_ = calc_elem_en[125] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4480" *) calc_data_13[175:154] : calc_op0_int_125_d1;
  assign _0149_ = calc_elem_en[124] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4470" *) calc_data_12[175:154] : calc_op0_int_124_d1;
  assign _0148_ = calc_elem_en[123] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4460" *) calc_data_11[175:154] : calc_op0_int_123_d1;
  assign _0147_ = calc_elem_en[122] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4450" *) calc_data_10[175:154] : calc_op0_int_122_d1;
  assign _0146_ = calc_elem_en[121] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4440" *) calc_data_9[175:154] : calc_op0_int_121_d1;
  assign _0145_ = calc_elem_en[120] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4430" *) calc_data_8[175:154] : calc_op0_int_120_d1;
  assign _0143_ = calc_elem_en[119] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4420" *) calc_data_7[175:154] : calc_op0_int_119_d1;
  assign _0142_ = calc_elem_en[118] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4410" *) calc_data_6[175:154] : calc_op0_int_118_d1;
  assign _0141_ = calc_elem_en[117] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4400" *) calc_data_5[175:154] : calc_op0_int_117_d1;
  assign _0140_ = calc_elem_en[116] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4390" *) calc_data_4[175:154] : calc_op0_int_116_d1;
  assign _0139_ = calc_elem_en[115] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4380" *) calc_data_3[175:154] : calc_op0_int_115_d1;
  assign _0138_ = calc_elem_en[114] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4370" *) calc_data_2[175:154] : calc_op0_int_114_d1;
  assign _0137_ = calc_elem_en[113] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4360" *) calc_data_1[175:154] : calc_op0_int_113_d1;
  assign _0136_ = calc_elem_en[112] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4350" *) calc_data_0[175:154] : calc_op0_int_112_d1;
  assign _0135_ = calc_elem_en[111] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4340" *) calc_data_15[131:110] : calc_op0_int_111_d1;
  assign _0134_ = calc_elem_en[110] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4330" *) calc_data_14[131:110] : calc_op0_int_110_d1;
  assign _0132_ = calc_elem_en[109] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4320" *) calc_data_13[131:110] : calc_op0_int_109_d1;
  assign _0131_ = calc_elem_en[108] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4310" *) calc_data_12[131:110] : calc_op0_int_108_d1;
  assign _0130_ = calc_elem_en[107] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4300" *) calc_data_11[131:110] : calc_op0_int_107_d1;
  assign _0129_ = calc_elem_en[106] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4290" *) calc_data_10[131:110] : calc_op0_int_106_d1;
  assign _0128_ = calc_elem_en[105] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4280" *) calc_data_9[131:110] : calc_op0_int_105_d1;
  assign _0127_ = calc_elem_en[104] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4270" *) calc_data_8[131:110] : calc_op0_int_104_d1;
  assign _0126_ = calc_elem_en[103] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4260" *) calc_data_7[131:110] : calc_op0_int_103_d1;
  assign _0125_ = calc_elem_en[102] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4250" *) calc_data_6[131:110] : calc_op0_int_102_d1;
  assign _0124_ = calc_elem_en[101] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4240" *) calc_data_5[131:110] : calc_op0_int_101_d1;
  assign _0123_ = calc_elem_en[100] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4230" *) calc_data_4[131:110] : calc_op0_int_100_d1;
  assign _0248_ = calc_elem_en[99] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4220" *) calc_data_3[131:110] : calc_op0_int_99_d1;
  assign _0247_ = calc_elem_en[98] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4210" *) calc_data_2[131:110] : calc_op0_int_98_d1;
  assign _0246_ = calc_elem_en[97] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4200" *) calc_data_1[131:110] : calc_op0_int_97_d1;
  assign _0245_ = calc_elem_en[96] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4190" *) calc_data_0[131:110] : calc_op0_int_96_d1;
  assign _0244_ = calc_elem_en[95] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4180" *) calc_data_15[87:66] : calc_op0_int_95_d1;
  assign _0243_ = calc_elem_en[94] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4170" *) calc_data_14[87:66] : calc_op0_int_94_d1;
  assign _0242_ = calc_elem_en[93] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4160" *) calc_data_13[87:66] : calc_op0_int_93_d1;
  assign _0241_ = calc_elem_en[92] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4150" *) calc_data_12[87:66] : calc_op0_int_92_d1;
  assign _0240_ = calc_elem_en[91] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4140" *) calc_data_11[87:66] : calc_op0_int_91_d1;
  assign _0239_ = calc_elem_en[90] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4130" *) calc_data_10[87:66] : calc_op0_int_90_d1;
  assign _0237_ = calc_elem_en[89] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4120" *) calc_data_9[87:66] : calc_op0_int_89_d1;
  assign _0236_ = calc_elem_en[88] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4110" *) calc_data_8[87:66] : calc_op0_int_88_d1;
  assign _0235_ = calc_elem_en[87] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4100" *) calc_data_7[87:66] : calc_op0_int_87_d1;
  assign _0234_ = calc_elem_en[86] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4090" *) calc_data_6[87:66] : calc_op0_int_86_d1;
  assign _0233_ = calc_elem_en[85] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4080" *) calc_data_5[87:66] : calc_op0_int_85_d1;
  assign _0232_ = calc_elem_en[84] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4070" *) calc_data_4[87:66] : calc_op0_int_84_d1;
  assign _0231_ = calc_elem_en[83] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4060" *) calc_data_3[87:66] : calc_op0_int_83_d1;
  assign _0230_ = calc_elem_en[82] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4050" *) calc_data_2[87:66] : calc_op0_int_82_d1;
  assign _0229_ = calc_elem_en[81] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4040" *) calc_data_1[87:66] : calc_op0_int_81_d1;
  assign _0228_ = calc_elem_en[80] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4030" *) calc_data_0[87:66] : calc_op0_int_80_d1;
  assign _0226_ = calc_elem_en[79] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4020" *) calc_data_15[43:22] : calc_op0_int_79_d1;
  assign _0225_ = calc_elem_en[78] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4010" *) calc_data_14[43:22] : calc_op0_int_78_d1;
  assign _0224_ = calc_elem_en[77] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:4000" *) calc_data_13[43:22] : calc_op0_int_77_d1;
  assign _0223_ = calc_elem_en[76] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3990" *) calc_data_12[43:22] : calc_op0_int_76_d1;
  assign _0222_ = calc_elem_en[75] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3980" *) calc_data_11[43:22] : calc_op0_int_75_d1;
  assign _0221_ = calc_elem_en[74] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3970" *) calc_data_10[43:22] : calc_op0_int_74_d1;
  assign _0220_ = calc_elem_en[73] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3960" *) calc_data_9[43:22] : calc_op0_int_73_d1;
  assign _0219_ = calc_elem_en[72] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3950" *) calc_data_8[43:22] : calc_op0_int_72_d1;
  assign _0218_ = calc_elem_en[71] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3940" *) calc_data_7[43:22] : calc_op0_int_71_d1;
  assign _0217_ = calc_elem_en[70] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3930" *) calc_data_6[43:22] : calc_op0_int_70_d1;
  assign _0215_ = calc_elem_en[69] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3920" *) calc_data_5[43:22] : calc_op0_int_69_d1;
  assign _0214_ = calc_elem_en[68] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3910" *) calc_data_4[43:22] : calc_op0_int_68_d1;
  assign _0213_ = calc_elem_en[67] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3900" *) calc_data_3[43:22] : calc_op0_int_67_d1;
  assign _0212_ = calc_elem_en[66] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3890" *) calc_data_2[43:22] : calc_op0_int_66_d1;
  assign _0211_ = calc_elem_en[65] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3880" *) calc_data_1[43:22] : calc_op0_int_65_d1;
  assign _0210_ = calc_elem_en[64] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3870" *) calc_data_0[43:22] : calc_op0_int_64_d1;
  assign _0209_ = calc_elem_en[63] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3860" *) calc_elem_63_w[37:0] : calc_op0_int_63_d1;
  assign _0208_ = calc_elem_en[62] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3850" *) calc_elem_62_w[37:0] : calc_op0_int_62_d1;
  assign _0207_ = calc_elem_en[61] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3840" *) calc_elem_61_w[37:0] : calc_op0_int_61_d1;
  assign _0206_ = calc_elem_en[60] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3830" *) calc_elem_60_w[37:0] : calc_op0_int_60_d1;
  assign _0204_ = calc_elem_en[59] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3820" *) calc_elem_59_w[37:0] : calc_op0_int_59_d1;
  assign _0203_ = calc_elem_en[58] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3810" *) calc_elem_58_w[37:0] : calc_op0_int_58_d1;
  assign _0202_ = calc_elem_en[57] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3800" *) calc_elem_57_w[37:0] : calc_op0_int_57_d1;
  assign _0201_ = calc_elem_en[56] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3790" *) calc_elem_56_w[37:0] : calc_op0_int_56_d1;
  assign _0200_ = calc_elem_en[55] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3780" *) calc_elem_55_w[37:0] : calc_op0_int_55_d1;
  assign _0199_ = calc_elem_en[54] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3770" *) calc_elem_54_w[37:0] : calc_op0_int_54_d1;
  assign _0198_ = calc_elem_en[53] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3760" *) calc_elem_53_w[37:0] : calc_op0_int_53_d1;
  assign _0197_ = calc_elem_en[52] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3750" *) calc_elem_52_w[37:0] : calc_op0_int_52_d1;
  assign _0196_ = calc_elem_en[51] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3740" *) calc_elem_51_w[37:0] : calc_op0_int_51_d1;
  assign _0195_ = calc_elem_en[50] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3730" *) calc_elem_50_w[37:0] : calc_op0_int_50_d1;
  assign _0193_ = calc_elem_en[49] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3720" *) calc_elem_49_w[37:0] : calc_op0_int_49_d1;
  assign _0192_ = calc_elem_en[48] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3710" *) calc_elem_48_w[37:0] : calc_op0_int_48_d1;
  assign _0191_ = calc_elem_en[47] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3700" *) calc_elem_47_w[37:0] : calc_op0_int_47_d1;
  assign _0190_ = calc_elem_en[46] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3690" *) calc_elem_46_w[37:0] : calc_op0_int_46_d1;
  assign _0189_ = calc_elem_en[45] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3680" *) calc_elem_45_w[37:0] : calc_op0_int_45_d1;
  assign _0188_ = calc_elem_en[44] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3670" *) calc_elem_44_w[37:0] : calc_op0_int_44_d1;
  assign _0187_ = calc_elem_en[43] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3660" *) calc_elem_43_w[37:0] : calc_op0_int_43_d1;
  assign _0186_ = calc_elem_en[42] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3650" *) calc_elem_42_w[37:0] : calc_op0_int_42_d1;
  assign _0185_ = calc_elem_en[41] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3640" *) calc_elem_41_w[37:0] : calc_op0_int_41_d1;
  assign _0184_ = calc_elem_en[40] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3630" *) calc_elem_40_w[37:0] : calc_op0_int_40_d1;
  assign _0182_ = calc_elem_en[39] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3620" *) calc_elem_39_w[37:0] : calc_op0_int_39_d1;
  assign _0181_ = calc_elem_en[38] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3610" *) calc_elem_38_w[37:0] : calc_op0_int_38_d1;
  assign _0180_ = calc_elem_en[37] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3600" *) calc_elem_37_w[37:0] : calc_op0_int_37_d1;
  assign _0179_ = calc_elem_en[36] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3590" *) calc_elem_36_w[37:0] : calc_op0_int_36_d1;
  assign _0178_ = calc_elem_en[35] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3580" *) calc_elem_35_w[37:0] : calc_op0_int_35_d1;
  assign _0177_ = calc_elem_en[34] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3570" *) calc_elem_34_w[37:0] : calc_op0_int_34_d1;
  assign _0176_ = calc_elem_en[33] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3560" *) calc_elem_33_w[37:0] : calc_op0_int_33_d1;
  assign _0175_ = calc_elem_en[32] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3550" *) calc_elem_32_w[37:0] : calc_op0_int_32_d1;
  assign _0174_ = calc_elem_en[31] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3540" *) calc_elem_31_w[37:0] : calc_op0_int_31_d1;
  assign _0173_ = calc_elem_en[30] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3530" *) calc_elem_30_w[37:0] : calc_op0_int_30_d1;
  assign _0171_ = calc_elem_en[29] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3520" *) calc_elem_29_w[37:0] : calc_op0_int_29_d1;
  assign _0170_ = calc_elem_en[28] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3510" *) calc_elem_28_w[37:0] : calc_op0_int_28_d1;
  assign _0169_ = calc_elem_en[27] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3500" *) calc_elem_27_w[37:0] : calc_op0_int_27_d1;
  assign _0168_ = calc_elem_en[26] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3490" *) calc_elem_26_w[37:0] : calc_op0_int_26_d1;
  assign _0167_ = calc_elem_en[25] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3480" *) calc_elem_25_w[37:0] : calc_op0_int_25_d1;
  assign _0166_ = calc_elem_en[24] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3470" *) calc_elem_24_w[37:0] : calc_op0_int_24_d1;
  assign _0165_ = calc_elem_en[23] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3460" *) calc_elem_23_w[37:0] : calc_op0_int_23_d1;
  assign _0164_ = calc_elem_en[22] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3450" *) calc_elem_22_w[37:0] : calc_op0_int_22_d1;
  assign _0163_ = calc_elem_en[21] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3440" *) calc_elem_21_w[37:0] : calc_op0_int_21_d1;
  assign _0162_ = calc_elem_en[20] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3430" *) calc_elem_20_w[37:0] : calc_op0_int_20_d1;
  assign _0160_ = calc_elem_en[19] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3420" *) calc_elem_19_w[37:0] : calc_op0_int_19_d1;
  assign _0159_ = calc_elem_en[18] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3410" *) calc_elem_18_w[37:0] : calc_op0_int_18_d1;
  assign _0158_ = calc_elem_en[17] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3400" *) calc_elem_17_w[37:0] : calc_op0_int_17_d1;
  assign _0157_ = calc_elem_en[16] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3390" *) calc_elem_16_w[37:0] : calc_op0_int_16_d1;
  assign _0156_ = calc_elem_en[15] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3380" *) calc_elem_15_w[37:0] : calc_op0_int_15_d1;
  assign _0155_ = calc_elem_en[14] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3370" *) calc_elem_14_w[37:0] : calc_op0_int_14_d1;
  assign _0154_ = calc_elem_en[13] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3360" *) calc_elem_13_w[37:0] : calc_op0_int_13_d1;
  assign _0153_ = calc_elem_en[12] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3350" *) calc_elem_12_w[37:0] : calc_op0_int_12_d1;
  assign _0144_ = calc_elem_en[11] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3340" *) calc_elem_11_w[37:0] : calc_op0_int_11_d1;
  assign _0133_ = calc_elem_en[10] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3330" *) calc_elem_10_w[37:0] : calc_op0_int_10_d1;
  assign _0249_ = calc_elem_en[9] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3320" *) calc_elem_9_w[37:0] : calc_op0_int_9_d1;
  assign _0238_ = calc_elem_en[8] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3310" *) calc_elem_8_w[37:0] : calc_op0_int_8_d1;
  assign _0227_ = calc_elem_en[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3300" *) calc_elem_7_w[37:0] : calc_op0_int_7_d1;
  assign _0216_ = calc_elem_en[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3290" *) calc_elem_6_w[37:0] : calc_op0_int_6_d1;
  assign _0205_ = calc_elem_en[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3280" *) calc_elem_5_w[37:0] : calc_op0_int_5_d1;
  assign _0194_ = calc_elem_en[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3270" *) calc_elem_4_w[37:0] : calc_op0_int_4_d1;
  assign _0183_ = calc_elem_en[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3260" *) calc_elem_3_w[37:0] : calc_op0_int_3_d1;
  assign _0172_ = calc_elem_en[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3250" *) calc_elem_2_w[37:0] : calc_op0_int_2_d1;
  assign _0161_ = calc_elem_en[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3240" *) calc_elem_1_w[37:0] : calc_op0_int_1_d1;
  assign _0122_ = calc_elem_en[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3230" *) calc_elem_0_w[37:0] : calc_op0_int_0_d1;
  assign _0052_ = _0896_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2616" *) { mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask, mac_b2accu_mask, mac_a2accu_mask } : calc_in_mask;
  assign _0025_ = _0879_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2580" *) mac_b2accu_data7[175:44] : calc_data_15[175:44];
  assign _0026_ = mac_b2accu_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2570" *) mac_b2accu_data7[43:0] : calc_data_15[43:0];
  assign _0023_ = _0878_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2560" *) mac_b2accu_data6[175:44] : calc_data_14[175:44];
  assign _0024_ = mac_b2accu_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2550" *) mac_b2accu_data6[43:0] : calc_data_14[43:0];
  assign _0021_ = _0877_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2540" *) mac_b2accu_data5[175:44] : calc_data_13[175:44];
  assign _0022_ = mac_b2accu_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2530" *) mac_b2accu_data5[43:0] : calc_data_13[43:0];
  assign _0019_ = _0876_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2520" *) mac_b2accu_data4[175:44] : calc_data_12[175:44];
  assign _0020_ = mac_b2accu_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2510" *) mac_b2accu_data4[43:0] : calc_data_12[43:0];
  assign _0017_ = _0875_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2500" *) mac_b2accu_data3[175:44] : calc_data_11[175:44];
  assign _0018_ = mac_b2accu_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2490" *) mac_b2accu_data3[43:0] : calc_data_11[43:0];
  assign _0015_ = _0874_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2480" *) mac_b2accu_data2[175:44] : calc_data_10[175:44];
  assign _0016_ = mac_b2accu_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2470" *) mac_b2accu_data2[43:0] : calc_data_10[43:0];
  assign _0043_ = _0873_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2460" *) mac_b2accu_data1[175:44] : calc_data_9[175:44];
  assign _0044_ = mac_b2accu_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2450" *) mac_b2accu_data1[43:0] : calc_data_9[43:0];
  assign _0041_ = _0872_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2440" *) mac_b2accu_data0[175:44] : calc_data_8[175:44];
  assign _0042_ = mac_b2accu_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2430" *) mac_b2accu_data0[43:0] : calc_data_8[43:0];
  assign _0039_ = _0871_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2420" *) mac_a2accu_data7[175:44] : calc_data_7[175:44];
  assign _0040_ = mac_a2accu_mask[7] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2410" *) mac_a2accu_data7[43:0] : calc_data_7[43:0];
  assign _0037_ = _0870_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2400" *) mac_a2accu_data6[175:44] : calc_data_6[175:44];
  assign _0038_ = mac_a2accu_mask[6] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2390" *) mac_a2accu_data6[43:0] : calc_data_6[43:0];
  assign _0035_ = _0869_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2380" *) mac_a2accu_data5[175:44] : calc_data_5[175:44];
  assign _0036_ = mac_a2accu_mask[5] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2370" *) mac_a2accu_data5[43:0] : calc_data_5[43:0];
  assign _0033_ = _0868_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2360" *) mac_a2accu_data4[175:44] : calc_data_4[175:44];
  assign _0034_ = mac_a2accu_mask[4] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2350" *) mac_a2accu_data4[43:0] : calc_data_4[43:0];
  assign _0031_ = _0867_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2340" *) mac_a2accu_data3[175:44] : calc_data_3[175:44];
  assign _0032_ = mac_a2accu_mask[3] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2330" *) mac_a2accu_data3[43:0] : calc_data_3[43:0];
  assign _0029_ = _0866_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2320" *) mac_a2accu_data2[175:44] : calc_data_2[175:44];
  assign _0030_ = mac_a2accu_mask[2] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2310" *) mac_a2accu_data2[43:0] : calc_data_2[43:0];
  assign _0027_ = _0865_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2300" *) mac_a2accu_data1[175:44] : calc_data_1[175:44];
  assign _0028_ = mac_a2accu_mask[1] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2290" *) mac_a2accu_data1[43:0] : calc_data_1[43:0];
  assign _0013_ = _0864_ ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2280" *) mac_a2accu_data0[175:44] : calc_data_0[175:44];
  assign _0014_ = mac_a2accu_mask[0] ? (* full_case = 32'd1 *) (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2270" *) mac_a2accu_data0[43:0] : calc_data_0[43:0];
  assign _0895_ = | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12588" *) { calc_wr_en_out[0], calc_wr_en_out[1], calc_wr_en_out[2], calc_wr_en_out[3], calc_wr_en_out[4], calc_wr_en_out[5], calc_wr_en_out[6], calc_wr_en_out[7] };
  assign _0909_ = | (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13420" *) { sat_sum[0], sat_sum[1], sat_sum[2], sat_sum[3], sat_sum[4], sat_sum[5], sat_sum[6], sat_sum[7] };
  assign abuf_wr_elem_16 = cfg_is_wg[0] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12332" *) calc_pout_16 : calc_pout_0;
  assign abuf_wr_elem_17 = cfg_is_wg[1] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12333" *) calc_pout_17 : calc_pout_1;
  assign abuf_wr_elem_18 = cfg_is_wg[2] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12334" *) calc_pout_18 : calc_pout_2;
  assign abuf_wr_elem_19 = cfg_is_wg[3] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12335" *) calc_pout_19 : calc_pout_3;
  assign abuf_wr_elem_20 = cfg_is_wg[4] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12336" *) calc_pout_20 : calc_pout_4;
  assign abuf_wr_elem_21 = cfg_is_wg[5] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12337" *) calc_pout_21 : calc_pout_5;
  assign abuf_wr_elem_22 = cfg_is_wg[6] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12338" *) calc_pout_22 : calc_pout_6;
  assign abuf_wr_elem_23 = cfg_is_wg[7] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12339" *) calc_pout_23 : calc_pout_7;
  assign abuf_wr_elem_24 = cfg_is_wg[8] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12340" *) calc_pout_24 : calc_pout_8;
  assign abuf_wr_elem_25 = cfg_is_wg[9] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12341" *) calc_pout_25 : calc_pout_9;
  assign abuf_wr_elem_26 = cfg_is_wg[10] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12342" *) calc_pout_26 : calc_pout_10;
  assign abuf_wr_elem_27 = cfg_is_wg[11] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12343" *) calc_pout_27 : calc_pout_11;
  assign abuf_wr_elem_28 = cfg_is_wg[12] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12344" *) calc_pout_28 : calc_pout_12;
  assign abuf_wr_elem_29 = cfg_is_wg[13] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12345" *) calc_pout_29 : calc_pout_13;
  assign abuf_wr_elem_30 = cfg_is_wg[14] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12346" *) calc_pout_30 : calc_pout_14;
  assign abuf_wr_elem_31 = cfg_is_wg[15] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12347" *) calc_pout_31 : calc_pout_15;
  assign abuf_wr_elem_32 = cfg_is_wg[16] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12348" *) calc_pout_32 : calc_pout_0;
  assign abuf_wr_elem_33 = cfg_is_wg[17] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12349" *) calc_pout_33 : calc_pout_1;
  assign abuf_wr_elem_34 = cfg_is_wg[18] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12350" *) calc_pout_34 : calc_pout_2;
  assign abuf_wr_elem_35 = cfg_is_wg[19] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12351" *) calc_pout_35 : calc_pout_3;
  assign abuf_wr_elem_36 = cfg_is_wg[20] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12352" *) calc_pout_36 : calc_pout_4;
  assign abuf_wr_elem_37 = cfg_is_wg[21] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12353" *) calc_pout_37 : calc_pout_5;
  assign abuf_wr_elem_38 = cfg_is_wg[22] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12354" *) calc_pout_38 : calc_pout_6;
  assign abuf_wr_elem_39 = cfg_is_wg[23] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12355" *) calc_pout_39 : calc_pout_7;
  assign abuf_wr_elem_40 = cfg_is_wg[24] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12356" *) calc_pout_40 : calc_pout_8;
  assign abuf_wr_elem_41 = cfg_is_wg[25] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12357" *) calc_pout_41 : calc_pout_9;
  assign abuf_wr_elem_42 = cfg_is_wg[26] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12358" *) calc_pout_42 : calc_pout_10;
  assign abuf_wr_elem_43 = cfg_is_wg[27] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12359" *) calc_pout_43 : calc_pout_11;
  assign abuf_wr_elem_44 = cfg_is_wg[28] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12360" *) calc_pout_44 : calc_pout_12;
  assign abuf_wr_elem_45 = cfg_is_wg[29] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12361" *) calc_pout_45 : calc_pout_13;
  assign abuf_wr_elem_46 = cfg_is_wg[30] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12362" *) calc_pout_46 : calc_pout_14;
  assign abuf_wr_elem_47 = cfg_is_wg[31] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12363" *) calc_pout_47 : calc_pout_15;
  assign abuf_wr_elem_48 = cfg_is_wg[32] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12364" *) calc_pout_48 : calc_pout_0;
  assign abuf_wr_elem_49 = cfg_is_wg[33] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12365" *) calc_pout_49 : calc_pout_1;
  assign abuf_wr_elem_50 = cfg_is_wg[34] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12366" *) calc_pout_50 : calc_pout_2;
  assign abuf_wr_elem_51 = cfg_is_wg[35] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12367" *) calc_pout_51 : calc_pout_3;
  assign abuf_wr_elem_52 = cfg_is_wg[36] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12368" *) calc_pout_52 : calc_pout_4;
  assign abuf_wr_elem_53 = cfg_is_wg[37] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12369" *) calc_pout_53 : calc_pout_5;
  assign abuf_wr_elem_54 = cfg_is_wg[38] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12370" *) calc_pout_54 : calc_pout_6;
  assign abuf_wr_elem_55 = cfg_is_wg[39] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12371" *) calc_pout_55 : calc_pout_7;
  assign abuf_wr_elem_56 = cfg_is_wg[40] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12372" *) calc_pout_56 : calc_pout_8;
  assign abuf_wr_elem_57 = cfg_is_wg[41] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12373" *) calc_pout_57 : calc_pout_9;
  assign abuf_wr_elem_58 = cfg_is_wg[42] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12374" *) calc_pout_58 : calc_pout_10;
  assign abuf_wr_elem_59 = cfg_is_wg[43] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12375" *) calc_pout_59 : calc_pout_11;
  assign abuf_wr_elem_60 = cfg_is_wg[44] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12376" *) calc_pout_60 : calc_pout_12;
  assign abuf_wr_elem_61 = cfg_is_wg[45] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12377" *) calc_pout_61 : calc_pout_13;
  assign abuf_wr_elem_62 = cfg_is_wg[46] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12378" *) calc_pout_62 : calc_pout_14;
  assign abuf_wr_elem_63 = cfg_is_wg[47] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12379" *) calc_pout_63 : calc_pout_15;
  assign abuf_wr_elem_80 = cfg_is_wg[48] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12396" *) calc_pout_80 : calc_pout_64;
  assign abuf_wr_elem_81 = cfg_is_wg[49] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12397" *) calc_pout_81 : calc_pout_65;
  assign abuf_wr_elem_82 = cfg_is_wg[50] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12398" *) calc_pout_82 : calc_pout_66;
  assign abuf_wr_elem_83 = cfg_is_wg[51] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12399" *) calc_pout_83 : calc_pout_67;
  assign abuf_wr_elem_84 = cfg_is_wg[52] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12400" *) calc_pout_84 : calc_pout_68;
  assign abuf_wr_elem_85 = cfg_is_wg[53] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12401" *) calc_pout_85 : calc_pout_69;
  assign abuf_wr_elem_86 = cfg_is_wg[54] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12402" *) calc_pout_86 : calc_pout_70;
  assign abuf_wr_elem_87 = cfg_is_wg[55] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12403" *) calc_pout_87 : calc_pout_71;
  assign abuf_wr_elem_88 = cfg_is_wg[56] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12404" *) calc_pout_88 : calc_pout_72;
  assign abuf_wr_elem_89 = cfg_is_wg[57] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12405" *) calc_pout_89 : calc_pout_73;
  assign abuf_wr_elem_90 = cfg_is_wg[58] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12406" *) calc_pout_90 : calc_pout_74;
  assign abuf_wr_elem_91 = cfg_is_wg[59] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12407" *) calc_pout_91 : calc_pout_75;
  assign abuf_wr_elem_92 = cfg_is_wg[60] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12408" *) calc_pout_92 : calc_pout_76;
  assign abuf_wr_elem_93 = cfg_is_wg[61] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12409" *) calc_pout_93 : calc_pout_77;
  assign abuf_wr_elem_94 = cfg_is_wg[62] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12410" *) calc_pout_94 : calc_pout_78;
  assign abuf_wr_elem_95 = cfg_is_wg[63] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12411" *) calc_pout_95 : calc_pout_79;
  assign abuf_wr_elem_96 = cfg_is_wg[64] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12412" *) calc_pout_96 : calc_pout_64;
  assign abuf_wr_elem_97 = cfg_is_wg[65] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12413" *) calc_pout_97 : calc_pout_65;
  assign abuf_wr_elem_98 = cfg_is_wg[66] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12414" *) calc_pout_98 : calc_pout_66;
  assign abuf_wr_elem_99 = cfg_is_wg[67] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12415" *) calc_pout_99 : calc_pout_67;
  assign abuf_wr_elem_100 = cfg_is_wg[68] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12416" *) calc_pout_100 : calc_pout_68;
  assign abuf_wr_elem_101 = cfg_is_wg[69] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12417" *) calc_pout_101 : calc_pout_69;
  assign abuf_wr_elem_102 = cfg_is_wg[70] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12418" *) calc_pout_102 : calc_pout_70;
  assign abuf_wr_elem_103 = cfg_is_wg[71] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12419" *) calc_pout_103 : calc_pout_71;
  assign abuf_wr_elem_104 = cfg_is_wg[72] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12420" *) calc_pout_104 : calc_pout_72;
  assign abuf_wr_elem_105 = cfg_is_wg[73] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12421" *) calc_pout_105 : calc_pout_73;
  assign abuf_wr_elem_106 = cfg_is_wg[74] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12422" *) calc_pout_106 : calc_pout_74;
  assign abuf_wr_elem_107 = cfg_is_wg[75] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12423" *) calc_pout_107 : calc_pout_75;
  assign abuf_wr_elem_108 = cfg_is_wg[76] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12424" *) calc_pout_108 : calc_pout_76;
  assign abuf_wr_elem_109 = cfg_is_wg[77] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12425" *) calc_pout_109 : calc_pout_77;
  assign abuf_wr_elem_110 = cfg_is_wg[78] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12426" *) calc_pout_110 : calc_pout_78;
  assign abuf_wr_elem_111 = cfg_is_wg[79] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12427" *) calc_pout_111 : calc_pout_79;
  assign abuf_wr_elem_112 = cfg_is_wg[80] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12428" *) calc_pout_112 : calc_pout_64;
  assign abuf_wr_elem_113 = cfg_is_wg[81] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12429" *) calc_pout_113 : calc_pout_65;
  assign abuf_wr_elem_114 = cfg_is_wg[82] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12430" *) calc_pout_114 : calc_pout_66;
  assign abuf_wr_elem_115 = cfg_is_wg[83] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12431" *) calc_pout_115 : calc_pout_67;
  assign abuf_wr_elem_116 = cfg_is_wg[84] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12432" *) calc_pout_116 : calc_pout_68;
  assign abuf_wr_elem_117 = cfg_is_wg[85] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12433" *) calc_pout_117 : calc_pout_69;
  assign abuf_wr_elem_118 = cfg_is_wg[86] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12434" *) calc_pout_118 : calc_pout_70;
  assign abuf_wr_elem_119 = cfg_is_wg[87] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12435" *) calc_pout_119 : calc_pout_71;
  assign abuf_wr_elem_120 = cfg_is_wg[88] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12436" *) calc_pout_120 : calc_pout_72;
  assign abuf_wr_elem_121 = cfg_is_wg[89] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12437" *) calc_pout_121 : calc_pout_73;
  assign abuf_wr_elem_122 = cfg_is_wg[90] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12438" *) calc_pout_122 : calc_pout_74;
  assign abuf_wr_elem_123 = cfg_is_wg[91] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12439" *) calc_pout_123 : calc_pout_75;
  assign abuf_wr_elem_124 = cfg_is_wg[92] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12440" *) calc_pout_124 : calc_pout_76;
  assign abuf_wr_elem_125 = cfg_is_wg[93] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12441" *) calc_pout_125 : calc_pout_77;
  assign abuf_wr_elem_126 = cfg_is_wg[94] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12442" *) calc_pout_126 : calc_pout_78;
  assign abuf_wr_elem_127 = cfg_is_wg[95] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12443" *) calc_pout_127 : calc_pout_79;
  assign calc_dlv_elem_1 = cfg_is_int8[64] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12729" *) calc_fout_64 : calc_fout_1;
  assign calc_dlv_elem_2 = cfg_is_int8[65] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12730" *) calc_fout_1 : calc_fout_2;
  assign calc_dlv_elem_3 = cfg_is_int8[66] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12731" *) calc_fout_65 : calc_fout_3;
  assign calc_dlv_elem_4 = cfg_is_int8[67] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12732" *) calc_fout_2 : calc_fout_4;
  assign calc_dlv_elem_5 = cfg_is_int8[68] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12733" *) calc_fout_66 : calc_fout_5;
  assign calc_dlv_elem_6 = cfg_is_int8[69] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12734" *) calc_fout_3 : calc_fout_6;
  assign calc_dlv_elem_7 = cfg_is_int8[70] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12735" *) calc_fout_67 : calc_fout_7;
  assign calc_dlv_elem_8 = cfg_is_int8[71] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12736" *) calc_fout_4 : calc_fout_8;
  assign calc_dlv_elem_9 = cfg_is_int8[72] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12737" *) calc_fout_68 : calc_fout_9;
  assign calc_dlv_elem_10 = cfg_is_int8[73] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12738" *) calc_fout_5 : calc_fout_10;
  assign calc_dlv_elem_11 = cfg_is_int8[74] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12739" *) calc_fout_69 : calc_fout_11;
  assign calc_dlv_elem_12 = cfg_is_int8[75] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12740" *) calc_fout_6 : calc_fout_12;
  assign calc_dlv_elem_13 = cfg_is_int8[76] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12741" *) calc_fout_70 : calc_fout_13;
  assign calc_dlv_elem_14 = cfg_is_int8[77] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12742" *) calc_fout_7 : calc_fout_14;
  assign calc_dlv_elem_15 = cfg_is_int8[78] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12743" *) calc_fout_71 : calc_fout_15;
  assign calc_dlv_elem_16 = cfg_is_int8[79] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12744" *) calc_fout_8 : calc_fout_16;
  assign calc_dlv_elem_17 = cfg_is_int8[80] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12745" *) calc_fout_72 : calc_fout_17;
  assign calc_dlv_elem_18 = cfg_is_int8[81] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12746" *) calc_fout_9 : calc_fout_18;
  assign calc_dlv_elem_19 = cfg_is_int8[82] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12747" *) calc_fout_73 : calc_fout_19;
  assign calc_dlv_elem_20 = cfg_is_int8[83] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12748" *) calc_fout_10 : calc_fout_20;
  assign calc_dlv_elem_21 = cfg_is_int8[84] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12749" *) calc_fout_74 : calc_fout_21;
  assign calc_dlv_elem_22 = cfg_is_int8[85] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12750" *) calc_fout_11 : calc_fout_22;
  assign calc_dlv_elem_23 = cfg_is_int8[86] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12751" *) calc_fout_75 : calc_fout_23;
  assign calc_dlv_elem_24 = cfg_is_int8[87] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12752" *) calc_fout_12 : calc_fout_24;
  assign calc_dlv_elem_25 = cfg_is_int8[88] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12753" *) calc_fout_76 : calc_fout_25;
  assign calc_dlv_elem_26 = cfg_is_int8[89] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12754" *) calc_fout_13 : calc_fout_26;
  assign calc_dlv_elem_27 = cfg_is_int8[90] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12755" *) calc_fout_77 : calc_fout_27;
  assign calc_dlv_elem_28 = cfg_is_int8[91] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12756" *) calc_fout_14 : calc_fout_28;
  assign calc_dlv_elem_29 = cfg_is_int8[92] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12757" *) calc_fout_78 : calc_fout_29;
  assign calc_dlv_elem_30 = cfg_is_int8[93] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12758" *) calc_fout_15 : calc_fout_30;
  assign calc_dlv_elem_31 = cfg_is_int8[94] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12759" *) calc_fout_79 : calc_fout_31;
  assign calc_dlv_elem_32 = cfg_is_int8[95] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12760" *) calc_fout_16 : calc_fout_32;
  assign calc_dlv_elem_33 = cfg_is_int8[96] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12761" *) calc_fout_80 : calc_fout_33;
  assign calc_dlv_elem_34 = cfg_is_int8[97] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12762" *) calc_fout_17 : calc_fout_34;
  assign calc_dlv_elem_35 = cfg_is_int8[98] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12763" *) calc_fout_81 : calc_fout_35;
  assign calc_dlv_elem_36 = cfg_is_int8[99] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12764" *) calc_fout_18 : calc_fout_36;
  assign calc_dlv_elem_37 = cfg_is_int8[100] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12765" *) calc_fout_82 : calc_fout_37;
  assign calc_dlv_elem_38 = cfg_is_int8[101] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12766" *) calc_fout_19 : calc_fout_38;
  assign calc_dlv_elem_39 = cfg_is_int8[102] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12767" *) calc_fout_83 : calc_fout_39;
  assign calc_dlv_elem_40 = cfg_is_int8[103] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12768" *) calc_fout_20 : calc_fout_40;
  assign calc_dlv_elem_41 = cfg_is_int8[104] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12769" *) calc_fout_84 : calc_fout_41;
  assign calc_dlv_elem_42 = cfg_is_int8[105] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12770" *) calc_fout_21 : calc_fout_42;
  assign calc_dlv_elem_43 = cfg_is_int8[106] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12771" *) calc_fout_85 : calc_fout_43;
  assign calc_dlv_elem_44 = cfg_is_int8[107] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12772" *) calc_fout_22 : calc_fout_44;
  assign calc_dlv_elem_45 = cfg_is_int8[108] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12773" *) calc_fout_86 : calc_fout_45;
  assign calc_dlv_elem_46 = cfg_is_int8[109] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12774" *) calc_fout_23 : calc_fout_46;
  assign calc_dlv_elem_47 = cfg_is_int8[110] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12775" *) calc_fout_87 : calc_fout_47;
  assign calc_dlv_elem_48 = cfg_is_int8[111] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12776" *) calc_fout_24 : calc_fout_48;
  assign calc_dlv_elem_49 = cfg_is_int8[112] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12777" *) calc_fout_88 : calc_fout_49;
  assign calc_dlv_elem_50 = cfg_is_int8[113] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12778" *) calc_fout_25 : calc_fout_50;
  assign calc_dlv_elem_51 = cfg_is_int8[114] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12779" *) calc_fout_89 : calc_fout_51;
  assign calc_dlv_elem_52 = cfg_is_int8[115] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12780" *) calc_fout_26 : calc_fout_52;
  assign calc_dlv_elem_53 = cfg_is_int8[116] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12781" *) calc_fout_90 : calc_fout_53;
  assign calc_dlv_elem_54 = cfg_is_int8[117] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12782" *) calc_fout_27 : calc_fout_54;
  assign calc_dlv_elem_55 = cfg_is_int8[118] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12783" *) calc_fout_91 : calc_fout_55;
  assign calc_dlv_elem_56 = cfg_is_int8[119] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12784" *) calc_fout_28 : calc_fout_56;
  assign calc_dlv_elem_57 = cfg_is_int8[120] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12785" *) calc_fout_92 : calc_fout_57;
  assign calc_dlv_elem_58 = cfg_is_int8[121] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12786" *) calc_fout_29 : calc_fout_58;
  assign calc_dlv_elem_59 = cfg_is_int8[122] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12787" *) calc_fout_93 : calc_fout_59;
  assign calc_dlv_elem_60 = cfg_is_int8[123] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12788" *) calc_fout_30 : calc_fout_60;
  assign calc_dlv_elem_61 = cfg_is_int8[124] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12789" *) calc_fout_94 : calc_fout_61;
  assign calc_dlv_elem_62 = cfg_is_int8[125] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12790" *) calc_fout_31 : calc_fout_62;
  assign calc_dlv_elem_63 = cfg_is_int8[126] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:12791" *) calc_fout_95 : calc_fout_63;
  assign _0910_ = sat_carry ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13419" *) 32'd4294967295 : sat_count_inc;
  assign sat_count_w = dlv_sat_clr_d1 ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:13419" *) { 24'b000000000000000000000000, sat_sum } : _0910_;
  assign calc_elem_0_w = cfg_is_int8[0] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2989" *) { calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21:0] } : calc_data_0[43:0];
  assign calc_elem_1_w = cfg_is_int8[1] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2990" *) { calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21:0] } : calc_data_1[43:0];
  assign calc_elem_2_w = cfg_is_int8[2] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2991" *) { calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21:0] } : calc_data_2[43:0];
  assign calc_elem_3_w = cfg_is_int8[3] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2992" *) { calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21:0] } : calc_data_3[43:0];
  assign calc_elem_4_w = cfg_is_int8[4] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2993" *) { calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21:0] } : calc_data_4[43:0];
  assign calc_elem_5_w = cfg_is_int8[5] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2994" *) { calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21:0] } : calc_data_5[43:0];
  assign calc_elem_6_w = cfg_is_int8[6] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2995" *) { calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21:0] } : calc_data_6[43:0];
  assign calc_elem_7_w = cfg_is_int8[7] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2996" *) { calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21:0] } : calc_data_7[43:0];
  assign calc_elem_8_w = cfg_is_int8[8] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2997" *) { calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21:0] } : calc_data_8[43:0];
  assign calc_elem_9_w = cfg_is_int8[9] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2998" *) { calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21:0] } : calc_data_9[43:0];
  assign calc_elem_10_w = cfg_is_int8[10] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:2999" *) { calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21:0] } : calc_data_10[43:0];
  assign calc_elem_11_w = cfg_is_int8[11] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3000" *) { calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21:0] } : calc_data_11[43:0];
  assign calc_elem_12_w = cfg_is_int8[12] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3001" *) { calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21:0] } : calc_data_12[43:0];
  assign calc_elem_13_w = cfg_is_int8[13] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3002" *) { calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21:0] } : calc_data_13[43:0];
  assign calc_elem_14_w = cfg_is_int8[14] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3003" *) { calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21:0] } : calc_data_14[43:0];
  assign calc_elem_15_w = cfg_is_int8[15] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3004" *) { calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21:0] } : calc_data_15[43:0];
  assign calc_elem_16_w = cfg_is_int8[16] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3005" *) { calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65:44] } : calc_data_0[87:44];
  assign calc_elem_17_w = cfg_is_int8[17] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3006" *) { calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65:44] } : calc_data_1[87:44];
  assign calc_elem_18_w = cfg_is_int8[18] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3007" *) { calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65:44] } : calc_data_2[87:44];
  assign calc_elem_19_w = cfg_is_int8[19] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3008" *) { calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65:44] } : calc_data_3[87:44];
  assign calc_elem_20_w = cfg_is_int8[20] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3009" *) { calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65:44] } : calc_data_4[87:44];
  assign calc_elem_21_w = cfg_is_int8[21] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3010" *) { calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65:44] } : calc_data_5[87:44];
  assign calc_elem_22_w = cfg_is_int8[22] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3011" *) { calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65:44] } : calc_data_6[87:44];
  assign calc_elem_23_w = cfg_is_int8[23] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3012" *) { calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65:44] } : calc_data_7[87:44];
  assign calc_elem_24_w = cfg_is_int8[24] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3013" *) { calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65:44] } : calc_data_8[87:44];
  assign calc_elem_25_w = cfg_is_int8[25] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3014" *) { calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65:44] } : calc_data_9[87:44];
  assign calc_elem_26_w = cfg_is_int8[26] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3015" *) { calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65:44] } : calc_data_10[87:44];
  assign calc_elem_27_w = cfg_is_int8[27] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3016" *) { calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65:44] } : calc_data_11[87:44];
  assign calc_elem_28_w = cfg_is_int8[28] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3017" *) { calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65:44] } : calc_data_12[87:44];
  assign calc_elem_29_w = cfg_is_int8[29] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3018" *) { calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65:44] } : calc_data_13[87:44];
  assign calc_elem_30_w = cfg_is_int8[30] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3019" *) { calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65:44] } : calc_data_14[87:44];
  assign calc_elem_31_w = cfg_is_int8[31] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3020" *) { calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65:44] } : calc_data_15[87:44];
  assign calc_elem_32_w = cfg_is_int8[32] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3021" *) { calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109:88] } : calc_data_0[131:88];
  assign calc_elem_33_w = cfg_is_int8[33] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3022" *) { calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109:88] } : calc_data_1[131:88];
  assign calc_elem_34_w = cfg_is_int8[34] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3023" *) { calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109:88] } : calc_data_2[131:88];
  assign calc_elem_35_w = cfg_is_int8[35] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3024" *) { calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109:88] } : calc_data_3[131:88];
  assign calc_elem_36_w = cfg_is_int8[36] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3025" *) { calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109:88] } : calc_data_4[131:88];
  assign calc_elem_37_w = cfg_is_int8[37] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3026" *) { calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109:88] } : calc_data_5[131:88];
  assign calc_elem_38_w = cfg_is_int8[38] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3027" *) { calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109:88] } : calc_data_6[131:88];
  assign calc_elem_39_w = cfg_is_int8[39] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3028" *) { calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109:88] } : calc_data_7[131:88];
  assign calc_elem_40_w = cfg_is_int8[40] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3029" *) { calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109:88] } : calc_data_8[131:88];
  assign calc_elem_41_w = cfg_is_int8[41] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3030" *) { calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109:88] } : calc_data_9[131:88];
  assign calc_elem_42_w = cfg_is_int8[42] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3031" *) { calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109:88] } : calc_data_10[131:88];
  assign calc_elem_43_w = cfg_is_int8[43] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3032" *) { calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109:88] } : calc_data_11[131:88];
  assign calc_elem_44_w = cfg_is_int8[44] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3033" *) { calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109:88] } : calc_data_12[131:88];
  assign calc_elem_45_w = cfg_is_int8[45] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3034" *) { calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109:88] } : calc_data_13[131:88];
  assign calc_elem_46_w = cfg_is_int8[46] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3035" *) { calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109:88] } : calc_data_14[131:88];
  assign calc_elem_47_w = cfg_is_int8[47] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3036" *) { calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109:88] } : calc_data_15[131:88];
  assign calc_elem_48_w = cfg_is_int8[48] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3037" *) { calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153:132] } : calc_data_0[175:132];
  assign calc_elem_49_w = cfg_is_int8[49] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3038" *) { calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153:132] } : calc_data_1[175:132];
  assign calc_elem_50_w = cfg_is_int8[50] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3039" *) { calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153:132] } : calc_data_2[175:132];
  assign calc_elem_51_w = cfg_is_int8[51] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3040" *) { calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153:132] } : calc_data_3[175:132];
  assign calc_elem_52_w = cfg_is_int8[52] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3041" *) { calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153:132] } : calc_data_4[175:132];
  assign calc_elem_53_w = cfg_is_int8[53] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3042" *) { calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153:132] } : calc_data_5[175:132];
  assign calc_elem_54_w = cfg_is_int8[54] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3043" *) { calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153:132] } : calc_data_6[175:132];
  assign calc_elem_55_w = cfg_is_int8[55] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3044" *) { calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153:132] } : calc_data_7[175:132];
  assign calc_elem_56_w = cfg_is_int8[56] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3045" *) { calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153:132] } : calc_data_8[175:132];
  assign calc_elem_57_w = cfg_is_int8[57] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3046" *) { calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153:132] } : calc_data_9[175:132];
  assign calc_elem_58_w = cfg_is_int8[58] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3047" *) { calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153:132] } : calc_data_10[175:132];
  assign calc_elem_59_w = cfg_is_int8[59] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3048" *) { calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153:132] } : calc_data_11[175:132];
  assign calc_elem_60_w = cfg_is_int8[60] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3049" *) { calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153:132] } : calc_data_12[175:132];
  assign calc_elem_61_w = cfg_is_int8[61] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3050" *) { calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153:132] } : calc_data_13[175:132];
  assign calc_elem_62_w = cfg_is_int8[62] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3051" *) { calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153:132] } : calc_data_14[175:132];
  assign calc_elem_63_w = cfg_is_int8[63] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3052" *) { calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153:132] } : calc_data_15[175:132];
  assign _0911_ = accu_ctrl_pd[7] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *) 8'b00001111 : 8'b11111111;
  assign _0912_ = accu_ctrl_pd[6] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *) 8'b00000011 : _0911_;
  assign _0913_ = accu_ctrl_pd[5] ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *) 8'b00000001 : _0912_;
  assign calc_dlv_en = _0907_ ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3209" *) 8'b00000000 : _0913_;
  assign calc_wr_en = _0908_ ? (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:3217" *) 8'b00000000 : accu_ctrl_pd[16:9];
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9678" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_0 (
    .in_data(calc_op0_fp_0_d1),
    .in_op(calc_op1_fp_0_d1),
    .in_op_valid(calc_op1_vld_fp_d1[0]),
    .in_sel(calc_dlv_en_fp_d1[0]),
    .in_valid(calc_op_en_fp_d1[0]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_0_sum),
    .out_final_valid(calc_fout_fp_vld[0]),
    .out_partial_data(calc_pout_fp_0_sum),
    .out_partial_valid(calc_pout_fp_vld[0])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9691" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_1 (
    .in_data(calc_op0_fp_1_d1),
    .in_op(calc_op1_fp_1_d1),
    .in_op_valid(calc_op1_vld_fp_d1[1]),
    .in_sel(calc_dlv_en_fp_d1[1]),
    .in_valid(calc_op_en_fp_d1[1]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_1_sum),
    .out_final_valid(calc_fout_fp_vld[1]),
    .out_partial_data(calc_pout_fp_1_sum),
    .out_partial_valid(calc_pout_fp_vld[1])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9808" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_10 (
    .in_data(calc_op0_fp_10_d1),
    .in_op(calc_op1_fp_10_d1),
    .in_op_valid(calc_op1_vld_fp_d1[10]),
    .in_sel(calc_dlv_en_fp_d1[10]),
    .in_valid(calc_op_en_fp_d1[10]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_10_sum),
    .out_final_valid(calc_fout_fp_vld[10]),
    .out_partial_data(calc_pout_fp_10_sum),
    .out_partial_valid(calc_pout_fp_vld[10])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9821" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_11 (
    .in_data(calc_op0_fp_11_d1),
    .in_op(calc_op1_fp_11_d1),
    .in_op_valid(calc_op1_vld_fp_d1[11]),
    .in_sel(calc_dlv_en_fp_d1[11]),
    .in_valid(calc_op_en_fp_d1[11]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_11_sum),
    .out_final_valid(calc_fout_fp_vld[11]),
    .out_partial_data(calc_pout_fp_11_sum),
    .out_partial_valid(calc_pout_fp_vld[11])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9834" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_12 (
    .in_data(calc_op0_fp_12_d1),
    .in_op(calc_op1_fp_12_d1),
    .in_op_valid(calc_op1_vld_fp_d1[12]),
    .in_sel(calc_dlv_en_fp_d1[12]),
    .in_valid(calc_op_en_fp_d1[12]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_12_sum),
    .out_final_valid(calc_fout_fp_vld[12]),
    .out_partial_data(calc_pout_fp_12_sum),
    .out_partial_valid(calc_pout_fp_vld[12])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9847" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_13 (
    .in_data(calc_op0_fp_13_d1),
    .in_op(calc_op1_fp_13_d1),
    .in_op_valid(calc_op1_vld_fp_d1[13]),
    .in_sel(calc_dlv_en_fp_d1[13]),
    .in_valid(calc_op_en_fp_d1[13]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_13_sum),
    .out_final_valid(calc_fout_fp_vld[13]),
    .out_partial_data(calc_pout_fp_13_sum),
    .out_partial_valid(calc_pout_fp_vld[13])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9860" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_14 (
    .in_data(calc_op0_fp_14_d1),
    .in_op(calc_op1_fp_14_d1),
    .in_op_valid(calc_op1_vld_fp_d1[14]),
    .in_sel(calc_dlv_en_fp_d1[14]),
    .in_valid(calc_op_en_fp_d1[14]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_14_sum),
    .out_final_valid(calc_fout_fp_vld[14]),
    .out_partial_data(calc_pout_fp_14_sum),
    .out_partial_valid(calc_pout_fp_vld[14])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9873" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_15 (
    .in_data(calc_op0_fp_15_d1),
    .in_op(calc_op1_fp_15_d1),
    .in_op_valid(calc_op1_vld_fp_d1[15]),
    .in_sel(calc_dlv_en_fp_d1[15]),
    .in_valid(calc_op_en_fp_d1[15]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_15_sum),
    .out_final_valid(calc_fout_fp_vld[15]),
    .out_partial_data(calc_pout_fp_15_sum),
    .out_partial_valid(calc_pout_fp_vld[15])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9886" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_16 (
    .in_data(calc_op0_fp_16_d1),
    .in_op(calc_op1_fp_16_d1),
    .in_op_valid(calc_op1_vld_fp_d1[16]),
    .in_sel(calc_dlv_en_fp_d1[16]),
    .in_valid(calc_op_en_fp_d1[16]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_16_sum),
    .out_final_valid(calc_fout_fp_vld[16]),
    .out_partial_data(calc_pout_fp_16_sum),
    .out_partial_valid(calc_pout_fp_vld[16])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9899" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_17 (
    .in_data(calc_op0_fp_17_d1),
    .in_op(calc_op1_fp_17_d1),
    .in_op_valid(calc_op1_vld_fp_d1[17]),
    .in_sel(calc_dlv_en_fp_d1[17]),
    .in_valid(calc_op_en_fp_d1[17]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_17_sum),
    .out_final_valid(calc_fout_fp_vld[17]),
    .out_partial_data(calc_pout_fp_17_sum),
    .out_partial_valid(calc_pout_fp_vld[17])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9912" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_18 (
    .in_data(calc_op0_fp_18_d1),
    .in_op(calc_op1_fp_18_d1),
    .in_op_valid(calc_op1_vld_fp_d1[18]),
    .in_sel(calc_dlv_en_fp_d1[18]),
    .in_valid(calc_op_en_fp_d1[18]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_18_sum),
    .out_final_valid(calc_fout_fp_vld[18]),
    .out_partial_data(calc_pout_fp_18_sum),
    .out_partial_valid(calc_pout_fp_vld[18])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9925" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_19 (
    .in_data(calc_op0_fp_19_d1),
    .in_op(calc_op1_fp_19_d1),
    .in_op_valid(calc_op1_vld_fp_d1[19]),
    .in_sel(calc_dlv_en_fp_d1[19]),
    .in_valid(calc_op_en_fp_d1[19]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_19_sum),
    .out_final_valid(calc_fout_fp_vld[19]),
    .out_partial_data(calc_pout_fp_19_sum),
    .out_partial_valid(calc_pout_fp_vld[19])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9704" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_2 (
    .in_data(calc_op0_fp_2_d1),
    .in_op(calc_op1_fp_2_d1),
    .in_op_valid(calc_op1_vld_fp_d1[2]),
    .in_sel(calc_dlv_en_fp_d1[2]),
    .in_valid(calc_op_en_fp_d1[2]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_2_sum),
    .out_final_valid(calc_fout_fp_vld[2]),
    .out_partial_data(calc_pout_fp_2_sum),
    .out_partial_valid(calc_pout_fp_vld[2])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9938" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_20 (
    .in_data(calc_op0_fp_20_d1),
    .in_op(calc_op1_fp_20_d1),
    .in_op_valid(calc_op1_vld_fp_d1[20]),
    .in_sel(calc_dlv_en_fp_d1[20]),
    .in_valid(calc_op_en_fp_d1[20]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_20_sum),
    .out_final_valid(calc_fout_fp_vld[20]),
    .out_partial_data(calc_pout_fp_20_sum),
    .out_partial_valid(calc_pout_fp_vld[20])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9951" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_21 (
    .in_data(calc_op0_fp_21_d1),
    .in_op(calc_op1_fp_21_d1),
    .in_op_valid(calc_op1_vld_fp_d1[21]),
    .in_sel(calc_dlv_en_fp_d1[21]),
    .in_valid(calc_op_en_fp_d1[21]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_21_sum),
    .out_final_valid(calc_fout_fp_vld[21]),
    .out_partial_data(calc_pout_fp_21_sum),
    .out_partial_valid(calc_pout_fp_vld[21])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9964" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_22 (
    .in_data(calc_op0_fp_22_d1),
    .in_op(calc_op1_fp_22_d1),
    .in_op_valid(calc_op1_vld_fp_d1[22]),
    .in_sel(calc_dlv_en_fp_d1[22]),
    .in_valid(calc_op_en_fp_d1[22]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_22_sum),
    .out_final_valid(calc_fout_fp_vld[22]),
    .out_partial_data(calc_pout_fp_22_sum),
    .out_partial_valid(calc_pout_fp_vld[22])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9977" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_23 (
    .in_data(calc_op0_fp_23_d1),
    .in_op(calc_op1_fp_23_d1),
    .in_op_valid(calc_op1_vld_fp_d1[23]),
    .in_sel(calc_dlv_en_fp_d1[23]),
    .in_valid(calc_op_en_fp_d1[23]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_23_sum),
    .out_final_valid(calc_fout_fp_vld[23]),
    .out_partial_data(calc_pout_fp_23_sum),
    .out_partial_valid(calc_pout_fp_vld[23])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9990" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_24 (
    .in_data(calc_op0_fp_24_d1),
    .in_op(calc_op1_fp_24_d1),
    .in_op_valid(calc_op1_vld_fp_d1[24]),
    .in_sel(calc_dlv_en_fp_d1[24]),
    .in_valid(calc_op_en_fp_d1[24]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_24_sum),
    .out_final_valid(calc_fout_fp_vld[24]),
    .out_partial_data(calc_pout_fp_24_sum),
    .out_partial_valid(calc_pout_fp_vld[24])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10003" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_25 (
    .in_data(calc_op0_fp_25_d1),
    .in_op(calc_op1_fp_25_d1),
    .in_op_valid(calc_op1_vld_fp_d1[25]),
    .in_sel(calc_dlv_en_fp_d1[25]),
    .in_valid(calc_op_en_fp_d1[25]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_25_sum),
    .out_final_valid(calc_fout_fp_vld[25]),
    .out_partial_data(calc_pout_fp_25_sum),
    .out_partial_valid(calc_pout_fp_vld[25])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10016" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_26 (
    .in_data(calc_op0_fp_26_d1),
    .in_op(calc_op1_fp_26_d1),
    .in_op_valid(calc_op1_vld_fp_d1[26]),
    .in_sel(calc_dlv_en_fp_d1[26]),
    .in_valid(calc_op_en_fp_d1[26]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_26_sum),
    .out_final_valid(calc_fout_fp_vld[26]),
    .out_partial_data(calc_pout_fp_26_sum),
    .out_partial_valid(calc_pout_fp_vld[26])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10029" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_27 (
    .in_data(calc_op0_fp_27_d1),
    .in_op(calc_op1_fp_27_d1),
    .in_op_valid(calc_op1_vld_fp_d1[27]),
    .in_sel(calc_dlv_en_fp_d1[27]),
    .in_valid(calc_op_en_fp_d1[27]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_27_sum),
    .out_final_valid(calc_fout_fp_vld[27]),
    .out_partial_data(calc_pout_fp_27_sum),
    .out_partial_valid(calc_pout_fp_vld[27])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10042" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_28 (
    .in_data(calc_op0_fp_28_d1),
    .in_op(calc_op1_fp_28_d1),
    .in_op_valid(calc_op1_vld_fp_d1[28]),
    .in_sel(calc_dlv_en_fp_d1[28]),
    .in_valid(calc_op_en_fp_d1[28]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_28_sum),
    .out_final_valid(calc_fout_fp_vld[28]),
    .out_partial_data(calc_pout_fp_28_sum),
    .out_partial_valid(calc_pout_fp_vld[28])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10055" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_29 (
    .in_data(calc_op0_fp_29_d1),
    .in_op(calc_op1_fp_29_d1),
    .in_op_valid(calc_op1_vld_fp_d1[29]),
    .in_sel(calc_dlv_en_fp_d1[29]),
    .in_valid(calc_op_en_fp_d1[29]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_29_sum),
    .out_final_valid(calc_fout_fp_vld[29]),
    .out_partial_data(calc_pout_fp_29_sum),
    .out_partial_valid(calc_pout_fp_vld[29])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9717" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_3 (
    .in_data(calc_op0_fp_3_d1),
    .in_op(calc_op1_fp_3_d1),
    .in_op_valid(calc_op1_vld_fp_d1[3]),
    .in_sel(calc_dlv_en_fp_d1[3]),
    .in_valid(calc_op_en_fp_d1[3]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_3_sum),
    .out_final_valid(calc_fout_fp_vld[3]),
    .out_partial_data(calc_pout_fp_3_sum),
    .out_partial_valid(calc_pout_fp_vld[3])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10068" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_30 (
    .in_data(calc_op0_fp_30_d1),
    .in_op(calc_op1_fp_30_d1),
    .in_op_valid(calc_op1_vld_fp_d1[30]),
    .in_sel(calc_dlv_en_fp_d1[30]),
    .in_valid(calc_op_en_fp_d1[30]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_30_sum),
    .out_final_valid(calc_fout_fp_vld[30]),
    .out_partial_data(calc_pout_fp_30_sum),
    .out_partial_valid(calc_pout_fp_vld[30])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10081" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_31 (
    .in_data(calc_op0_fp_31_d1),
    .in_op(calc_op1_fp_31_d1),
    .in_op_valid(calc_op1_vld_fp_d1[31]),
    .in_sel(calc_dlv_en_fp_d1[31]),
    .in_valid(calc_op_en_fp_d1[31]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_31_sum),
    .out_final_valid(calc_fout_fp_vld[31]),
    .out_partial_data(calc_pout_fp_31_sum),
    .out_partial_valid(calc_pout_fp_vld[31])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10094" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_32 (
    .in_data(calc_op0_fp_32_d1),
    .in_op(calc_op1_fp_32_d1),
    .in_op_valid(calc_op1_vld_fp_d1[32]),
    .in_sel(calc_dlv_en_fp_d1[32]),
    .in_valid(calc_op_en_fp_d1[32]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_32_sum),
    .out_final_valid(calc_fout_fp_vld[32]),
    .out_partial_data(calc_pout_fp_32_sum),
    .out_partial_valid(calc_pout_fp_vld[32])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10107" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_33 (
    .in_data(calc_op0_fp_33_d1),
    .in_op(calc_op1_fp_33_d1),
    .in_op_valid(calc_op1_vld_fp_d1[33]),
    .in_sel(calc_dlv_en_fp_d1[33]),
    .in_valid(calc_op_en_fp_d1[33]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_33_sum),
    .out_final_valid(calc_fout_fp_vld[33]),
    .out_partial_data(calc_pout_fp_33_sum),
    .out_partial_valid(calc_pout_fp_vld[33])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10120" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_34 (
    .in_data(calc_op0_fp_34_d1),
    .in_op(calc_op1_fp_34_d1),
    .in_op_valid(calc_op1_vld_fp_d1[34]),
    .in_sel(calc_dlv_en_fp_d1[34]),
    .in_valid(calc_op_en_fp_d1[34]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_34_sum),
    .out_final_valid(calc_fout_fp_vld[34]),
    .out_partial_data(calc_pout_fp_34_sum),
    .out_partial_valid(calc_pout_fp_vld[34])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10133" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_35 (
    .in_data(calc_op0_fp_35_d1),
    .in_op(calc_op1_fp_35_d1),
    .in_op_valid(calc_op1_vld_fp_d1[35]),
    .in_sel(calc_dlv_en_fp_d1[35]),
    .in_valid(calc_op_en_fp_d1[35]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_35_sum),
    .out_final_valid(calc_fout_fp_vld[35]),
    .out_partial_data(calc_pout_fp_35_sum),
    .out_partial_valid(calc_pout_fp_vld[35])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10146" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_36 (
    .in_data(calc_op0_fp_36_d1),
    .in_op(calc_op1_fp_36_d1),
    .in_op_valid(calc_op1_vld_fp_d1[36]),
    .in_sel(calc_dlv_en_fp_d1[36]),
    .in_valid(calc_op_en_fp_d1[36]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_36_sum),
    .out_final_valid(calc_fout_fp_vld[36]),
    .out_partial_data(calc_pout_fp_36_sum),
    .out_partial_valid(calc_pout_fp_vld[36])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10159" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_37 (
    .in_data(calc_op0_fp_37_d1),
    .in_op(calc_op1_fp_37_d1),
    .in_op_valid(calc_op1_vld_fp_d1[37]),
    .in_sel(calc_dlv_en_fp_d1[37]),
    .in_valid(calc_op_en_fp_d1[37]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_37_sum),
    .out_final_valid(calc_fout_fp_vld[37]),
    .out_partial_data(calc_pout_fp_37_sum),
    .out_partial_valid(calc_pout_fp_vld[37])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10172" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_38 (
    .in_data(calc_op0_fp_38_d1),
    .in_op(calc_op1_fp_38_d1),
    .in_op_valid(calc_op1_vld_fp_d1[38]),
    .in_sel(calc_dlv_en_fp_d1[38]),
    .in_valid(calc_op_en_fp_d1[38]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_38_sum),
    .out_final_valid(calc_fout_fp_vld[38]),
    .out_partial_data(calc_pout_fp_38_sum),
    .out_partial_valid(calc_pout_fp_vld[38])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10185" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_39 (
    .in_data(calc_op0_fp_39_d1),
    .in_op(calc_op1_fp_39_d1),
    .in_op_valid(calc_op1_vld_fp_d1[39]),
    .in_sel(calc_dlv_en_fp_d1[39]),
    .in_valid(calc_op_en_fp_d1[39]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_39_sum),
    .out_final_valid(calc_fout_fp_vld[39]),
    .out_partial_data(calc_pout_fp_39_sum),
    .out_partial_valid(calc_pout_fp_vld[39])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9730" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_4 (
    .in_data(calc_op0_fp_4_d1),
    .in_op(calc_op1_fp_4_d1),
    .in_op_valid(calc_op1_vld_fp_d1[4]),
    .in_sel(calc_dlv_en_fp_d1[4]),
    .in_valid(calc_op_en_fp_d1[4]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_4_sum),
    .out_final_valid(calc_fout_fp_vld[4]),
    .out_partial_data(calc_pout_fp_4_sum),
    .out_partial_valid(calc_pout_fp_vld[4])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10198" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_40 (
    .in_data(calc_op0_fp_40_d1),
    .in_op(calc_op1_fp_40_d1),
    .in_op_valid(calc_op1_vld_fp_d1[40]),
    .in_sel(calc_dlv_en_fp_d1[40]),
    .in_valid(calc_op_en_fp_d1[40]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_40_sum),
    .out_final_valid(calc_fout_fp_vld[40]),
    .out_partial_data(calc_pout_fp_40_sum),
    .out_partial_valid(calc_pout_fp_vld[40])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10211" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_41 (
    .in_data(calc_op0_fp_41_d1),
    .in_op(calc_op1_fp_41_d1),
    .in_op_valid(calc_op1_vld_fp_d1[41]),
    .in_sel(calc_dlv_en_fp_d1[41]),
    .in_valid(calc_op_en_fp_d1[41]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_41_sum),
    .out_final_valid(calc_fout_fp_vld[41]),
    .out_partial_data(calc_pout_fp_41_sum),
    .out_partial_valid(calc_pout_fp_vld[41])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10224" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_42 (
    .in_data(calc_op0_fp_42_d1),
    .in_op(calc_op1_fp_42_d1),
    .in_op_valid(calc_op1_vld_fp_d1[42]),
    .in_sel(calc_dlv_en_fp_d1[42]),
    .in_valid(calc_op_en_fp_d1[42]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_42_sum),
    .out_final_valid(calc_fout_fp_vld[42]),
    .out_partial_data(calc_pout_fp_42_sum),
    .out_partial_valid(calc_pout_fp_vld[42])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10237" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_43 (
    .in_data(calc_op0_fp_43_d1),
    .in_op(calc_op1_fp_43_d1),
    .in_op_valid(calc_op1_vld_fp_d1[43]),
    .in_sel(calc_dlv_en_fp_d1[43]),
    .in_valid(calc_op_en_fp_d1[43]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_43_sum),
    .out_final_valid(calc_fout_fp_vld[43]),
    .out_partial_data(calc_pout_fp_43_sum),
    .out_partial_valid(calc_pout_fp_vld[43])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10250" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_44 (
    .in_data(calc_op0_fp_44_d1),
    .in_op(calc_op1_fp_44_d1),
    .in_op_valid(calc_op1_vld_fp_d1[44]),
    .in_sel(calc_dlv_en_fp_d1[44]),
    .in_valid(calc_op_en_fp_d1[44]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_44_sum),
    .out_final_valid(calc_fout_fp_vld[44]),
    .out_partial_data(calc_pout_fp_44_sum),
    .out_partial_valid(calc_pout_fp_vld[44])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10263" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_45 (
    .in_data(calc_op0_fp_45_d1),
    .in_op(calc_op1_fp_45_d1),
    .in_op_valid(calc_op1_vld_fp_d1[45]),
    .in_sel(calc_dlv_en_fp_d1[45]),
    .in_valid(calc_op_en_fp_d1[45]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_45_sum),
    .out_final_valid(calc_fout_fp_vld[45]),
    .out_partial_data(calc_pout_fp_45_sum),
    .out_partial_valid(calc_pout_fp_vld[45])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10276" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_46 (
    .in_data(calc_op0_fp_46_d1),
    .in_op(calc_op1_fp_46_d1),
    .in_op_valid(calc_op1_vld_fp_d1[46]),
    .in_sel(calc_dlv_en_fp_d1[46]),
    .in_valid(calc_op_en_fp_d1[46]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_46_sum),
    .out_final_valid(calc_fout_fp_vld[46]),
    .out_partial_data(calc_pout_fp_46_sum),
    .out_partial_valid(calc_pout_fp_vld[46])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10289" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_47 (
    .in_data(calc_op0_fp_47_d1),
    .in_op(calc_op1_fp_47_d1),
    .in_op_valid(calc_op1_vld_fp_d1[47]),
    .in_sel(calc_dlv_en_fp_d1[47]),
    .in_valid(calc_op_en_fp_d1[47]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_47_sum),
    .out_final_valid(calc_fout_fp_vld[47]),
    .out_partial_data(calc_pout_fp_47_sum),
    .out_partial_valid(calc_pout_fp_vld[47])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10302" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_48 (
    .in_data(calc_op0_fp_48_d1),
    .in_op(calc_op1_fp_48_d1),
    .in_op_valid(calc_op1_vld_fp_d1[48]),
    .in_sel(calc_dlv_en_fp_d1[48]),
    .in_valid(calc_op_en_fp_d1[48]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_48_sum),
    .out_final_valid(calc_fout_fp_vld[48]),
    .out_partial_data(calc_pout_fp_48_sum),
    .out_partial_valid(calc_pout_fp_vld[48])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10315" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_49 (
    .in_data(calc_op0_fp_49_d1),
    .in_op(calc_op1_fp_49_d1),
    .in_op_valid(calc_op1_vld_fp_d1[49]),
    .in_sel(calc_dlv_en_fp_d1[49]),
    .in_valid(calc_op_en_fp_d1[49]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_49_sum),
    .out_final_valid(calc_fout_fp_vld[49]),
    .out_partial_data(calc_pout_fp_49_sum),
    .out_partial_valid(calc_pout_fp_vld[49])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9743" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_5 (
    .in_data(calc_op0_fp_5_d1),
    .in_op(calc_op1_fp_5_d1),
    .in_op_valid(calc_op1_vld_fp_d1[5]),
    .in_sel(calc_dlv_en_fp_d1[5]),
    .in_valid(calc_op_en_fp_d1[5]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_5_sum),
    .out_final_valid(calc_fout_fp_vld[5]),
    .out_partial_data(calc_pout_fp_5_sum),
    .out_partial_valid(calc_pout_fp_vld[5])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10328" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_50 (
    .in_data(calc_op0_fp_50_d1),
    .in_op(calc_op1_fp_50_d1),
    .in_op_valid(calc_op1_vld_fp_d1[50]),
    .in_sel(calc_dlv_en_fp_d1[50]),
    .in_valid(calc_op_en_fp_d1[50]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_50_sum),
    .out_final_valid(calc_fout_fp_vld[50]),
    .out_partial_data(calc_pout_fp_50_sum),
    .out_partial_valid(calc_pout_fp_vld[50])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10341" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_51 (
    .in_data(calc_op0_fp_51_d1),
    .in_op(calc_op1_fp_51_d1),
    .in_op_valid(calc_op1_vld_fp_d1[51]),
    .in_sel(calc_dlv_en_fp_d1[51]),
    .in_valid(calc_op_en_fp_d1[51]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_51_sum),
    .out_final_valid(calc_fout_fp_vld[51]),
    .out_partial_data(calc_pout_fp_51_sum),
    .out_partial_valid(calc_pout_fp_vld[51])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10354" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_52 (
    .in_data(calc_op0_fp_52_d1),
    .in_op(calc_op1_fp_52_d1),
    .in_op_valid(calc_op1_vld_fp_d1[52]),
    .in_sel(calc_dlv_en_fp_d1[52]),
    .in_valid(calc_op_en_fp_d1[52]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_52_sum),
    .out_final_valid(calc_fout_fp_vld[52]),
    .out_partial_data(calc_pout_fp_52_sum),
    .out_partial_valid(calc_pout_fp_vld[52])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10367" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_53 (
    .in_data(calc_op0_fp_53_d1),
    .in_op(calc_op1_fp_53_d1),
    .in_op_valid(calc_op1_vld_fp_d1[53]),
    .in_sel(calc_dlv_en_fp_d1[53]),
    .in_valid(calc_op_en_fp_d1[53]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_53_sum),
    .out_final_valid(calc_fout_fp_vld[53]),
    .out_partial_data(calc_pout_fp_53_sum),
    .out_partial_valid(calc_pout_fp_vld[53])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10380" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_54 (
    .in_data(calc_op0_fp_54_d1),
    .in_op(calc_op1_fp_54_d1),
    .in_op_valid(calc_op1_vld_fp_d1[54]),
    .in_sel(calc_dlv_en_fp_d1[54]),
    .in_valid(calc_op_en_fp_d1[54]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_54_sum),
    .out_final_valid(calc_fout_fp_vld[54]),
    .out_partial_data(calc_pout_fp_54_sum),
    .out_partial_valid(calc_pout_fp_vld[54])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10393" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_55 (
    .in_data(calc_op0_fp_55_d1),
    .in_op(calc_op1_fp_55_d1),
    .in_op_valid(calc_op1_vld_fp_d1[55]),
    .in_sel(calc_dlv_en_fp_d1[55]),
    .in_valid(calc_op_en_fp_d1[55]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_55_sum),
    .out_final_valid(calc_fout_fp_vld[55]),
    .out_partial_data(calc_pout_fp_55_sum),
    .out_partial_valid(calc_pout_fp_vld[55])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10406" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_56 (
    .in_data(calc_op0_fp_56_d1),
    .in_op(calc_op1_fp_56_d1),
    .in_op_valid(calc_op1_vld_fp_d1[56]),
    .in_sel(calc_dlv_en_fp_d1[56]),
    .in_valid(calc_op_en_fp_d1[56]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_56_sum),
    .out_final_valid(calc_fout_fp_vld[56]),
    .out_partial_data(calc_pout_fp_56_sum),
    .out_partial_valid(calc_pout_fp_vld[56])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10419" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_57 (
    .in_data(calc_op0_fp_57_d1),
    .in_op(calc_op1_fp_57_d1),
    .in_op_valid(calc_op1_vld_fp_d1[57]),
    .in_sel(calc_dlv_en_fp_d1[57]),
    .in_valid(calc_op_en_fp_d1[57]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_57_sum),
    .out_final_valid(calc_fout_fp_vld[57]),
    .out_partial_data(calc_pout_fp_57_sum),
    .out_partial_valid(calc_pout_fp_vld[57])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10432" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_58 (
    .in_data(calc_op0_fp_58_d1),
    .in_op(calc_op1_fp_58_d1),
    .in_op_valid(calc_op1_vld_fp_d1[58]),
    .in_sel(calc_dlv_en_fp_d1[58]),
    .in_valid(calc_op_en_fp_d1[58]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_58_sum),
    .out_final_valid(calc_fout_fp_vld[58]),
    .out_partial_data(calc_pout_fp_58_sum),
    .out_partial_valid(calc_pout_fp_vld[58])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10445" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_59 (
    .in_data(calc_op0_fp_59_d1),
    .in_op(calc_op1_fp_59_d1),
    .in_op_valid(calc_op1_vld_fp_d1[59]),
    .in_sel(calc_dlv_en_fp_d1[59]),
    .in_valid(calc_op_en_fp_d1[59]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_59_sum),
    .out_final_valid(calc_fout_fp_vld[59]),
    .out_partial_data(calc_pout_fp_59_sum),
    .out_partial_valid(calc_pout_fp_vld[59])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9756" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_6 (
    .in_data(calc_op0_fp_6_d1),
    .in_op(calc_op1_fp_6_d1),
    .in_op_valid(calc_op1_vld_fp_d1[6]),
    .in_sel(calc_dlv_en_fp_d1[6]),
    .in_valid(calc_op_en_fp_d1[6]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_6_sum),
    .out_final_valid(calc_fout_fp_vld[6]),
    .out_partial_data(calc_pout_fp_6_sum),
    .out_partial_valid(calc_pout_fp_vld[6])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10458" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_60 (
    .in_data(calc_op0_fp_60_d1),
    .in_op(calc_op1_fp_60_d1),
    .in_op_valid(calc_op1_vld_fp_d1[60]),
    .in_sel(calc_dlv_en_fp_d1[60]),
    .in_valid(calc_op_en_fp_d1[60]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_60_sum),
    .out_final_valid(calc_fout_fp_vld[60]),
    .out_partial_data(calc_pout_fp_60_sum),
    .out_partial_valid(calc_pout_fp_vld[60])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10471" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_61 (
    .in_data(calc_op0_fp_61_d1),
    .in_op(calc_op1_fp_61_d1),
    .in_op_valid(calc_op1_vld_fp_d1[61]),
    .in_sel(calc_dlv_en_fp_d1[61]),
    .in_valid(calc_op_en_fp_d1[61]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_61_sum),
    .out_final_valid(calc_fout_fp_vld[61]),
    .out_partial_data(calc_pout_fp_61_sum),
    .out_partial_valid(calc_pout_fp_vld[61])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10484" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_62 (
    .in_data(calc_op0_fp_62_d1),
    .in_op(calc_op1_fp_62_d1),
    .in_op_valid(calc_op1_vld_fp_d1[62]),
    .in_sel(calc_dlv_en_fp_d1[62]),
    .in_valid(calc_op_en_fp_d1[62]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_62_sum),
    .out_final_valid(calc_fout_fp_vld[62]),
    .out_partial_data(calc_pout_fp_62_sum),
    .out_partial_valid(calc_pout_fp_vld[62])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:10497" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_63 (
    .in_data(calc_op0_fp_63_d1),
    .in_op(calc_op1_fp_63_d1),
    .in_op_valid(calc_op1_vld_fp_d1[63]),
    .in_sel(calc_dlv_en_fp_d1[63]),
    .in_valid(calc_op_en_fp_d1[63]),
    .nvdla_core_clk(nvdla_cell_clk_3),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_63_sum),
    .out_final_valid(calc_fout_fp_vld[63]),
    .out_partial_data(calc_pout_fp_63_sum),
    .out_partial_valid(calc_pout_fp_vld[63])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9769" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_7 (
    .in_data(calc_op0_fp_7_d1),
    .in_op(calc_op1_fp_7_d1),
    .in_op_valid(calc_op1_vld_fp_d1[7]),
    .in_sel(calc_dlv_en_fp_d1[7]),
    .in_valid(calc_op_en_fp_d1[7]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_7_sum),
    .out_final_valid(calc_fout_fp_vld[7]),
    .out_partial_data(calc_pout_fp_7_sum),
    .out_partial_valid(calc_pout_fp_vld[7])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9782" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_8 (
    .in_data(calc_op0_fp_8_d1),
    .in_op(calc_op1_fp_8_d1),
    .in_op_valid(calc_op1_vld_fp_d1[8]),
    .in_sel(calc_dlv_en_fp_d1[8]),
    .in_valid(calc_op_en_fp_d1[8]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_8_sum),
    .out_final_valid(calc_fout_fp_vld[8]),
    .out_partial_data(calc_pout_fp_8_sum),
    .out_partial_valid(calc_pout_fp_vld[8])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9795" *)
  NV_NVDLA_CACC_CALC_fp_48b u_cell_fp_9 (
    .in_data(calc_op0_fp_9_d1),
    .in_op(calc_op1_fp_9_d1),
    .in_op_valid(calc_op1_vld_fp_d1[9]),
    .in_sel(calc_dlv_en_fp_d1[9]),
    .in_valid(calc_op_en_fp_d1[9]),
    .nvdla_core_clk(nvdla_cell_clk_2),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_fp_9_sum),
    .out_final_valid(calc_fout_fp_vld[9]),
    .out_partial_data(calc_pout_fp_9_sum),
    .out_partial_valid(calc_pout_fp_vld[9])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7758" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_0 (
    .cfg_truncate(cfg_truncate[4:0]),
    .in_data(calc_op0_int_0_d1),
    .in_op(calc_op1_int_0_d1),
    .in_op_valid(calc_op1_vld_int_d1[0]),
    .in_sel(calc_dlv_en_int_d1[0]),
    .in_valid(calc_op_en_int_d1[0]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_0_sum),
    .out_final_sat(calc_fout_int_sat[0]),
    .out_final_valid(calc_fout_int_vld[0]),
    .out_partial_data(calc_pout_int_0_sum),
    .out_partial_valid(calc_pout_int_vld[0])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7773" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_1 (
    .cfg_truncate(cfg_truncate[9:5]),
    .in_data(calc_op0_int_1_d1),
    .in_op(calc_op1_int_1_d1),
    .in_op_valid(calc_op1_vld_int_d1[1]),
    .in_sel(calc_dlv_en_int_d1[1]),
    .in_valid(calc_op_en_int_d1[1]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_1_sum),
    .out_final_sat(calc_fout_int_sat[1]),
    .out_final_valid(calc_fout_int_vld[1]),
    .out_partial_data(calc_pout_int_1_sum),
    .out_partial_valid(calc_pout_int_vld[1])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7908" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_10 (
    .cfg_truncate(cfg_truncate[54:50]),
    .in_data(calc_op0_int_10_d1),
    .in_op(calc_op1_int_10_d1),
    .in_op_valid(calc_op1_vld_int_d1[10]),
    .in_sel(calc_dlv_en_int_d1[10]),
    .in_valid(calc_op_en_int_d1[10]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_10_sum),
    .out_final_sat(calc_fout_int_sat[10]),
    .out_final_valid(calc_fout_int_vld[10]),
    .out_partial_data(calc_pout_int_10_sum),
    .out_partial_valid(calc_pout_int_vld[10])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9258" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_100 (
    .cfg_truncate(cfg_truncate[504:500]),
    .in_data(calc_op0_int_100_d1),
    .in_op(calc_op1_int_100_d1),
    .in_op_valid(calc_op1_vld_int_d1[100]),
    .in_sel(calc_dlv_en_int_d1[100]),
    .in_valid(calc_op_en_int_d1[100]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_100_sum),
    .out_final_sat(calc_fout_int_sat[100]),
    .out_final_valid(calc_fout_int_vld[100]),
    .out_partial_data(calc_pout_int_100_sum),
    .out_partial_valid(calc_pout_int_vld[100])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9273" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_101 (
    .cfg_truncate(cfg_truncate[509:505]),
    .in_data(calc_op0_int_101_d1),
    .in_op(calc_op1_int_101_d1),
    .in_op_valid(calc_op1_vld_int_d1[101]),
    .in_sel(calc_dlv_en_int_d1[101]),
    .in_valid(calc_op_en_int_d1[101]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_101_sum),
    .out_final_sat(calc_fout_int_sat[101]),
    .out_final_valid(calc_fout_int_vld[101]),
    .out_partial_data(calc_pout_int_101_sum),
    .out_partial_valid(calc_pout_int_vld[101])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9288" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_102 (
    .cfg_truncate(cfg_truncate[514:510]),
    .in_data(calc_op0_int_102_d1),
    .in_op(calc_op1_int_102_d1),
    .in_op_valid(calc_op1_vld_int_d1[102]),
    .in_sel(calc_dlv_en_int_d1[102]),
    .in_valid(calc_op_en_int_d1[102]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_102_sum),
    .out_final_sat(calc_fout_int_sat[102]),
    .out_final_valid(calc_fout_int_vld[102]),
    .out_partial_data(calc_pout_int_102_sum),
    .out_partial_valid(calc_pout_int_vld[102])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9303" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_103 (
    .cfg_truncate(cfg_truncate[519:515]),
    .in_data(calc_op0_int_103_d1),
    .in_op(calc_op1_int_103_d1),
    .in_op_valid(calc_op1_vld_int_d1[103]),
    .in_sel(calc_dlv_en_int_d1[103]),
    .in_valid(calc_op_en_int_d1[103]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_103_sum),
    .out_final_sat(calc_fout_int_sat[103]),
    .out_final_valid(calc_fout_int_vld[103]),
    .out_partial_data(calc_pout_int_103_sum),
    .out_partial_valid(calc_pout_int_vld[103])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9318" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_104 (
    .cfg_truncate(cfg_truncate[524:520]),
    .in_data(calc_op0_int_104_d1),
    .in_op(calc_op1_int_104_d1),
    .in_op_valid(calc_op1_vld_int_d1[104]),
    .in_sel(calc_dlv_en_int_d1[104]),
    .in_valid(calc_op_en_int_d1[104]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_104_sum),
    .out_final_sat(calc_fout_int_sat[104]),
    .out_final_valid(calc_fout_int_vld[104]),
    .out_partial_data(calc_pout_int_104_sum),
    .out_partial_valid(calc_pout_int_vld[104])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9333" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_105 (
    .cfg_truncate(cfg_truncate[529:525]),
    .in_data(calc_op0_int_105_d1),
    .in_op(calc_op1_int_105_d1),
    .in_op_valid(calc_op1_vld_int_d1[105]),
    .in_sel(calc_dlv_en_int_d1[105]),
    .in_valid(calc_op_en_int_d1[105]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_105_sum),
    .out_final_sat(calc_fout_int_sat[105]),
    .out_final_valid(calc_fout_int_vld[105]),
    .out_partial_data(calc_pout_int_105_sum),
    .out_partial_valid(calc_pout_int_vld[105])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9348" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_106 (
    .cfg_truncate(cfg_truncate[534:530]),
    .in_data(calc_op0_int_106_d1),
    .in_op(calc_op1_int_106_d1),
    .in_op_valid(calc_op1_vld_int_d1[106]),
    .in_sel(calc_dlv_en_int_d1[106]),
    .in_valid(calc_op_en_int_d1[106]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_106_sum),
    .out_final_sat(calc_fout_int_sat[106]),
    .out_final_valid(calc_fout_int_vld[106]),
    .out_partial_data(calc_pout_int_106_sum),
    .out_partial_valid(calc_pout_int_vld[106])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9363" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_107 (
    .cfg_truncate(cfg_truncate[539:535]),
    .in_data(calc_op0_int_107_d1),
    .in_op(calc_op1_int_107_d1),
    .in_op_valid(calc_op1_vld_int_d1[107]),
    .in_sel(calc_dlv_en_int_d1[107]),
    .in_valid(calc_op_en_int_d1[107]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_107_sum),
    .out_final_sat(calc_fout_int_sat[107]),
    .out_final_valid(calc_fout_int_vld[107]),
    .out_partial_data(calc_pout_int_107_sum),
    .out_partial_valid(calc_pout_int_vld[107])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9378" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_108 (
    .cfg_truncate(cfg_truncate[544:540]),
    .in_data(calc_op0_int_108_d1),
    .in_op(calc_op1_int_108_d1),
    .in_op_valid(calc_op1_vld_int_d1[108]),
    .in_sel(calc_dlv_en_int_d1[108]),
    .in_valid(calc_op_en_int_d1[108]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_108_sum),
    .out_final_sat(calc_fout_int_sat[108]),
    .out_final_valid(calc_fout_int_vld[108]),
    .out_partial_data(calc_pout_int_108_sum),
    .out_partial_valid(calc_pout_int_vld[108])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9393" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_109 (
    .cfg_truncate(cfg_truncate[549:545]),
    .in_data(calc_op0_int_109_d1),
    .in_op(calc_op1_int_109_d1),
    .in_op_valid(calc_op1_vld_int_d1[109]),
    .in_sel(calc_dlv_en_int_d1[109]),
    .in_valid(calc_op_en_int_d1[109]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_109_sum),
    .out_final_sat(calc_fout_int_sat[109]),
    .out_final_valid(calc_fout_int_vld[109]),
    .out_partial_data(calc_pout_int_109_sum),
    .out_partial_valid(calc_pout_int_vld[109])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7923" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_11 (
    .cfg_truncate(cfg_truncate[59:55]),
    .in_data(calc_op0_int_11_d1),
    .in_op(calc_op1_int_11_d1),
    .in_op_valid(calc_op1_vld_int_d1[11]),
    .in_sel(calc_dlv_en_int_d1[11]),
    .in_valid(calc_op_en_int_d1[11]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_11_sum),
    .out_final_sat(calc_fout_int_sat[11]),
    .out_final_valid(calc_fout_int_vld[11]),
    .out_partial_data(calc_pout_int_11_sum),
    .out_partial_valid(calc_pout_int_vld[11])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9408" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_110 (
    .cfg_truncate(cfg_truncate[554:550]),
    .in_data(calc_op0_int_110_d1),
    .in_op(calc_op1_int_110_d1),
    .in_op_valid(calc_op1_vld_int_d1[110]),
    .in_sel(calc_dlv_en_int_d1[110]),
    .in_valid(calc_op_en_int_d1[110]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_110_sum),
    .out_final_sat(calc_fout_int_sat[110]),
    .out_final_valid(calc_fout_int_vld[110]),
    .out_partial_data(calc_pout_int_110_sum),
    .out_partial_valid(calc_pout_int_vld[110])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9423" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_111 (
    .cfg_truncate(cfg_truncate[559:555]),
    .in_data(calc_op0_int_111_d1),
    .in_op(calc_op1_int_111_d1),
    .in_op_valid(calc_op1_vld_int_d1[111]),
    .in_sel(calc_dlv_en_int_d1[111]),
    .in_valid(calc_op_en_int_d1[111]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_111_sum),
    .out_final_sat(calc_fout_int_sat[111]),
    .out_final_valid(calc_fout_int_vld[111]),
    .out_partial_data(calc_pout_int_111_sum),
    .out_partial_valid(calc_pout_int_vld[111])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9438" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_112 (
    .cfg_truncate(cfg_truncate[564:560]),
    .in_data(calc_op0_int_112_d1),
    .in_op(calc_op1_int_112_d1),
    .in_op_valid(calc_op1_vld_int_d1[112]),
    .in_sel(calc_dlv_en_int_d1[112]),
    .in_valid(calc_op_en_int_d1[112]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_112_sum),
    .out_final_sat(calc_fout_int_sat[112]),
    .out_final_valid(calc_fout_int_vld[112]),
    .out_partial_data(calc_pout_int_112_sum),
    .out_partial_valid(calc_pout_int_vld[112])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9453" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_113 (
    .cfg_truncate(cfg_truncate[569:565]),
    .in_data(calc_op0_int_113_d1),
    .in_op(calc_op1_int_113_d1),
    .in_op_valid(calc_op1_vld_int_d1[113]),
    .in_sel(calc_dlv_en_int_d1[113]),
    .in_valid(calc_op_en_int_d1[113]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_113_sum),
    .out_final_sat(calc_fout_int_sat[113]),
    .out_final_valid(calc_fout_int_vld[113]),
    .out_partial_data(calc_pout_int_113_sum),
    .out_partial_valid(calc_pout_int_vld[113])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9468" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_114 (
    .cfg_truncate(cfg_truncate[574:570]),
    .in_data(calc_op0_int_114_d1),
    .in_op(calc_op1_int_114_d1),
    .in_op_valid(calc_op1_vld_int_d1[114]),
    .in_sel(calc_dlv_en_int_d1[114]),
    .in_valid(calc_op_en_int_d1[114]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_114_sum),
    .out_final_sat(calc_fout_int_sat[114]),
    .out_final_valid(calc_fout_int_vld[114]),
    .out_partial_data(calc_pout_int_114_sum),
    .out_partial_valid(calc_pout_int_vld[114])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9483" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_115 (
    .cfg_truncate(cfg_truncate[579:575]),
    .in_data(calc_op0_int_115_d1),
    .in_op(calc_op1_int_115_d1),
    .in_op_valid(calc_op1_vld_int_d1[115]),
    .in_sel(calc_dlv_en_int_d1[115]),
    .in_valid(calc_op_en_int_d1[115]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_115_sum),
    .out_final_sat(calc_fout_int_sat[115]),
    .out_final_valid(calc_fout_int_vld[115]),
    .out_partial_data(calc_pout_int_115_sum),
    .out_partial_valid(calc_pout_int_vld[115])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9498" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_116 (
    .cfg_truncate(cfg_truncate[584:580]),
    .in_data(calc_op0_int_116_d1),
    .in_op(calc_op1_int_116_d1),
    .in_op_valid(calc_op1_vld_int_d1[116]),
    .in_sel(calc_dlv_en_int_d1[116]),
    .in_valid(calc_op_en_int_d1[116]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_116_sum),
    .out_final_sat(calc_fout_int_sat[116]),
    .out_final_valid(calc_fout_int_vld[116]),
    .out_partial_data(calc_pout_int_116_sum),
    .out_partial_valid(calc_pout_int_vld[116])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9513" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_117 (
    .cfg_truncate(cfg_truncate[589:585]),
    .in_data(calc_op0_int_117_d1),
    .in_op(calc_op1_int_117_d1),
    .in_op_valid(calc_op1_vld_int_d1[117]),
    .in_sel(calc_dlv_en_int_d1[117]),
    .in_valid(calc_op_en_int_d1[117]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_117_sum),
    .out_final_sat(calc_fout_int_sat[117]),
    .out_final_valid(calc_fout_int_vld[117]),
    .out_partial_data(calc_pout_int_117_sum),
    .out_partial_valid(calc_pout_int_vld[117])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9528" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_118 (
    .cfg_truncate(cfg_truncate[594:590]),
    .in_data(calc_op0_int_118_d1),
    .in_op(calc_op1_int_118_d1),
    .in_op_valid(calc_op1_vld_int_d1[118]),
    .in_sel(calc_dlv_en_int_d1[118]),
    .in_valid(calc_op_en_int_d1[118]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_118_sum),
    .out_final_sat(calc_fout_int_sat[118]),
    .out_final_valid(calc_fout_int_vld[118]),
    .out_partial_data(calc_pout_int_118_sum),
    .out_partial_valid(calc_pout_int_vld[118])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9543" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_119 (
    .cfg_truncate(cfg_truncate[599:595]),
    .in_data(calc_op0_int_119_d1),
    .in_op(calc_op1_int_119_d1),
    .in_op_valid(calc_op1_vld_int_d1[119]),
    .in_sel(calc_dlv_en_int_d1[119]),
    .in_valid(calc_op_en_int_d1[119]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_119_sum),
    .out_final_sat(calc_fout_int_sat[119]),
    .out_final_valid(calc_fout_int_vld[119]),
    .out_partial_data(calc_pout_int_119_sum),
    .out_partial_valid(calc_pout_int_vld[119])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7938" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_12 (
    .cfg_truncate(cfg_truncate[64:60]),
    .in_data(calc_op0_int_12_d1),
    .in_op(calc_op1_int_12_d1),
    .in_op_valid(calc_op1_vld_int_d1[12]),
    .in_sel(calc_dlv_en_int_d1[12]),
    .in_valid(calc_op_en_int_d1[12]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_12_sum),
    .out_final_sat(calc_fout_int_sat[12]),
    .out_final_valid(calc_fout_int_vld[12]),
    .out_partial_data(calc_pout_int_12_sum),
    .out_partial_valid(calc_pout_int_vld[12])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9558" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_120 (
    .cfg_truncate(cfg_truncate[604:600]),
    .in_data(calc_op0_int_120_d1),
    .in_op(calc_op1_int_120_d1),
    .in_op_valid(calc_op1_vld_int_d1[120]),
    .in_sel(calc_dlv_en_int_d1[120]),
    .in_valid(calc_op_en_int_d1[120]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_120_sum),
    .out_final_sat(calc_fout_int_sat[120]),
    .out_final_valid(calc_fout_int_vld[120]),
    .out_partial_data(calc_pout_int_120_sum),
    .out_partial_valid(calc_pout_int_vld[120])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9573" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_121 (
    .cfg_truncate(cfg_truncate[609:605]),
    .in_data(calc_op0_int_121_d1),
    .in_op(calc_op1_int_121_d1),
    .in_op_valid(calc_op1_vld_int_d1[121]),
    .in_sel(calc_dlv_en_int_d1[121]),
    .in_valid(calc_op_en_int_d1[121]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_121_sum),
    .out_final_sat(calc_fout_int_sat[121]),
    .out_final_valid(calc_fout_int_vld[121]),
    .out_partial_data(calc_pout_int_121_sum),
    .out_partial_valid(calc_pout_int_vld[121])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9588" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_122 (
    .cfg_truncate(cfg_truncate[614:610]),
    .in_data(calc_op0_int_122_d1),
    .in_op(calc_op1_int_122_d1),
    .in_op_valid(calc_op1_vld_int_d1[122]),
    .in_sel(calc_dlv_en_int_d1[122]),
    .in_valid(calc_op_en_int_d1[122]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_122_sum),
    .out_final_sat(calc_fout_int_sat[122]),
    .out_final_valid(calc_fout_int_vld[122]),
    .out_partial_data(calc_pout_int_122_sum),
    .out_partial_valid(calc_pout_int_vld[122])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9603" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_123 (
    .cfg_truncate(cfg_truncate[619:615]),
    .in_data(calc_op0_int_123_d1),
    .in_op(calc_op1_int_123_d1),
    .in_op_valid(calc_op1_vld_int_d1[123]),
    .in_sel(calc_dlv_en_int_d1[123]),
    .in_valid(calc_op_en_int_d1[123]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_123_sum),
    .out_final_sat(calc_fout_int_sat[123]),
    .out_final_valid(calc_fout_int_vld[123]),
    .out_partial_data(calc_pout_int_123_sum),
    .out_partial_valid(calc_pout_int_vld[123])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9618" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_124 (
    .cfg_truncate(cfg_truncate[624:620]),
    .in_data(calc_op0_int_124_d1),
    .in_op(calc_op1_int_124_d1),
    .in_op_valid(calc_op1_vld_int_d1[124]),
    .in_sel(calc_dlv_en_int_d1[124]),
    .in_valid(calc_op_en_int_d1[124]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_124_sum),
    .out_final_sat(calc_fout_int_sat[124]),
    .out_final_valid(calc_fout_int_vld[124]),
    .out_partial_data(calc_pout_int_124_sum),
    .out_partial_valid(calc_pout_int_vld[124])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9633" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_125 (
    .cfg_truncate(cfg_truncate[629:625]),
    .in_data(calc_op0_int_125_d1),
    .in_op(calc_op1_int_125_d1),
    .in_op_valid(calc_op1_vld_int_d1[125]),
    .in_sel(calc_dlv_en_int_d1[125]),
    .in_valid(calc_op_en_int_d1[125]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_125_sum),
    .out_final_sat(calc_fout_int_sat[125]),
    .out_final_valid(calc_fout_int_vld[125]),
    .out_partial_data(calc_pout_int_125_sum),
    .out_partial_valid(calc_pout_int_vld[125])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9648" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_126 (
    .cfg_truncate(cfg_truncate[634:630]),
    .in_data(calc_op0_int_126_d1),
    .in_op(calc_op1_int_126_d1),
    .in_op_valid(calc_op1_vld_int_d1[126]),
    .in_sel(calc_dlv_en_int_d1[126]),
    .in_valid(calc_op_en_int_d1[126]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_126_sum),
    .out_final_sat(calc_fout_int_sat[126]),
    .out_final_valid(calc_fout_int_vld[126]),
    .out_partial_data(calc_pout_int_126_sum),
    .out_partial_valid(calc_pout_int_vld[126])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9663" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_127 (
    .cfg_truncate(cfg_truncate[639:635]),
    .in_data(calc_op0_int_127_d1),
    .in_op(calc_op1_int_127_d1),
    .in_op_valid(calc_op1_vld_int_d1[127]),
    .in_sel(calc_dlv_en_int_d1[127]),
    .in_valid(calc_op_en_int_d1[127]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_127_sum),
    .out_final_sat(calc_fout_int_sat[127]),
    .out_final_valid(calc_fout_int_vld[127]),
    .out_partial_data(calc_pout_int_127_sum),
    .out_partial_valid(calc_pout_int_vld[127])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7953" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_13 (
    .cfg_truncate(cfg_truncate[69:65]),
    .in_data(calc_op0_int_13_d1),
    .in_op(calc_op1_int_13_d1),
    .in_op_valid(calc_op1_vld_int_d1[13]),
    .in_sel(calc_dlv_en_int_d1[13]),
    .in_valid(calc_op_en_int_d1[13]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_13_sum),
    .out_final_sat(calc_fout_int_sat[13]),
    .out_final_valid(calc_fout_int_vld[13]),
    .out_partial_data(calc_pout_int_13_sum),
    .out_partial_valid(calc_pout_int_vld[13])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7968" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_14 (
    .cfg_truncate(cfg_truncate[74:70]),
    .in_data(calc_op0_int_14_d1),
    .in_op(calc_op1_int_14_d1),
    .in_op_valid(calc_op1_vld_int_d1[14]),
    .in_sel(calc_dlv_en_int_d1[14]),
    .in_valid(calc_op_en_int_d1[14]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_14_sum),
    .out_final_sat(calc_fout_int_sat[14]),
    .out_final_valid(calc_fout_int_vld[14]),
    .out_partial_data(calc_pout_int_14_sum),
    .out_partial_valid(calc_pout_int_vld[14])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7983" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_15 (
    .cfg_truncate(cfg_truncate[79:75]),
    .in_data(calc_op0_int_15_d1),
    .in_op(calc_op1_int_15_d1),
    .in_op_valid(calc_op1_vld_int_d1[15]),
    .in_sel(calc_dlv_en_int_d1[15]),
    .in_valid(calc_op_en_int_d1[15]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_15_sum),
    .out_final_sat(calc_fout_int_sat[15]),
    .out_final_valid(calc_fout_int_vld[15]),
    .out_partial_data(calc_pout_int_15_sum),
    .out_partial_valid(calc_pout_int_vld[15])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7998" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_16 (
    .cfg_truncate(cfg_truncate[84:80]),
    .in_data(calc_op0_int_16_d1),
    .in_op(calc_op1_int_16_d1),
    .in_op_valid(calc_op1_vld_int_d1[16]),
    .in_sel(calc_dlv_en_int_d1[16]),
    .in_valid(calc_op_en_int_d1[16]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_16_sum),
    .out_final_sat(calc_fout_int_sat[16]),
    .out_final_valid(calc_fout_int_vld[16]),
    .out_partial_data(calc_pout_int_16_sum),
    .out_partial_valid(calc_pout_int_vld[16])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8013" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_17 (
    .cfg_truncate(cfg_truncate[89:85]),
    .in_data(calc_op0_int_17_d1),
    .in_op(calc_op1_int_17_d1),
    .in_op_valid(calc_op1_vld_int_d1[17]),
    .in_sel(calc_dlv_en_int_d1[17]),
    .in_valid(calc_op_en_int_d1[17]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_17_sum),
    .out_final_sat(calc_fout_int_sat[17]),
    .out_final_valid(calc_fout_int_vld[17]),
    .out_partial_data(calc_pout_int_17_sum),
    .out_partial_valid(calc_pout_int_vld[17])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8028" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_18 (
    .cfg_truncate(cfg_truncate[94:90]),
    .in_data(calc_op0_int_18_d1),
    .in_op(calc_op1_int_18_d1),
    .in_op_valid(calc_op1_vld_int_d1[18]),
    .in_sel(calc_dlv_en_int_d1[18]),
    .in_valid(calc_op_en_int_d1[18]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_18_sum),
    .out_final_sat(calc_fout_int_sat[18]),
    .out_final_valid(calc_fout_int_vld[18]),
    .out_partial_data(calc_pout_int_18_sum),
    .out_partial_valid(calc_pout_int_vld[18])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8043" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_19 (
    .cfg_truncate(cfg_truncate[99:95]),
    .in_data(calc_op0_int_19_d1),
    .in_op(calc_op1_int_19_d1),
    .in_op_valid(calc_op1_vld_int_d1[19]),
    .in_sel(calc_dlv_en_int_d1[19]),
    .in_valid(calc_op_en_int_d1[19]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_19_sum),
    .out_final_sat(calc_fout_int_sat[19]),
    .out_final_valid(calc_fout_int_vld[19]),
    .out_partial_data(calc_pout_int_19_sum),
    .out_partial_valid(calc_pout_int_vld[19])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7788" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_2 (
    .cfg_truncate(cfg_truncate[14:10]),
    .in_data(calc_op0_int_2_d1),
    .in_op(calc_op1_int_2_d1),
    .in_op_valid(calc_op1_vld_int_d1[2]),
    .in_sel(calc_dlv_en_int_d1[2]),
    .in_valid(calc_op_en_int_d1[2]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_2_sum),
    .out_final_sat(calc_fout_int_sat[2]),
    .out_final_valid(calc_fout_int_vld[2]),
    .out_partial_data(calc_pout_int_2_sum),
    .out_partial_valid(calc_pout_int_vld[2])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8058" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_20 (
    .cfg_truncate(cfg_truncate[104:100]),
    .in_data(calc_op0_int_20_d1),
    .in_op(calc_op1_int_20_d1),
    .in_op_valid(calc_op1_vld_int_d1[20]),
    .in_sel(calc_dlv_en_int_d1[20]),
    .in_valid(calc_op_en_int_d1[20]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_20_sum),
    .out_final_sat(calc_fout_int_sat[20]),
    .out_final_valid(calc_fout_int_vld[20]),
    .out_partial_data(calc_pout_int_20_sum),
    .out_partial_valid(calc_pout_int_vld[20])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8073" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_21 (
    .cfg_truncate(cfg_truncate[109:105]),
    .in_data(calc_op0_int_21_d1),
    .in_op(calc_op1_int_21_d1),
    .in_op_valid(calc_op1_vld_int_d1[21]),
    .in_sel(calc_dlv_en_int_d1[21]),
    .in_valid(calc_op_en_int_d1[21]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_21_sum),
    .out_final_sat(calc_fout_int_sat[21]),
    .out_final_valid(calc_fout_int_vld[21]),
    .out_partial_data(calc_pout_int_21_sum),
    .out_partial_valid(calc_pout_int_vld[21])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8088" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_22 (
    .cfg_truncate(cfg_truncate[114:110]),
    .in_data(calc_op0_int_22_d1),
    .in_op(calc_op1_int_22_d1),
    .in_op_valid(calc_op1_vld_int_d1[22]),
    .in_sel(calc_dlv_en_int_d1[22]),
    .in_valid(calc_op_en_int_d1[22]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_22_sum),
    .out_final_sat(calc_fout_int_sat[22]),
    .out_final_valid(calc_fout_int_vld[22]),
    .out_partial_data(calc_pout_int_22_sum),
    .out_partial_valid(calc_pout_int_vld[22])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8103" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_23 (
    .cfg_truncate(cfg_truncate[119:115]),
    .in_data(calc_op0_int_23_d1),
    .in_op(calc_op1_int_23_d1),
    .in_op_valid(calc_op1_vld_int_d1[23]),
    .in_sel(calc_dlv_en_int_d1[23]),
    .in_valid(calc_op_en_int_d1[23]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_23_sum),
    .out_final_sat(calc_fout_int_sat[23]),
    .out_final_valid(calc_fout_int_vld[23]),
    .out_partial_data(calc_pout_int_23_sum),
    .out_partial_valid(calc_pout_int_vld[23])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8118" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_24 (
    .cfg_truncate(cfg_truncate[124:120]),
    .in_data(calc_op0_int_24_d1),
    .in_op(calc_op1_int_24_d1),
    .in_op_valid(calc_op1_vld_int_d1[24]),
    .in_sel(calc_dlv_en_int_d1[24]),
    .in_valid(calc_op_en_int_d1[24]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_24_sum),
    .out_final_sat(calc_fout_int_sat[24]),
    .out_final_valid(calc_fout_int_vld[24]),
    .out_partial_data(calc_pout_int_24_sum),
    .out_partial_valid(calc_pout_int_vld[24])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8133" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_25 (
    .cfg_truncate(cfg_truncate[129:125]),
    .in_data(calc_op0_int_25_d1),
    .in_op(calc_op1_int_25_d1),
    .in_op_valid(calc_op1_vld_int_d1[25]),
    .in_sel(calc_dlv_en_int_d1[25]),
    .in_valid(calc_op_en_int_d1[25]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_25_sum),
    .out_final_sat(calc_fout_int_sat[25]),
    .out_final_valid(calc_fout_int_vld[25]),
    .out_partial_data(calc_pout_int_25_sum),
    .out_partial_valid(calc_pout_int_vld[25])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8148" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_26 (
    .cfg_truncate(cfg_truncate[134:130]),
    .in_data(calc_op0_int_26_d1),
    .in_op(calc_op1_int_26_d1),
    .in_op_valid(calc_op1_vld_int_d1[26]),
    .in_sel(calc_dlv_en_int_d1[26]),
    .in_valid(calc_op_en_int_d1[26]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_26_sum),
    .out_final_sat(calc_fout_int_sat[26]),
    .out_final_valid(calc_fout_int_vld[26]),
    .out_partial_data(calc_pout_int_26_sum),
    .out_partial_valid(calc_pout_int_vld[26])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8163" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_27 (
    .cfg_truncate(cfg_truncate[139:135]),
    .in_data(calc_op0_int_27_d1),
    .in_op(calc_op1_int_27_d1),
    .in_op_valid(calc_op1_vld_int_d1[27]),
    .in_sel(calc_dlv_en_int_d1[27]),
    .in_valid(calc_op_en_int_d1[27]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_27_sum),
    .out_final_sat(calc_fout_int_sat[27]),
    .out_final_valid(calc_fout_int_vld[27]),
    .out_partial_data(calc_pout_int_27_sum),
    .out_partial_valid(calc_pout_int_vld[27])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8178" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_28 (
    .cfg_truncate(cfg_truncate[144:140]),
    .in_data(calc_op0_int_28_d1),
    .in_op(calc_op1_int_28_d1),
    .in_op_valid(calc_op1_vld_int_d1[28]),
    .in_sel(calc_dlv_en_int_d1[28]),
    .in_valid(calc_op_en_int_d1[28]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_28_sum),
    .out_final_sat(calc_fout_int_sat[28]),
    .out_final_valid(calc_fout_int_vld[28]),
    .out_partial_data(calc_pout_int_28_sum),
    .out_partial_valid(calc_pout_int_vld[28])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8193" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_29 (
    .cfg_truncate(cfg_truncate[149:145]),
    .in_data(calc_op0_int_29_d1),
    .in_op(calc_op1_int_29_d1),
    .in_op_valid(calc_op1_vld_int_d1[29]),
    .in_sel(calc_dlv_en_int_d1[29]),
    .in_valid(calc_op_en_int_d1[29]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_29_sum),
    .out_final_sat(calc_fout_int_sat[29]),
    .out_final_valid(calc_fout_int_vld[29]),
    .out_partial_data(calc_pout_int_29_sum),
    .out_partial_valid(calc_pout_int_vld[29])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7803" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_3 (
    .cfg_truncate(cfg_truncate[19:15]),
    .in_data(calc_op0_int_3_d1),
    .in_op(calc_op1_int_3_d1),
    .in_op_valid(calc_op1_vld_int_d1[3]),
    .in_sel(calc_dlv_en_int_d1[3]),
    .in_valid(calc_op_en_int_d1[3]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_3_sum),
    .out_final_sat(calc_fout_int_sat[3]),
    .out_final_valid(calc_fout_int_vld[3]),
    .out_partial_data(calc_pout_int_3_sum),
    .out_partial_valid(calc_pout_int_vld[3])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8208" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_30 (
    .cfg_truncate(cfg_truncate[154:150]),
    .in_data(calc_op0_int_30_d1),
    .in_op(calc_op1_int_30_d1),
    .in_op_valid(calc_op1_vld_int_d1[30]),
    .in_sel(calc_dlv_en_int_d1[30]),
    .in_valid(calc_op_en_int_d1[30]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_30_sum),
    .out_final_sat(calc_fout_int_sat[30]),
    .out_final_valid(calc_fout_int_vld[30]),
    .out_partial_data(calc_pout_int_30_sum),
    .out_partial_valid(calc_pout_int_vld[30])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8223" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_31 (
    .cfg_truncate(cfg_truncate[159:155]),
    .in_data(calc_op0_int_31_d1),
    .in_op(calc_op1_int_31_d1),
    .in_op_valid(calc_op1_vld_int_d1[31]),
    .in_sel(calc_dlv_en_int_d1[31]),
    .in_valid(calc_op_en_int_d1[31]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_31_sum),
    .out_final_sat(calc_fout_int_sat[31]),
    .out_final_valid(calc_fout_int_vld[31]),
    .out_partial_data(calc_pout_int_31_sum),
    .out_partial_valid(calc_pout_int_vld[31])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8238" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_32 (
    .cfg_truncate(cfg_truncate[164:160]),
    .in_data(calc_op0_int_32_d1),
    .in_op(calc_op1_int_32_d1),
    .in_op_valid(calc_op1_vld_int_d1[32]),
    .in_sel(calc_dlv_en_int_d1[32]),
    .in_valid(calc_op_en_int_d1[32]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_32_sum),
    .out_final_sat(calc_fout_int_sat[32]),
    .out_final_valid(calc_fout_int_vld[32]),
    .out_partial_data(calc_pout_int_32_sum),
    .out_partial_valid(calc_pout_int_vld[32])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8253" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_33 (
    .cfg_truncate(cfg_truncate[169:165]),
    .in_data(calc_op0_int_33_d1),
    .in_op(calc_op1_int_33_d1),
    .in_op_valid(calc_op1_vld_int_d1[33]),
    .in_sel(calc_dlv_en_int_d1[33]),
    .in_valid(calc_op_en_int_d1[33]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_33_sum),
    .out_final_sat(calc_fout_int_sat[33]),
    .out_final_valid(calc_fout_int_vld[33]),
    .out_partial_data(calc_pout_int_33_sum),
    .out_partial_valid(calc_pout_int_vld[33])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8268" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_34 (
    .cfg_truncate(cfg_truncate[174:170]),
    .in_data(calc_op0_int_34_d1),
    .in_op(calc_op1_int_34_d1),
    .in_op_valid(calc_op1_vld_int_d1[34]),
    .in_sel(calc_dlv_en_int_d1[34]),
    .in_valid(calc_op_en_int_d1[34]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_34_sum),
    .out_final_sat(calc_fout_int_sat[34]),
    .out_final_valid(calc_fout_int_vld[34]),
    .out_partial_data(calc_pout_int_34_sum),
    .out_partial_valid(calc_pout_int_vld[34])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8283" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_35 (
    .cfg_truncate(cfg_truncate[179:175]),
    .in_data(calc_op0_int_35_d1),
    .in_op(calc_op1_int_35_d1),
    .in_op_valid(calc_op1_vld_int_d1[35]),
    .in_sel(calc_dlv_en_int_d1[35]),
    .in_valid(calc_op_en_int_d1[35]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_35_sum),
    .out_final_sat(calc_fout_int_sat[35]),
    .out_final_valid(calc_fout_int_vld[35]),
    .out_partial_data(calc_pout_int_35_sum),
    .out_partial_valid(calc_pout_int_vld[35])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8298" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_36 (
    .cfg_truncate(cfg_truncate[184:180]),
    .in_data(calc_op0_int_36_d1),
    .in_op(calc_op1_int_36_d1),
    .in_op_valid(calc_op1_vld_int_d1[36]),
    .in_sel(calc_dlv_en_int_d1[36]),
    .in_valid(calc_op_en_int_d1[36]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_36_sum),
    .out_final_sat(calc_fout_int_sat[36]),
    .out_final_valid(calc_fout_int_vld[36]),
    .out_partial_data(calc_pout_int_36_sum),
    .out_partial_valid(calc_pout_int_vld[36])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8313" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_37 (
    .cfg_truncate(cfg_truncate[189:185]),
    .in_data(calc_op0_int_37_d1),
    .in_op(calc_op1_int_37_d1),
    .in_op_valid(calc_op1_vld_int_d1[37]),
    .in_sel(calc_dlv_en_int_d1[37]),
    .in_valid(calc_op_en_int_d1[37]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_37_sum),
    .out_final_sat(calc_fout_int_sat[37]),
    .out_final_valid(calc_fout_int_vld[37]),
    .out_partial_data(calc_pout_int_37_sum),
    .out_partial_valid(calc_pout_int_vld[37])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8328" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_38 (
    .cfg_truncate(cfg_truncate[194:190]),
    .in_data(calc_op0_int_38_d1),
    .in_op(calc_op1_int_38_d1),
    .in_op_valid(calc_op1_vld_int_d1[38]),
    .in_sel(calc_dlv_en_int_d1[38]),
    .in_valid(calc_op_en_int_d1[38]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_38_sum),
    .out_final_sat(calc_fout_int_sat[38]),
    .out_final_valid(calc_fout_int_vld[38]),
    .out_partial_data(calc_pout_int_38_sum),
    .out_partial_valid(calc_pout_int_vld[38])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8343" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_39 (
    .cfg_truncate(cfg_truncate[199:195]),
    .in_data(calc_op0_int_39_d1),
    .in_op(calc_op1_int_39_d1),
    .in_op_valid(calc_op1_vld_int_d1[39]),
    .in_sel(calc_dlv_en_int_d1[39]),
    .in_valid(calc_op_en_int_d1[39]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_39_sum),
    .out_final_sat(calc_fout_int_sat[39]),
    .out_final_valid(calc_fout_int_vld[39]),
    .out_partial_data(calc_pout_int_39_sum),
    .out_partial_valid(calc_pout_int_vld[39])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7818" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_4 (
    .cfg_truncate(cfg_truncate[24:20]),
    .in_data(calc_op0_int_4_d1),
    .in_op(calc_op1_int_4_d1),
    .in_op_valid(calc_op1_vld_int_d1[4]),
    .in_sel(calc_dlv_en_int_d1[4]),
    .in_valid(calc_op_en_int_d1[4]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_4_sum),
    .out_final_sat(calc_fout_int_sat[4]),
    .out_final_valid(calc_fout_int_vld[4]),
    .out_partial_data(calc_pout_int_4_sum),
    .out_partial_valid(calc_pout_int_vld[4])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8358" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_40 (
    .cfg_truncate(cfg_truncate[204:200]),
    .in_data(calc_op0_int_40_d1),
    .in_op(calc_op1_int_40_d1),
    .in_op_valid(calc_op1_vld_int_d1[40]),
    .in_sel(calc_dlv_en_int_d1[40]),
    .in_valid(calc_op_en_int_d1[40]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_40_sum),
    .out_final_sat(calc_fout_int_sat[40]),
    .out_final_valid(calc_fout_int_vld[40]),
    .out_partial_data(calc_pout_int_40_sum),
    .out_partial_valid(calc_pout_int_vld[40])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8373" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_41 (
    .cfg_truncate(cfg_truncate[209:205]),
    .in_data(calc_op0_int_41_d1),
    .in_op(calc_op1_int_41_d1),
    .in_op_valid(calc_op1_vld_int_d1[41]),
    .in_sel(calc_dlv_en_int_d1[41]),
    .in_valid(calc_op_en_int_d1[41]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_41_sum),
    .out_final_sat(calc_fout_int_sat[41]),
    .out_final_valid(calc_fout_int_vld[41]),
    .out_partial_data(calc_pout_int_41_sum),
    .out_partial_valid(calc_pout_int_vld[41])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8388" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_42 (
    .cfg_truncate(cfg_truncate[214:210]),
    .in_data(calc_op0_int_42_d1),
    .in_op(calc_op1_int_42_d1),
    .in_op_valid(calc_op1_vld_int_d1[42]),
    .in_sel(calc_dlv_en_int_d1[42]),
    .in_valid(calc_op_en_int_d1[42]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_42_sum),
    .out_final_sat(calc_fout_int_sat[42]),
    .out_final_valid(calc_fout_int_vld[42]),
    .out_partial_data(calc_pout_int_42_sum),
    .out_partial_valid(calc_pout_int_vld[42])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8403" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_43 (
    .cfg_truncate(cfg_truncate[219:215]),
    .in_data(calc_op0_int_43_d1),
    .in_op(calc_op1_int_43_d1),
    .in_op_valid(calc_op1_vld_int_d1[43]),
    .in_sel(calc_dlv_en_int_d1[43]),
    .in_valid(calc_op_en_int_d1[43]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_43_sum),
    .out_final_sat(calc_fout_int_sat[43]),
    .out_final_valid(calc_fout_int_vld[43]),
    .out_partial_data(calc_pout_int_43_sum),
    .out_partial_valid(calc_pout_int_vld[43])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8418" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_44 (
    .cfg_truncate(cfg_truncate[224:220]),
    .in_data(calc_op0_int_44_d1),
    .in_op(calc_op1_int_44_d1),
    .in_op_valid(calc_op1_vld_int_d1[44]),
    .in_sel(calc_dlv_en_int_d1[44]),
    .in_valid(calc_op_en_int_d1[44]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_44_sum),
    .out_final_sat(calc_fout_int_sat[44]),
    .out_final_valid(calc_fout_int_vld[44]),
    .out_partial_data(calc_pout_int_44_sum),
    .out_partial_valid(calc_pout_int_vld[44])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8433" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_45 (
    .cfg_truncate(cfg_truncate[229:225]),
    .in_data(calc_op0_int_45_d1),
    .in_op(calc_op1_int_45_d1),
    .in_op_valid(calc_op1_vld_int_d1[45]),
    .in_sel(calc_dlv_en_int_d1[45]),
    .in_valid(calc_op_en_int_d1[45]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_45_sum),
    .out_final_sat(calc_fout_int_sat[45]),
    .out_final_valid(calc_fout_int_vld[45]),
    .out_partial_data(calc_pout_int_45_sum),
    .out_partial_valid(calc_pout_int_vld[45])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8448" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_46 (
    .cfg_truncate(cfg_truncate[234:230]),
    .in_data(calc_op0_int_46_d1),
    .in_op(calc_op1_int_46_d1),
    .in_op_valid(calc_op1_vld_int_d1[46]),
    .in_sel(calc_dlv_en_int_d1[46]),
    .in_valid(calc_op_en_int_d1[46]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_46_sum),
    .out_final_sat(calc_fout_int_sat[46]),
    .out_final_valid(calc_fout_int_vld[46]),
    .out_partial_data(calc_pout_int_46_sum),
    .out_partial_valid(calc_pout_int_vld[46])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8463" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_47 (
    .cfg_truncate(cfg_truncate[239:235]),
    .in_data(calc_op0_int_47_d1),
    .in_op(calc_op1_int_47_d1),
    .in_op_valid(calc_op1_vld_int_d1[47]),
    .in_sel(calc_dlv_en_int_d1[47]),
    .in_valid(calc_op_en_int_d1[47]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_47_sum),
    .out_final_sat(calc_fout_int_sat[47]),
    .out_final_valid(calc_fout_int_vld[47]),
    .out_partial_data(calc_pout_int_47_sum),
    .out_partial_valid(calc_pout_int_vld[47])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8478" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_48 (
    .cfg_truncate(cfg_truncate[244:240]),
    .in_data(calc_op0_int_48_d1),
    .in_op(calc_op1_int_48_d1),
    .in_op_valid(calc_op1_vld_int_d1[48]),
    .in_sel(calc_dlv_en_int_d1[48]),
    .in_valid(calc_op_en_int_d1[48]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_48_sum),
    .out_final_sat(calc_fout_int_sat[48]),
    .out_final_valid(calc_fout_int_vld[48]),
    .out_partial_data(calc_pout_int_48_sum),
    .out_partial_valid(calc_pout_int_vld[48])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8493" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_49 (
    .cfg_truncate(cfg_truncate[249:245]),
    .in_data(calc_op0_int_49_d1),
    .in_op(calc_op1_int_49_d1),
    .in_op_valid(calc_op1_vld_int_d1[49]),
    .in_sel(calc_dlv_en_int_d1[49]),
    .in_valid(calc_op_en_int_d1[49]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_49_sum),
    .out_final_sat(calc_fout_int_sat[49]),
    .out_final_valid(calc_fout_int_vld[49]),
    .out_partial_data(calc_pout_int_49_sum),
    .out_partial_valid(calc_pout_int_vld[49])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7833" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_5 (
    .cfg_truncate(cfg_truncate[29:25]),
    .in_data(calc_op0_int_5_d1),
    .in_op(calc_op1_int_5_d1),
    .in_op_valid(calc_op1_vld_int_d1[5]),
    .in_sel(calc_dlv_en_int_d1[5]),
    .in_valid(calc_op_en_int_d1[5]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_5_sum),
    .out_final_sat(calc_fout_int_sat[5]),
    .out_final_valid(calc_fout_int_vld[5]),
    .out_partial_data(calc_pout_int_5_sum),
    .out_partial_valid(calc_pout_int_vld[5])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8508" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_50 (
    .cfg_truncate(cfg_truncate[254:250]),
    .in_data(calc_op0_int_50_d1),
    .in_op(calc_op1_int_50_d1),
    .in_op_valid(calc_op1_vld_int_d1[50]),
    .in_sel(calc_dlv_en_int_d1[50]),
    .in_valid(calc_op_en_int_d1[50]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_50_sum),
    .out_final_sat(calc_fout_int_sat[50]),
    .out_final_valid(calc_fout_int_vld[50]),
    .out_partial_data(calc_pout_int_50_sum),
    .out_partial_valid(calc_pout_int_vld[50])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8523" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_51 (
    .cfg_truncate(cfg_truncate[259:255]),
    .in_data(calc_op0_int_51_d1),
    .in_op(calc_op1_int_51_d1),
    .in_op_valid(calc_op1_vld_int_d1[51]),
    .in_sel(calc_dlv_en_int_d1[51]),
    .in_valid(calc_op_en_int_d1[51]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_51_sum),
    .out_final_sat(calc_fout_int_sat[51]),
    .out_final_valid(calc_fout_int_vld[51]),
    .out_partial_data(calc_pout_int_51_sum),
    .out_partial_valid(calc_pout_int_vld[51])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8538" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_52 (
    .cfg_truncate(cfg_truncate[264:260]),
    .in_data(calc_op0_int_52_d1),
    .in_op(calc_op1_int_52_d1),
    .in_op_valid(calc_op1_vld_int_d1[52]),
    .in_sel(calc_dlv_en_int_d1[52]),
    .in_valid(calc_op_en_int_d1[52]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_52_sum),
    .out_final_sat(calc_fout_int_sat[52]),
    .out_final_valid(calc_fout_int_vld[52]),
    .out_partial_data(calc_pout_int_52_sum),
    .out_partial_valid(calc_pout_int_vld[52])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8553" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_53 (
    .cfg_truncate(cfg_truncate[269:265]),
    .in_data(calc_op0_int_53_d1),
    .in_op(calc_op1_int_53_d1),
    .in_op_valid(calc_op1_vld_int_d1[53]),
    .in_sel(calc_dlv_en_int_d1[53]),
    .in_valid(calc_op_en_int_d1[53]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_53_sum),
    .out_final_sat(calc_fout_int_sat[53]),
    .out_final_valid(calc_fout_int_vld[53]),
    .out_partial_data(calc_pout_int_53_sum),
    .out_partial_valid(calc_pout_int_vld[53])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8568" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_54 (
    .cfg_truncate(cfg_truncate[274:270]),
    .in_data(calc_op0_int_54_d1),
    .in_op(calc_op1_int_54_d1),
    .in_op_valid(calc_op1_vld_int_d1[54]),
    .in_sel(calc_dlv_en_int_d1[54]),
    .in_valid(calc_op_en_int_d1[54]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_54_sum),
    .out_final_sat(calc_fout_int_sat[54]),
    .out_final_valid(calc_fout_int_vld[54]),
    .out_partial_data(calc_pout_int_54_sum),
    .out_partial_valid(calc_pout_int_vld[54])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8583" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_55 (
    .cfg_truncate(cfg_truncate[279:275]),
    .in_data(calc_op0_int_55_d1),
    .in_op(calc_op1_int_55_d1),
    .in_op_valid(calc_op1_vld_int_d1[55]),
    .in_sel(calc_dlv_en_int_d1[55]),
    .in_valid(calc_op_en_int_d1[55]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_55_sum),
    .out_final_sat(calc_fout_int_sat[55]),
    .out_final_valid(calc_fout_int_vld[55]),
    .out_partial_data(calc_pout_int_55_sum),
    .out_partial_valid(calc_pout_int_vld[55])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8598" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_56 (
    .cfg_truncate(cfg_truncate[284:280]),
    .in_data(calc_op0_int_56_d1),
    .in_op(calc_op1_int_56_d1),
    .in_op_valid(calc_op1_vld_int_d1[56]),
    .in_sel(calc_dlv_en_int_d1[56]),
    .in_valid(calc_op_en_int_d1[56]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_56_sum),
    .out_final_sat(calc_fout_int_sat[56]),
    .out_final_valid(calc_fout_int_vld[56]),
    .out_partial_data(calc_pout_int_56_sum),
    .out_partial_valid(calc_pout_int_vld[56])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8613" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_57 (
    .cfg_truncate(cfg_truncate[289:285]),
    .in_data(calc_op0_int_57_d1),
    .in_op(calc_op1_int_57_d1),
    .in_op_valid(calc_op1_vld_int_d1[57]),
    .in_sel(calc_dlv_en_int_d1[57]),
    .in_valid(calc_op_en_int_d1[57]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_57_sum),
    .out_final_sat(calc_fout_int_sat[57]),
    .out_final_valid(calc_fout_int_vld[57]),
    .out_partial_data(calc_pout_int_57_sum),
    .out_partial_valid(calc_pout_int_vld[57])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8628" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_58 (
    .cfg_truncate(cfg_truncate[294:290]),
    .in_data(calc_op0_int_58_d1),
    .in_op(calc_op1_int_58_d1),
    .in_op_valid(calc_op1_vld_int_d1[58]),
    .in_sel(calc_dlv_en_int_d1[58]),
    .in_valid(calc_op_en_int_d1[58]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_58_sum),
    .out_final_sat(calc_fout_int_sat[58]),
    .out_final_valid(calc_fout_int_vld[58]),
    .out_partial_data(calc_pout_int_58_sum),
    .out_partial_valid(calc_pout_int_vld[58])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8643" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_59 (
    .cfg_truncate(cfg_truncate[299:295]),
    .in_data(calc_op0_int_59_d1),
    .in_op(calc_op1_int_59_d1),
    .in_op_valid(calc_op1_vld_int_d1[59]),
    .in_sel(calc_dlv_en_int_d1[59]),
    .in_valid(calc_op_en_int_d1[59]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_59_sum),
    .out_final_sat(calc_fout_int_sat[59]),
    .out_final_valid(calc_fout_int_vld[59]),
    .out_partial_data(calc_pout_int_59_sum),
    .out_partial_valid(calc_pout_int_vld[59])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7848" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_6 (
    .cfg_truncate(cfg_truncate[34:30]),
    .in_data(calc_op0_int_6_d1),
    .in_op(calc_op1_int_6_d1),
    .in_op_valid(calc_op1_vld_int_d1[6]),
    .in_sel(calc_dlv_en_int_d1[6]),
    .in_valid(calc_op_en_int_d1[6]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_6_sum),
    .out_final_sat(calc_fout_int_sat[6]),
    .out_final_valid(calc_fout_int_vld[6]),
    .out_partial_data(calc_pout_int_6_sum),
    .out_partial_valid(calc_pout_int_vld[6])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8658" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_60 (
    .cfg_truncate(cfg_truncate[304:300]),
    .in_data(calc_op0_int_60_d1),
    .in_op(calc_op1_int_60_d1),
    .in_op_valid(calc_op1_vld_int_d1[60]),
    .in_sel(calc_dlv_en_int_d1[60]),
    .in_valid(calc_op_en_int_d1[60]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_60_sum),
    .out_final_sat(calc_fout_int_sat[60]),
    .out_final_valid(calc_fout_int_vld[60]),
    .out_partial_data(calc_pout_int_60_sum),
    .out_partial_valid(calc_pout_int_vld[60])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8673" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_61 (
    .cfg_truncate(cfg_truncate[309:305]),
    .in_data(calc_op0_int_61_d1),
    .in_op(calc_op1_int_61_d1),
    .in_op_valid(calc_op1_vld_int_d1[61]),
    .in_sel(calc_dlv_en_int_d1[61]),
    .in_valid(calc_op_en_int_d1[61]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_61_sum),
    .out_final_sat(calc_fout_int_sat[61]),
    .out_final_valid(calc_fout_int_vld[61]),
    .out_partial_data(calc_pout_int_61_sum),
    .out_partial_valid(calc_pout_int_vld[61])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8688" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_62 (
    .cfg_truncate(cfg_truncate[314:310]),
    .in_data(calc_op0_int_62_d1),
    .in_op(calc_op1_int_62_d1),
    .in_op_valid(calc_op1_vld_int_d1[62]),
    .in_sel(calc_dlv_en_int_d1[62]),
    .in_valid(calc_op_en_int_d1[62]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_62_sum),
    .out_final_sat(calc_fout_int_sat[62]),
    .out_final_valid(calc_fout_int_vld[62]),
    .out_partial_data(calc_pout_int_62_sum),
    .out_partial_valid(calc_pout_int_vld[62])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8703" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_63 (
    .cfg_truncate(cfg_truncate[319:315]),
    .in_data(calc_op0_int_63_d1),
    .in_op(calc_op1_int_63_d1),
    .in_op_valid(calc_op1_vld_int_d1[63]),
    .in_sel(calc_dlv_en_int_d1[63]),
    .in_valid(calc_op_en_int_d1[63]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_63_sum),
    .out_final_sat(calc_fout_int_sat[63]),
    .out_final_valid(calc_fout_int_vld[63]),
    .out_partial_data(calc_pout_int_63_sum),
    .out_partial_valid(calc_pout_int_vld[63])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8718" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_64 (
    .cfg_truncate(cfg_truncate[324:320]),
    .in_data(calc_op0_int_64_d1),
    .in_op(calc_op1_int_64_d1),
    .in_op_valid(calc_op1_vld_int_d1[64]),
    .in_sel(calc_dlv_en_int_d1[64]),
    .in_valid(calc_op_en_int_d1[64]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_64_sum),
    .out_final_sat(calc_fout_int_sat[64]),
    .out_final_valid(calc_fout_int_vld[64]),
    .out_partial_data(calc_pout_int_64_sum),
    .out_partial_valid(calc_pout_int_vld[64])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8733" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_65 (
    .cfg_truncate(cfg_truncate[329:325]),
    .in_data(calc_op0_int_65_d1),
    .in_op(calc_op1_int_65_d1),
    .in_op_valid(calc_op1_vld_int_d1[65]),
    .in_sel(calc_dlv_en_int_d1[65]),
    .in_valid(calc_op_en_int_d1[65]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_65_sum),
    .out_final_sat(calc_fout_int_sat[65]),
    .out_final_valid(calc_fout_int_vld[65]),
    .out_partial_data(calc_pout_int_65_sum),
    .out_partial_valid(calc_pout_int_vld[65])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8748" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_66 (
    .cfg_truncate(cfg_truncate[334:330]),
    .in_data(calc_op0_int_66_d1),
    .in_op(calc_op1_int_66_d1),
    .in_op_valid(calc_op1_vld_int_d1[66]),
    .in_sel(calc_dlv_en_int_d1[66]),
    .in_valid(calc_op_en_int_d1[66]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_66_sum),
    .out_final_sat(calc_fout_int_sat[66]),
    .out_final_valid(calc_fout_int_vld[66]),
    .out_partial_data(calc_pout_int_66_sum),
    .out_partial_valid(calc_pout_int_vld[66])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8763" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_67 (
    .cfg_truncate(cfg_truncate[339:335]),
    .in_data(calc_op0_int_67_d1),
    .in_op(calc_op1_int_67_d1),
    .in_op_valid(calc_op1_vld_int_d1[67]),
    .in_sel(calc_dlv_en_int_d1[67]),
    .in_valid(calc_op_en_int_d1[67]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_67_sum),
    .out_final_sat(calc_fout_int_sat[67]),
    .out_final_valid(calc_fout_int_vld[67]),
    .out_partial_data(calc_pout_int_67_sum),
    .out_partial_valid(calc_pout_int_vld[67])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8778" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_68 (
    .cfg_truncate(cfg_truncate[344:340]),
    .in_data(calc_op0_int_68_d1),
    .in_op(calc_op1_int_68_d1),
    .in_op_valid(calc_op1_vld_int_d1[68]),
    .in_sel(calc_dlv_en_int_d1[68]),
    .in_valid(calc_op_en_int_d1[68]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_68_sum),
    .out_final_sat(calc_fout_int_sat[68]),
    .out_final_valid(calc_fout_int_vld[68]),
    .out_partial_data(calc_pout_int_68_sum),
    .out_partial_valid(calc_pout_int_vld[68])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8793" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_69 (
    .cfg_truncate(cfg_truncate[349:345]),
    .in_data(calc_op0_int_69_d1),
    .in_op(calc_op1_int_69_d1),
    .in_op_valid(calc_op1_vld_int_d1[69]),
    .in_sel(calc_dlv_en_int_d1[69]),
    .in_valid(calc_op_en_int_d1[69]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_69_sum),
    .out_final_sat(calc_fout_int_sat[69]),
    .out_final_valid(calc_fout_int_vld[69]),
    .out_partial_data(calc_pout_int_69_sum),
    .out_partial_valid(calc_pout_int_vld[69])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7863" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_7 (
    .cfg_truncate(cfg_truncate[39:35]),
    .in_data(calc_op0_int_7_d1),
    .in_op(calc_op1_int_7_d1),
    .in_op_valid(calc_op1_vld_int_d1[7]),
    .in_sel(calc_dlv_en_int_d1[7]),
    .in_valid(calc_op_en_int_d1[7]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_7_sum),
    .out_final_sat(calc_fout_int_sat[7]),
    .out_final_valid(calc_fout_int_vld[7]),
    .out_partial_data(calc_pout_int_7_sum),
    .out_partial_valid(calc_pout_int_vld[7])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8808" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_70 (
    .cfg_truncate(cfg_truncate[354:350]),
    .in_data(calc_op0_int_70_d1),
    .in_op(calc_op1_int_70_d1),
    .in_op_valid(calc_op1_vld_int_d1[70]),
    .in_sel(calc_dlv_en_int_d1[70]),
    .in_valid(calc_op_en_int_d1[70]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_70_sum),
    .out_final_sat(calc_fout_int_sat[70]),
    .out_final_valid(calc_fout_int_vld[70]),
    .out_partial_data(calc_pout_int_70_sum),
    .out_partial_valid(calc_pout_int_vld[70])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8823" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_71 (
    .cfg_truncate(cfg_truncate[359:355]),
    .in_data(calc_op0_int_71_d1),
    .in_op(calc_op1_int_71_d1),
    .in_op_valid(calc_op1_vld_int_d1[71]),
    .in_sel(calc_dlv_en_int_d1[71]),
    .in_valid(calc_op_en_int_d1[71]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_71_sum),
    .out_final_sat(calc_fout_int_sat[71]),
    .out_final_valid(calc_fout_int_vld[71]),
    .out_partial_data(calc_pout_int_71_sum),
    .out_partial_valid(calc_pout_int_vld[71])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8838" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_72 (
    .cfg_truncate(cfg_truncate[364:360]),
    .in_data(calc_op0_int_72_d1),
    .in_op(calc_op1_int_72_d1),
    .in_op_valid(calc_op1_vld_int_d1[72]),
    .in_sel(calc_dlv_en_int_d1[72]),
    .in_valid(calc_op_en_int_d1[72]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_72_sum),
    .out_final_sat(calc_fout_int_sat[72]),
    .out_final_valid(calc_fout_int_vld[72]),
    .out_partial_data(calc_pout_int_72_sum),
    .out_partial_valid(calc_pout_int_vld[72])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8853" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_73 (
    .cfg_truncate(cfg_truncate[369:365]),
    .in_data(calc_op0_int_73_d1),
    .in_op(calc_op1_int_73_d1),
    .in_op_valid(calc_op1_vld_int_d1[73]),
    .in_sel(calc_dlv_en_int_d1[73]),
    .in_valid(calc_op_en_int_d1[73]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_73_sum),
    .out_final_sat(calc_fout_int_sat[73]),
    .out_final_valid(calc_fout_int_vld[73]),
    .out_partial_data(calc_pout_int_73_sum),
    .out_partial_valid(calc_pout_int_vld[73])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8868" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_74 (
    .cfg_truncate(cfg_truncate[374:370]),
    .in_data(calc_op0_int_74_d1),
    .in_op(calc_op1_int_74_d1),
    .in_op_valid(calc_op1_vld_int_d1[74]),
    .in_sel(calc_dlv_en_int_d1[74]),
    .in_valid(calc_op_en_int_d1[74]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_74_sum),
    .out_final_sat(calc_fout_int_sat[74]),
    .out_final_valid(calc_fout_int_vld[74]),
    .out_partial_data(calc_pout_int_74_sum),
    .out_partial_valid(calc_pout_int_vld[74])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8883" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_75 (
    .cfg_truncate(cfg_truncate[379:375]),
    .in_data(calc_op0_int_75_d1),
    .in_op(calc_op1_int_75_d1),
    .in_op_valid(calc_op1_vld_int_d1[75]),
    .in_sel(calc_dlv_en_int_d1[75]),
    .in_valid(calc_op_en_int_d1[75]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_75_sum),
    .out_final_sat(calc_fout_int_sat[75]),
    .out_final_valid(calc_fout_int_vld[75]),
    .out_partial_data(calc_pout_int_75_sum),
    .out_partial_valid(calc_pout_int_vld[75])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8898" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_76 (
    .cfg_truncate(cfg_truncate[384:380]),
    .in_data(calc_op0_int_76_d1),
    .in_op(calc_op1_int_76_d1),
    .in_op_valid(calc_op1_vld_int_d1[76]),
    .in_sel(calc_dlv_en_int_d1[76]),
    .in_valid(calc_op_en_int_d1[76]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_76_sum),
    .out_final_sat(calc_fout_int_sat[76]),
    .out_final_valid(calc_fout_int_vld[76]),
    .out_partial_data(calc_pout_int_76_sum),
    .out_partial_valid(calc_pout_int_vld[76])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8913" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_77 (
    .cfg_truncate(cfg_truncate[389:385]),
    .in_data(calc_op0_int_77_d1),
    .in_op(calc_op1_int_77_d1),
    .in_op_valid(calc_op1_vld_int_d1[77]),
    .in_sel(calc_dlv_en_int_d1[77]),
    .in_valid(calc_op_en_int_d1[77]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_77_sum),
    .out_final_sat(calc_fout_int_sat[77]),
    .out_final_valid(calc_fout_int_vld[77]),
    .out_partial_data(calc_pout_int_77_sum),
    .out_partial_valid(calc_pout_int_vld[77])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8928" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_78 (
    .cfg_truncate(cfg_truncate[394:390]),
    .in_data(calc_op0_int_78_d1),
    .in_op(calc_op1_int_78_d1),
    .in_op_valid(calc_op1_vld_int_d1[78]),
    .in_sel(calc_dlv_en_int_d1[78]),
    .in_valid(calc_op_en_int_d1[78]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_78_sum),
    .out_final_sat(calc_fout_int_sat[78]),
    .out_final_valid(calc_fout_int_vld[78]),
    .out_partial_data(calc_pout_int_78_sum),
    .out_partial_valid(calc_pout_int_vld[78])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8943" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_79 (
    .cfg_truncate(cfg_truncate[399:395]),
    .in_data(calc_op0_int_79_d1),
    .in_op(calc_op1_int_79_d1),
    .in_op_valid(calc_op1_vld_int_d1[79]),
    .in_sel(calc_dlv_en_int_d1[79]),
    .in_valid(calc_op_en_int_d1[79]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_79_sum),
    .out_final_sat(calc_fout_int_sat[79]),
    .out_final_valid(calc_fout_int_vld[79]),
    .out_partial_data(calc_pout_int_79_sum),
    .out_partial_valid(calc_pout_int_vld[79])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7878" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_8 (
    .cfg_truncate(cfg_truncate[44:40]),
    .in_data(calc_op0_int_8_d1),
    .in_op(calc_op1_int_8_d1),
    .in_op_valid(calc_op1_vld_int_d1[8]),
    .in_sel(calc_dlv_en_int_d1[8]),
    .in_valid(calc_op_en_int_d1[8]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_8_sum),
    .out_final_sat(calc_fout_int_sat[8]),
    .out_final_valid(calc_fout_int_vld[8]),
    .out_partial_data(calc_pout_int_8_sum),
    .out_partial_valid(calc_pout_int_vld[8])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8958" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_80 (
    .cfg_truncate(cfg_truncate[404:400]),
    .in_data(calc_op0_int_80_d1),
    .in_op(calc_op1_int_80_d1),
    .in_op_valid(calc_op1_vld_int_d1[80]),
    .in_sel(calc_dlv_en_int_d1[80]),
    .in_valid(calc_op_en_int_d1[80]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_80_sum),
    .out_final_sat(calc_fout_int_sat[80]),
    .out_final_valid(calc_fout_int_vld[80]),
    .out_partial_data(calc_pout_int_80_sum),
    .out_partial_valid(calc_pout_int_vld[80])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8973" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_81 (
    .cfg_truncate(cfg_truncate[409:405]),
    .in_data(calc_op0_int_81_d1),
    .in_op(calc_op1_int_81_d1),
    .in_op_valid(calc_op1_vld_int_d1[81]),
    .in_sel(calc_dlv_en_int_d1[81]),
    .in_valid(calc_op_en_int_d1[81]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_81_sum),
    .out_final_sat(calc_fout_int_sat[81]),
    .out_final_valid(calc_fout_int_vld[81]),
    .out_partial_data(calc_pout_int_81_sum),
    .out_partial_valid(calc_pout_int_vld[81])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:8988" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_82 (
    .cfg_truncate(cfg_truncate[414:410]),
    .in_data(calc_op0_int_82_d1),
    .in_op(calc_op1_int_82_d1),
    .in_op_valid(calc_op1_vld_int_d1[82]),
    .in_sel(calc_dlv_en_int_d1[82]),
    .in_valid(calc_op_en_int_d1[82]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_82_sum),
    .out_final_sat(calc_fout_int_sat[82]),
    .out_final_valid(calc_fout_int_vld[82]),
    .out_partial_data(calc_pout_int_82_sum),
    .out_partial_valid(calc_pout_int_vld[82])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9003" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_83 (
    .cfg_truncate(cfg_truncate[419:415]),
    .in_data(calc_op0_int_83_d1),
    .in_op(calc_op1_int_83_d1),
    .in_op_valid(calc_op1_vld_int_d1[83]),
    .in_sel(calc_dlv_en_int_d1[83]),
    .in_valid(calc_op_en_int_d1[83]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_83_sum),
    .out_final_sat(calc_fout_int_sat[83]),
    .out_final_valid(calc_fout_int_vld[83]),
    .out_partial_data(calc_pout_int_83_sum),
    .out_partial_valid(calc_pout_int_vld[83])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9018" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_84 (
    .cfg_truncate(cfg_truncate[424:420]),
    .in_data(calc_op0_int_84_d1),
    .in_op(calc_op1_int_84_d1),
    .in_op_valid(calc_op1_vld_int_d1[84]),
    .in_sel(calc_dlv_en_int_d1[84]),
    .in_valid(calc_op_en_int_d1[84]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_84_sum),
    .out_final_sat(calc_fout_int_sat[84]),
    .out_final_valid(calc_fout_int_vld[84]),
    .out_partial_data(calc_pout_int_84_sum),
    .out_partial_valid(calc_pout_int_vld[84])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9033" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_85 (
    .cfg_truncate(cfg_truncate[429:425]),
    .in_data(calc_op0_int_85_d1),
    .in_op(calc_op1_int_85_d1),
    .in_op_valid(calc_op1_vld_int_d1[85]),
    .in_sel(calc_dlv_en_int_d1[85]),
    .in_valid(calc_op_en_int_d1[85]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_85_sum),
    .out_final_sat(calc_fout_int_sat[85]),
    .out_final_valid(calc_fout_int_vld[85]),
    .out_partial_data(calc_pout_int_85_sum),
    .out_partial_valid(calc_pout_int_vld[85])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9048" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_86 (
    .cfg_truncate(cfg_truncate[434:430]),
    .in_data(calc_op0_int_86_d1),
    .in_op(calc_op1_int_86_d1),
    .in_op_valid(calc_op1_vld_int_d1[86]),
    .in_sel(calc_dlv_en_int_d1[86]),
    .in_valid(calc_op_en_int_d1[86]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_86_sum),
    .out_final_sat(calc_fout_int_sat[86]),
    .out_final_valid(calc_fout_int_vld[86]),
    .out_partial_data(calc_pout_int_86_sum),
    .out_partial_valid(calc_pout_int_vld[86])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9063" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_87 (
    .cfg_truncate(cfg_truncate[439:435]),
    .in_data(calc_op0_int_87_d1),
    .in_op(calc_op1_int_87_d1),
    .in_op_valid(calc_op1_vld_int_d1[87]),
    .in_sel(calc_dlv_en_int_d1[87]),
    .in_valid(calc_op_en_int_d1[87]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_87_sum),
    .out_final_sat(calc_fout_int_sat[87]),
    .out_final_valid(calc_fout_int_vld[87]),
    .out_partial_data(calc_pout_int_87_sum),
    .out_partial_valid(calc_pout_int_vld[87])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9078" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_88 (
    .cfg_truncate(cfg_truncate[444:440]),
    .in_data(calc_op0_int_88_d1),
    .in_op(calc_op1_int_88_d1),
    .in_op_valid(calc_op1_vld_int_d1[88]),
    .in_sel(calc_dlv_en_int_d1[88]),
    .in_valid(calc_op_en_int_d1[88]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_88_sum),
    .out_final_sat(calc_fout_int_sat[88]),
    .out_final_valid(calc_fout_int_vld[88]),
    .out_partial_data(calc_pout_int_88_sum),
    .out_partial_valid(calc_pout_int_vld[88])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9093" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_89 (
    .cfg_truncate(cfg_truncate[449:445]),
    .in_data(calc_op0_int_89_d1),
    .in_op(calc_op1_int_89_d1),
    .in_op_valid(calc_op1_vld_int_d1[89]),
    .in_sel(calc_dlv_en_int_d1[89]),
    .in_valid(calc_op_en_int_d1[89]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_89_sum),
    .out_final_sat(calc_fout_int_sat[89]),
    .out_final_valid(calc_fout_int_vld[89]),
    .out_partial_data(calc_pout_int_89_sum),
    .out_partial_valid(calc_pout_int_vld[89])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:7893" *)
  NV_NVDLA_CACC_CALC_int16 u_cell_int_9 (
    .cfg_truncate(cfg_truncate[49:45]),
    .in_data(calc_op0_int_9_d1),
    .in_op(calc_op1_int_9_d1),
    .in_op_valid(calc_op1_vld_int_d1[9]),
    .in_sel(calc_dlv_en_int_d1[9]),
    .in_valid(calc_op_en_int_d1[9]),
    .nvdla_core_clk(nvdla_cell_clk_0),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_9_sum),
    .out_final_sat(calc_fout_int_sat[9]),
    .out_final_valid(calc_fout_int_vld[9]),
    .out_partial_data(calc_pout_int_9_sum),
    .out_partial_valid(calc_pout_int_vld[9])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9108" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_90 (
    .cfg_truncate(cfg_truncate[454:450]),
    .in_data(calc_op0_int_90_d1),
    .in_op(calc_op1_int_90_d1),
    .in_op_valid(calc_op1_vld_int_d1[90]),
    .in_sel(calc_dlv_en_int_d1[90]),
    .in_valid(calc_op_en_int_d1[90]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_90_sum),
    .out_final_sat(calc_fout_int_sat[90]),
    .out_final_valid(calc_fout_int_vld[90]),
    .out_partial_data(calc_pout_int_90_sum),
    .out_partial_valid(calc_pout_int_vld[90])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9123" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_91 (
    .cfg_truncate(cfg_truncate[459:455]),
    .in_data(calc_op0_int_91_d1),
    .in_op(calc_op1_int_91_d1),
    .in_op_valid(calc_op1_vld_int_d1[91]),
    .in_sel(calc_dlv_en_int_d1[91]),
    .in_valid(calc_op_en_int_d1[91]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_91_sum),
    .out_final_sat(calc_fout_int_sat[91]),
    .out_final_valid(calc_fout_int_vld[91]),
    .out_partial_data(calc_pout_int_91_sum),
    .out_partial_valid(calc_pout_int_vld[91])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9138" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_92 (
    .cfg_truncate(cfg_truncate[464:460]),
    .in_data(calc_op0_int_92_d1),
    .in_op(calc_op1_int_92_d1),
    .in_op_valid(calc_op1_vld_int_d1[92]),
    .in_sel(calc_dlv_en_int_d1[92]),
    .in_valid(calc_op_en_int_d1[92]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_92_sum),
    .out_final_sat(calc_fout_int_sat[92]),
    .out_final_valid(calc_fout_int_vld[92]),
    .out_partial_data(calc_pout_int_92_sum),
    .out_partial_valid(calc_pout_int_vld[92])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9153" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_93 (
    .cfg_truncate(cfg_truncate[469:465]),
    .in_data(calc_op0_int_93_d1),
    .in_op(calc_op1_int_93_d1),
    .in_op_valid(calc_op1_vld_int_d1[93]),
    .in_sel(calc_dlv_en_int_d1[93]),
    .in_valid(calc_op_en_int_d1[93]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_93_sum),
    .out_final_sat(calc_fout_int_sat[93]),
    .out_final_valid(calc_fout_int_vld[93]),
    .out_partial_data(calc_pout_int_93_sum),
    .out_partial_valid(calc_pout_int_vld[93])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9168" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_94 (
    .cfg_truncate(cfg_truncate[474:470]),
    .in_data(calc_op0_int_94_d1),
    .in_op(calc_op1_int_94_d1),
    .in_op_valid(calc_op1_vld_int_d1[94]),
    .in_sel(calc_dlv_en_int_d1[94]),
    .in_valid(calc_op_en_int_d1[94]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_94_sum),
    .out_final_sat(calc_fout_int_sat[94]),
    .out_final_valid(calc_fout_int_vld[94]),
    .out_partial_data(calc_pout_int_94_sum),
    .out_partial_valid(calc_pout_int_vld[94])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9183" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_95 (
    .cfg_truncate(cfg_truncate[479:475]),
    .in_data(calc_op0_int_95_d1),
    .in_op(calc_op1_int_95_d1),
    .in_op_valid(calc_op1_vld_int_d1[95]),
    .in_sel(calc_dlv_en_int_d1[95]),
    .in_valid(calc_op_en_int_d1[95]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_95_sum),
    .out_final_sat(calc_fout_int_sat[95]),
    .out_final_valid(calc_fout_int_vld[95]),
    .out_partial_data(calc_pout_int_95_sum),
    .out_partial_valid(calc_pout_int_vld[95])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9198" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_96 (
    .cfg_truncate(cfg_truncate[484:480]),
    .in_data(calc_op0_int_96_d1),
    .in_op(calc_op1_int_96_d1),
    .in_op_valid(calc_op1_vld_int_d1[96]),
    .in_sel(calc_dlv_en_int_d1[96]),
    .in_valid(calc_op_en_int_d1[96]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_96_sum),
    .out_final_sat(calc_fout_int_sat[96]),
    .out_final_valid(calc_fout_int_vld[96]),
    .out_partial_data(calc_pout_int_96_sum),
    .out_partial_valid(calc_pout_int_vld[96])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9213" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_97 (
    .cfg_truncate(cfg_truncate[489:485]),
    .in_data(calc_op0_int_97_d1),
    .in_op(calc_op1_int_97_d1),
    .in_op_valid(calc_op1_vld_int_d1[97]),
    .in_sel(calc_dlv_en_int_d1[97]),
    .in_valid(calc_op_en_int_d1[97]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_97_sum),
    .out_final_sat(calc_fout_int_sat[97]),
    .out_final_valid(calc_fout_int_vld[97]),
    .out_partial_data(calc_pout_int_97_sum),
    .out_partial_valid(calc_pout_int_vld[97])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9228" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_98 (
    .cfg_truncate(cfg_truncate[494:490]),
    .in_data(calc_op0_int_98_d1),
    .in_op(calc_op1_int_98_d1),
    .in_op_valid(calc_op1_vld_int_d1[98]),
    .in_sel(calc_dlv_en_int_d1[98]),
    .in_valid(calc_op_en_int_d1[98]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_98_sum),
    .out_final_sat(calc_fout_int_sat[98]),
    .out_final_valid(calc_fout_int_vld[98]),
    .out_partial_data(calc_pout_int_98_sum),
    .out_partial_valid(calc_pout_int_vld[98])
  );
  (* module_not_derived = 32'd1 *)
  (* src = "./vmod/nvdla/cacc/NV_NVDLA_CACC_calculator.v:9243" *)
  NV_NVDLA_CACC_CALC_int8 u_cell_int_99 (
    .cfg_truncate(cfg_truncate[499:495]),
    .in_data(calc_op0_int_99_d1),
    .in_op(calc_op1_int_99_d1),
    .in_op_valid(calc_op1_vld_int_d1[99]),
    .in_sel(calc_dlv_en_int_d1[99]),
    .in_valid(calc_op_en_int_d1[99]),
    .nvdla_core_clk(nvdla_cell_clk_1),
    .nvdla_core_rstn(nvdla_core_rstn),
    .out_final_data(calc_fout_int_99_sum),
    .out_final_sat(calc_fout_int_sat[99]),
    .out_final_valid(calc_fout_int_vld[99]),
    .out_partial_data(calc_pout_int_99_sum),
    .out_partial_valid(calc_pout_int_vld[99])
  );
  assign abuf_in_data_0 = abuf_rd_data_0_sft[47:0];
  assign abuf_in_data_1 = abuf_rd_data_0_sft[95:48];
  assign abuf_in_data_10 = abuf_rd_data_0_sft[527:480];
  assign abuf_in_data_100 = abuf_rd_data_6[169:136];
  assign abuf_in_data_101 = abuf_rd_data_6[203:170];
  assign abuf_in_data_102 = abuf_rd_data_6[237:204];
  assign abuf_in_data_103 = abuf_rd_data_6[271:238];
  assign abuf_in_data_104 = abuf_rd_data_6[305:272];
  assign abuf_in_data_105 = abuf_rd_data_6[339:306];
  assign abuf_in_data_106 = abuf_rd_data_6[373:340];
  assign abuf_in_data_107 = abuf_rd_data_6[407:374];
  assign abuf_in_data_108 = abuf_rd_data_6[441:408];
  assign abuf_in_data_109 = abuf_rd_data_6[475:442];
  assign abuf_in_data_11 = abuf_rd_data_0_sft[575:528];
  assign abuf_in_data_110 = abuf_rd_data_6[509:476];
  assign abuf_in_data_111 = abuf_rd_data_6[543:510];
  assign abuf_in_data_112 = abuf_rd_data_7[33:0];
  assign abuf_in_data_113 = abuf_rd_data_7[67:34];
  assign abuf_in_data_114 = abuf_rd_data_7[101:68];
  assign abuf_in_data_115 = abuf_rd_data_7[135:102];
  assign abuf_in_data_116 = abuf_rd_data_7[169:136];
  assign abuf_in_data_117 = abuf_rd_data_7[203:170];
  assign abuf_in_data_118 = abuf_rd_data_7[237:204];
  assign abuf_in_data_119 = abuf_rd_data_7[271:238];
  assign abuf_in_data_12 = abuf_rd_data_0_sft[623:576];
  assign abuf_in_data_120 = abuf_rd_data_7[305:272];
  assign abuf_in_data_121 = abuf_rd_data_7[339:306];
  assign abuf_in_data_122 = abuf_rd_data_7[373:340];
  assign abuf_in_data_123 = abuf_rd_data_7[407:374];
  assign abuf_in_data_124 = abuf_rd_data_7[441:408];
  assign abuf_in_data_125 = abuf_rd_data_7[475:442];
  assign abuf_in_data_126 = abuf_rd_data_7[509:476];
  assign abuf_in_data_127 = abuf_rd_data_7[543:510];
  assign abuf_in_data_13 = abuf_rd_data_0_sft[671:624];
  assign abuf_in_data_14 = abuf_rd_data_0_sft[719:672];
  assign abuf_in_data_15 = abuf_rd_data_0_sft[767:720];
  assign abuf_in_data_16 = abuf_rd_data_1[47:0];
  assign abuf_in_data_17 = abuf_rd_data_1[95:48];
  assign abuf_in_data_18 = abuf_rd_data_1[143:96];
  assign abuf_in_data_19 = abuf_rd_data_1[191:144];
  assign abuf_in_data_2 = abuf_rd_data_0_sft[143:96];
  assign abuf_in_data_20 = abuf_rd_data_1[239:192];
  assign abuf_in_data_21 = abuf_rd_data_1[287:240];
  assign abuf_in_data_22 = abuf_rd_data_1[335:288];
  assign abuf_in_data_23 = abuf_rd_data_1[383:336];
  assign abuf_in_data_24 = abuf_rd_data_1[431:384];
  assign abuf_in_data_25 = abuf_rd_data_1[479:432];
  assign abuf_in_data_26 = abuf_rd_data_1[527:480];
  assign abuf_in_data_27 = abuf_rd_data_1[575:528];
  assign abuf_in_data_28 = abuf_rd_data_1[623:576];
  assign abuf_in_data_29 = abuf_rd_data_1[671:624];
  assign abuf_in_data_3 = abuf_rd_data_0_sft[191:144];
  assign abuf_in_data_30 = abuf_rd_data_1[719:672];
  assign abuf_in_data_31 = abuf_rd_data_1[767:720];
  assign abuf_in_data_32 = abuf_rd_data_2[47:0];
  assign abuf_in_data_33 = abuf_rd_data_2[95:48];
  assign abuf_in_data_34 = abuf_rd_data_2[143:96];
  assign abuf_in_data_35 = abuf_rd_data_2[191:144];
  assign abuf_in_data_36 = abuf_rd_data_2[239:192];
  assign abuf_in_data_37 = abuf_rd_data_2[287:240];
  assign abuf_in_data_38 = abuf_rd_data_2[335:288];
  assign abuf_in_data_39 = abuf_rd_data_2[383:336];
  assign abuf_in_data_4 = abuf_rd_data_0_sft[239:192];
  assign abuf_in_data_40 = abuf_rd_data_2[431:384];
  assign abuf_in_data_41 = abuf_rd_data_2[479:432];
  assign abuf_in_data_42 = abuf_rd_data_2[527:480];
  assign abuf_in_data_43 = abuf_rd_data_2[575:528];
  assign abuf_in_data_44 = abuf_rd_data_2[623:576];
  assign abuf_in_data_45 = abuf_rd_data_2[671:624];
  assign abuf_in_data_46 = abuf_rd_data_2[719:672];
  assign abuf_in_data_47 = abuf_rd_data_2[767:720];
  assign abuf_in_data_48 = abuf_rd_data_3[47:0];
  assign abuf_in_data_49 = abuf_rd_data_3[95:48];
  assign abuf_in_data_5 = abuf_rd_data_0_sft[287:240];
  assign abuf_in_data_50 = abuf_rd_data_3[143:96];
  assign abuf_in_data_51 = abuf_rd_data_3[191:144];
  assign abuf_in_data_52 = abuf_rd_data_3[239:192];
  assign abuf_in_data_53 = abuf_rd_data_3[287:240];
  assign abuf_in_data_54 = abuf_rd_data_3[335:288];
  assign abuf_in_data_55 = abuf_rd_data_3[383:336];
  assign abuf_in_data_56 = abuf_rd_data_3[431:384];
  assign abuf_in_data_57 = abuf_rd_data_3[479:432];
  assign abuf_in_data_58 = abuf_rd_data_3[527:480];
  assign abuf_in_data_59 = abuf_rd_data_3[575:528];
  assign abuf_in_data_6 = abuf_rd_data_0_sft[335:288];
  assign abuf_in_data_60 = abuf_rd_data_3[623:576];
  assign abuf_in_data_61 = abuf_rd_data_3[671:624];
  assign abuf_in_data_62 = abuf_rd_data_3[719:672];
  assign abuf_in_data_63 = abuf_rd_data_3[767:720];
  assign abuf_in_data_64 = abuf_rd_data_4_sft[33:0];
  assign abuf_in_data_65 = abuf_rd_data_4_sft[67:34];
  assign abuf_in_data_66 = abuf_rd_data_4_sft[101:68];
  assign abuf_in_data_67 = abuf_rd_data_4_sft[135:102];
  assign abuf_in_data_68 = abuf_rd_data_4_sft[169:136];
  assign abuf_in_data_69 = abuf_rd_data_4_sft[203:170];
  assign abuf_in_data_7 = abuf_rd_data_0_sft[383:336];
  assign abuf_in_data_70 = abuf_rd_data_4_sft[237:204];
  assign abuf_in_data_71 = abuf_rd_data_4_sft[271:238];
  assign abuf_in_data_72 = abuf_rd_data_4_sft[305:272];
  assign abuf_in_data_73 = abuf_rd_data_4_sft[339:306];
  assign abuf_in_data_74 = abuf_rd_data_4_sft[373:340];
  assign abuf_in_data_75 = abuf_rd_data_4_sft[407:374];
  assign abuf_in_data_76 = abuf_rd_data_4_sft[441:408];
  assign abuf_in_data_77 = abuf_rd_data_4_sft[475:442];
  assign abuf_in_data_78 = abuf_rd_data_4_sft[509:476];
  assign abuf_in_data_79 = abuf_rd_data_4_sft[543:510];
  assign abuf_in_data_8 = abuf_rd_data_0_sft[431:384];
  assign abuf_in_data_80 = abuf_rd_data_5[33:0];
  assign abuf_in_data_81 = abuf_rd_data_5[67:34];
  assign abuf_in_data_82 = abuf_rd_data_5[101:68];
  assign abuf_in_data_83 = abuf_rd_data_5[135:102];
  assign abuf_in_data_84 = abuf_rd_data_5[169:136];
  assign abuf_in_data_85 = abuf_rd_data_5[203:170];
  assign abuf_in_data_86 = abuf_rd_data_5[237:204];
  assign abuf_in_data_87 = abuf_rd_data_5[271:238];
  assign abuf_in_data_88 = abuf_rd_data_5[305:272];
  assign abuf_in_data_89 = abuf_rd_data_5[339:306];
  assign abuf_in_data_9 = abuf_rd_data_0_sft[479:432];
  assign abuf_in_data_90 = abuf_rd_data_5[373:340];
  assign abuf_in_data_91 = abuf_rd_data_5[407:374];
  assign abuf_in_data_92 = abuf_rd_data_5[441:408];
  assign abuf_in_data_93 = abuf_rd_data_5[475:442];
  assign abuf_in_data_94 = abuf_rd_data_5[509:476];
  assign abuf_in_data_95 = abuf_rd_data_5[543:510];
  assign abuf_in_data_96 = abuf_rd_data_6[33:0];
  assign abuf_in_data_97 = abuf_rd_data_6[67:34];
  assign abuf_in_data_98 = abuf_rd_data_6[101:68];
  assign abuf_in_data_99 = abuf_rd_data_6[135:102];
  assign abuf_rd_data_1_sft = abuf_rd_data_1;
  assign abuf_rd_data_2_sft = abuf_rd_data_2;
  assign abuf_rd_data_3_sft = abuf_rd_data_3;
  assign abuf_rd_data_5_sft = abuf_rd_data_5;
  assign abuf_rd_data_6_sft = abuf_rd_data_6;
  assign abuf_rd_data_7_sft = abuf_rd_data_7;
  assign abuf_wr_data_0_w = { calc_pout_15, calc_pout_14, calc_pout_13, calc_pout_12, calc_pout_11, calc_pout_10, calc_pout_9, calc_pout_8, calc_pout_7, calc_pout_6, calc_pout_5, calc_pout_4, calc_pout_3, calc_pout_2, calc_pout_1, calc_pout_0 };
  assign abuf_wr_data_1_w = { abuf_wr_elem_31, abuf_wr_elem_30, abuf_wr_elem_29, abuf_wr_elem_28, abuf_wr_elem_27, abuf_wr_elem_26, abuf_wr_elem_25, abuf_wr_elem_24, abuf_wr_elem_23, abuf_wr_elem_22, abuf_wr_elem_21, abuf_wr_elem_20, abuf_wr_elem_19, abuf_wr_elem_18, abuf_wr_elem_17, abuf_wr_elem_16 };
  assign abuf_wr_data_2_w = { abuf_wr_elem_47, abuf_wr_elem_46, abuf_wr_elem_45, abuf_wr_elem_44, abuf_wr_elem_43, abuf_wr_elem_42, abuf_wr_elem_41, abuf_wr_elem_40, abuf_wr_elem_39, abuf_wr_elem_38, abuf_wr_elem_37, abuf_wr_elem_36, abuf_wr_elem_35, abuf_wr_elem_34, abuf_wr_elem_33, abuf_wr_elem_32 };
  assign abuf_wr_data_3_w = { abuf_wr_elem_63, abuf_wr_elem_62, abuf_wr_elem_61, abuf_wr_elem_60, abuf_wr_elem_59, abuf_wr_elem_58, abuf_wr_elem_57, abuf_wr_elem_56, abuf_wr_elem_55, abuf_wr_elem_54, abuf_wr_elem_53, abuf_wr_elem_52, abuf_wr_elem_51, abuf_wr_elem_50, abuf_wr_elem_49, abuf_wr_elem_48 };
  assign abuf_wr_data_4_w = { calc_pout_79, calc_pout_78, calc_pout_77, calc_pout_76, calc_pout_75, calc_pout_74, calc_pout_73, calc_pout_72, calc_pout_71, calc_pout_70, calc_pout_69, calc_pout_68, calc_pout_67, calc_pout_66, calc_pout_65, calc_pout_64 };
  assign abuf_wr_data_5_w = { abuf_wr_elem_95, abuf_wr_elem_94, abuf_wr_elem_93, abuf_wr_elem_92, abuf_wr_elem_91, abuf_wr_elem_90, abuf_wr_elem_89, abuf_wr_elem_88, abuf_wr_elem_87, abuf_wr_elem_86, abuf_wr_elem_85, abuf_wr_elem_84, abuf_wr_elem_83, abuf_wr_elem_82, abuf_wr_elem_81, abuf_wr_elem_80 };
  assign abuf_wr_data_6_w = { abuf_wr_elem_111, abuf_wr_elem_110, abuf_wr_elem_109, abuf_wr_elem_108, abuf_wr_elem_107, abuf_wr_elem_106, abuf_wr_elem_105, abuf_wr_elem_104, abuf_wr_elem_103, abuf_wr_elem_102, abuf_wr_elem_101, abuf_wr_elem_100, abuf_wr_elem_99, abuf_wr_elem_98, abuf_wr_elem_97, abuf_wr_elem_96 };
  assign abuf_wr_data_7_w = { abuf_wr_elem_127, abuf_wr_elem_126, abuf_wr_elem_125, abuf_wr_elem_124, abuf_wr_elem_123, abuf_wr_elem_122, abuf_wr_elem_121, abuf_wr_elem_120, abuf_wr_elem_119, abuf_wr_elem_118, abuf_wr_elem_117, abuf_wr_elem_116, abuf_wr_elem_115, abuf_wr_elem_114, abuf_wr_elem_113, abuf_wr_elem_112 };
  assign abuf_wr_elem_0 = calc_pout_0;
  assign abuf_wr_elem_1 = calc_pout_1;
  assign abuf_wr_elem_10 = calc_pout_10;
  assign abuf_wr_elem_11 = calc_pout_11;
  assign abuf_wr_elem_12 = calc_pout_12;
  assign abuf_wr_elem_13 = calc_pout_13;
  assign abuf_wr_elem_14 = calc_pout_14;
  assign abuf_wr_elem_15 = calc_pout_15;
  assign abuf_wr_elem_2 = calc_pout_2;
  assign abuf_wr_elem_3 = calc_pout_3;
  assign abuf_wr_elem_4 = calc_pout_4;
  assign abuf_wr_elem_5 = calc_pout_5;
  assign abuf_wr_elem_6 = calc_pout_6;
  assign abuf_wr_elem_64 = calc_pout_64;
  assign abuf_wr_elem_65 = calc_pout_65;
  assign abuf_wr_elem_66 = calc_pout_66;
  assign abuf_wr_elem_67 = calc_pout_67;
  assign abuf_wr_elem_68 = calc_pout_68;
  assign abuf_wr_elem_69 = calc_pout_69;
  assign abuf_wr_elem_7 = calc_pout_7;
  assign abuf_wr_elem_70 = calc_pout_70;
  assign abuf_wr_elem_71 = calc_pout_71;
  assign abuf_wr_elem_72 = calc_pout_72;
  assign abuf_wr_elem_73 = calc_pout_73;
  assign abuf_wr_elem_74 = calc_pout_74;
  assign abuf_wr_elem_75 = calc_pout_75;
  assign abuf_wr_elem_76 = calc_pout_76;
  assign abuf_wr_elem_77 = calc_pout_77;
  assign abuf_wr_elem_78 = calc_pout_78;
  assign abuf_wr_elem_79 = calc_pout_79;
  assign abuf_wr_elem_8 = calc_pout_8;
  assign abuf_wr_elem_9 = calc_pout_9;
  assign calc_addr = accu_ctrl_pd[4:0];
  assign calc_channel_end = accu_ctrl_pd[18];
  assign calc_data_16_0 = calc_data_0[43:0];
  assign calc_data_16_1 = calc_data_0[87:44];
  assign calc_data_16_10 = calc_data_2[131:88];
  assign calc_data_16_11 = calc_data_2[175:132];
  assign calc_data_16_12 = calc_data_3[43:0];
  assign calc_data_16_13 = calc_data_3[87:44];
  assign calc_data_16_14 = calc_data_3[131:88];
  assign calc_data_16_15 = calc_data_3[175:132];
  assign calc_data_16_16 = calc_data_4[43:0];
  assign calc_data_16_17 = calc_data_4[87:44];
  assign calc_data_16_18 = calc_data_4[131:88];
  assign calc_data_16_19 = calc_data_4[175:132];
  assign calc_data_16_2 = calc_data_0[131:88];
  assign calc_data_16_20 = calc_data_5[43:0];
  assign calc_data_16_21 = calc_data_5[87:44];
  assign calc_data_16_22 = calc_data_5[131:88];
  assign calc_data_16_23 = calc_data_5[175:132];
  assign calc_data_16_24 = calc_data_6[43:0];
  assign calc_data_16_25 = calc_data_6[87:44];
  assign calc_data_16_26 = calc_data_6[131:88];
  assign calc_data_16_27 = calc_data_6[175:132];
  assign calc_data_16_28 = calc_data_7[43:0];
  assign calc_data_16_29 = calc_data_7[87:44];
  assign calc_data_16_3 = calc_data_0[175:132];
  assign calc_data_16_30 = calc_data_7[131:88];
  assign calc_data_16_31 = calc_data_7[175:132];
  assign calc_data_16_32 = calc_data_8[43:0];
  assign calc_data_16_33 = calc_data_8[87:44];
  assign calc_data_16_34 = calc_data_8[131:88];
  assign calc_data_16_35 = calc_data_8[175:132];
  assign calc_data_16_36 = calc_data_9[43:0];
  assign calc_data_16_37 = calc_data_9[87:44];
  assign calc_data_16_38 = calc_data_9[131:88];
  assign calc_data_16_39 = calc_data_9[175:132];
  assign calc_data_16_4 = calc_data_1[43:0];
  assign calc_data_16_40 = calc_data_10[43:0];
  assign calc_data_16_41 = calc_data_10[87:44];
  assign calc_data_16_42 = calc_data_10[131:88];
  assign calc_data_16_43 = calc_data_10[175:132];
  assign calc_data_16_44 = calc_data_11[43:0];
  assign calc_data_16_45 = calc_data_11[87:44];
  assign calc_data_16_46 = calc_data_11[131:88];
  assign calc_data_16_47 = calc_data_11[175:132];
  assign calc_data_16_48 = calc_data_12[43:0];
  assign calc_data_16_49 = calc_data_12[87:44];
  assign calc_data_16_5 = calc_data_1[87:44];
  assign calc_data_16_50 = calc_data_12[131:88];
  assign calc_data_16_51 = calc_data_12[175:132];
  assign calc_data_16_52 = calc_data_13[43:0];
  assign calc_data_16_53 = calc_data_13[87:44];
  assign calc_data_16_54 = calc_data_13[131:88];
  assign calc_data_16_55 = calc_data_13[175:132];
  assign calc_data_16_56 = calc_data_14[43:0];
  assign calc_data_16_57 = calc_data_14[87:44];
  assign calc_data_16_58 = calc_data_14[131:88];
  assign calc_data_16_59 = calc_data_14[175:132];
  assign calc_data_16_6 = calc_data_1[131:88];
  assign calc_data_16_60 = calc_data_15[43:0];
  assign calc_data_16_61 = calc_data_15[87:44];
  assign calc_data_16_62 = calc_data_15[131:88];
  assign calc_data_16_63 = calc_data_15[175:132];
  assign calc_data_16_7 = calc_data_1[175:132];
  assign calc_data_16_8 = calc_data_2[43:0];
  assign calc_data_16_9 = calc_data_2[87:44];
  assign calc_data_8_0 = { calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21], calc_data_0[21:0] };
  assign calc_data_8_1 = calc_data_0[43:22];
  assign calc_data_8_10 = { calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65], calc_data_1[65:44] };
  assign calc_data_8_100 = { calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109], calc_data_12[109:88] };
  assign calc_data_8_101 = calc_data_12[131:110];
  assign calc_data_8_102 = { calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153], calc_data_12[153:132] };
  assign calc_data_8_103 = calc_data_12[175:154];
  assign calc_data_8_104 = { calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21], calc_data_13[21:0] };
  assign calc_data_8_105 = calc_data_13[43:22];
  assign calc_data_8_106 = { calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65], calc_data_13[65:44] };
  assign calc_data_8_107 = calc_data_13[87:66];
  assign calc_data_8_108 = { calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109], calc_data_13[109:88] };
  assign calc_data_8_109 = calc_data_13[131:110];
  assign calc_data_8_11 = calc_data_1[87:66];
  assign calc_data_8_110 = { calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153], calc_data_13[153:132] };
  assign calc_data_8_111 = calc_data_13[175:154];
  assign calc_data_8_112 = { calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21], calc_data_14[21:0] };
  assign calc_data_8_113 = calc_data_14[43:22];
  assign calc_data_8_114 = { calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65], calc_data_14[65:44] };
  assign calc_data_8_115 = calc_data_14[87:66];
  assign calc_data_8_116 = { calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109], calc_data_14[109:88] };
  assign calc_data_8_117 = calc_data_14[131:110];
  assign calc_data_8_118 = { calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153], calc_data_14[153:132] };
  assign calc_data_8_119 = calc_data_14[175:154];
  assign calc_data_8_12 = { calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109], calc_data_1[109:88] };
  assign calc_data_8_120 = { calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21], calc_data_15[21:0] };
  assign calc_data_8_121 = calc_data_15[43:22];
  assign calc_data_8_122 = { calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65], calc_data_15[65:44] };
  assign calc_data_8_123 = calc_data_15[87:66];
  assign calc_data_8_124 = { calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109], calc_data_15[109:88] };
  assign calc_data_8_125 = calc_data_15[131:110];
  assign calc_data_8_126 = { calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153], calc_data_15[153:132] };
  assign calc_data_8_127 = calc_data_15[175:154];
  assign calc_data_8_13 = calc_data_1[131:110];
  assign calc_data_8_14 = { calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153], calc_data_1[153:132] };
  assign calc_data_8_15 = calc_data_1[175:154];
  assign calc_data_8_16 = { calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21], calc_data_2[21:0] };
  assign calc_data_8_17 = calc_data_2[43:22];
  assign calc_data_8_18 = { calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65], calc_data_2[65:44] };
  assign calc_data_8_19 = calc_data_2[87:66];
  assign calc_data_8_2 = { calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65], calc_data_0[65:44] };
  assign calc_data_8_20 = { calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109], calc_data_2[109:88] };
  assign calc_data_8_21 = calc_data_2[131:110];
  assign calc_data_8_22 = { calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153], calc_data_2[153:132] };
  assign calc_data_8_23 = calc_data_2[175:154];
  assign calc_data_8_24 = { calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21], calc_data_3[21:0] };
  assign calc_data_8_25 = calc_data_3[43:22];
  assign calc_data_8_26 = { calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65], calc_data_3[65:44] };
  assign calc_data_8_27 = calc_data_3[87:66];
  assign calc_data_8_28 = { calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109], calc_data_3[109:88] };
  assign calc_data_8_29 = calc_data_3[131:110];
  assign calc_data_8_3 = calc_data_0[87:66];
  assign calc_data_8_30 = { calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153], calc_data_3[153:132] };
  assign calc_data_8_31 = calc_data_3[175:154];
  assign calc_data_8_32 = { calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21], calc_data_4[21:0] };
  assign calc_data_8_33 = calc_data_4[43:22];
  assign calc_data_8_34 = { calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65], calc_data_4[65:44] };
  assign calc_data_8_35 = calc_data_4[87:66];
  assign calc_data_8_36 = { calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109], calc_data_4[109:88] };
  assign calc_data_8_37 = calc_data_4[131:110];
  assign calc_data_8_38 = { calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153], calc_data_4[153:132] };
  assign calc_data_8_39 = calc_data_4[175:154];
  assign calc_data_8_4 = { calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109], calc_data_0[109:88] };
  assign calc_data_8_40 = { calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21], calc_data_5[21:0] };
  assign calc_data_8_41 = calc_data_5[43:22];
  assign calc_data_8_42 = { calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65], calc_data_5[65:44] };
  assign calc_data_8_43 = calc_data_5[87:66];
  assign calc_data_8_44 = { calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109], calc_data_5[109:88] };
  assign calc_data_8_45 = calc_data_5[131:110];
  assign calc_data_8_46 = { calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153], calc_data_5[153:132] };
  assign calc_data_8_47 = calc_data_5[175:154];
  assign calc_data_8_48 = { calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21], calc_data_6[21:0] };
  assign calc_data_8_49 = calc_data_6[43:22];
  assign calc_data_8_5 = calc_data_0[131:110];
  assign calc_data_8_50 = { calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65], calc_data_6[65:44] };
  assign calc_data_8_51 = calc_data_6[87:66];
  assign calc_data_8_52 = { calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109], calc_data_6[109:88] };
  assign calc_data_8_53 = calc_data_6[131:110];
  assign calc_data_8_54 = { calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153], calc_data_6[153:132] };
  assign calc_data_8_55 = calc_data_6[175:154];
  assign calc_data_8_56 = { calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21], calc_data_7[21:0] };
  assign calc_data_8_57 = calc_data_7[43:22];
  assign calc_data_8_58 = { calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65], calc_data_7[65:44] };
  assign calc_data_8_59 = calc_data_7[87:66];
  assign calc_data_8_6 = { calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153], calc_data_0[153:132] };
  assign calc_data_8_60 = { calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109], calc_data_7[109:88] };
  assign calc_data_8_61 = calc_data_7[131:110];
  assign calc_data_8_62 = { calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153], calc_data_7[153:132] };
  assign calc_data_8_63 = calc_data_7[175:154];
  assign calc_data_8_64 = { calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21], calc_data_8[21:0] };
  assign calc_data_8_65 = calc_data_8[43:22];
  assign calc_data_8_66 = { calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65], calc_data_8[65:44] };
  assign calc_data_8_67 = calc_data_8[87:66];
  assign calc_data_8_68 = { calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109], calc_data_8[109:88] };
  assign calc_data_8_69 = calc_data_8[131:110];
  assign calc_data_8_7 = calc_data_0[175:154];
  assign calc_data_8_70 = { calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153], calc_data_8[153:132] };
  assign calc_data_8_71 = calc_data_8[175:154];
  assign calc_data_8_72 = { calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21], calc_data_9[21:0] };
  assign calc_data_8_73 = calc_data_9[43:22];
  assign calc_data_8_74 = { calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65], calc_data_9[65:44] };
  assign calc_data_8_75 = calc_data_9[87:66];
  assign calc_data_8_76 = { calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109], calc_data_9[109:88] };
  assign calc_data_8_77 = calc_data_9[131:110];
  assign calc_data_8_78 = { calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153], calc_data_9[153:132] };
  assign calc_data_8_79 = calc_data_9[175:154];
  assign calc_data_8_8 = { calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21], calc_data_1[21:0] };
  assign calc_data_8_80 = { calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21], calc_data_10[21:0] };
  assign calc_data_8_81 = calc_data_10[43:22];
  assign calc_data_8_82 = { calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65], calc_data_10[65:44] };
  assign calc_data_8_83 = calc_data_10[87:66];
  assign calc_data_8_84 = { calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109], calc_data_10[109:88] };
  assign calc_data_8_85 = calc_data_10[131:110];
  assign calc_data_8_86 = { calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153], calc_data_10[153:132] };
  assign calc_data_8_87 = calc_data_10[175:154];
  assign calc_data_8_88 = { calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21], calc_data_11[21:0] };
  assign calc_data_8_89 = calc_data_11[43:22];
  assign calc_data_8_9 = calc_data_1[43:22];
  assign calc_data_8_90 = { calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65], calc_data_11[65:44] };
  assign calc_data_8_91 = calc_data_11[87:66];
  assign calc_data_8_92 = { calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109], calc_data_11[109:88] };
  assign calc_data_8_93 = calc_data_11[131:110];
  assign calc_data_8_94 = { calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153], calc_data_11[153:132] };
  assign calc_data_8_95 = calc_data_11[175:154];
  assign calc_data_8_96 = { calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21], calc_data_12[21:0] };
  assign calc_data_8_97 = calc_data_12[43:22];
  assign calc_data_8_98 = { calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65], calc_data_12[65:44] };
  assign calc_data_8_99 = calc_data_12[87:66];
  assign calc_data_all = { calc_data_15, calc_data_14, calc_data_13, calc_data_12, calc_data_11, calc_data_10, calc_data_9, calc_data_8, calc_data_7, calc_data_6, calc_data_5, calc_data_4, calc_data_3, calc_data_2, calc_data_1, calc_data_0 };
  assign calc_dlv_elem_100 = calc_fout_50;
  assign calc_dlv_elem_102 = calc_fout_51;
  assign calc_dlv_elem_104 = calc_fout_52;
  assign calc_dlv_elem_106 = calc_fout_53;
  assign calc_dlv_elem_108 = calc_fout_54;
  assign calc_dlv_elem_110 = calc_fout_55;
  assign calc_dlv_elem_112 = calc_fout_56;
  assign calc_dlv_elem_114 = calc_fout_57;
  assign calc_dlv_elem_116 = calc_fout_58;
  assign calc_dlv_elem_118 = calc_fout_59;
  assign calc_dlv_elem_120 = calc_fout_60;
  assign calc_dlv_elem_122 = calc_fout_61;
  assign calc_dlv_elem_124 = calc_fout_62;
  assign calc_dlv_elem_126 = calc_fout_63;
  assign calc_dlv_elem_64 = calc_fout_32;
  assign calc_dlv_elem_66 = calc_fout_33;
  assign calc_dlv_elem_68 = calc_fout_34;
  assign calc_dlv_elem_70 = calc_fout_35;
  assign calc_dlv_elem_72 = calc_fout_36;
  assign calc_dlv_elem_74 = calc_fout_37;
  assign calc_dlv_elem_76 = calc_fout_38;
  assign calc_dlv_elem_78 = calc_fout_39;
  assign calc_dlv_elem_80 = calc_fout_40;
  assign calc_dlv_elem_82 = calc_fout_41;
  assign calc_dlv_elem_84 = calc_fout_42;
  assign calc_dlv_elem_86 = calc_fout_43;
  assign calc_dlv_elem_88 = calc_fout_44;
  assign calc_dlv_elem_90 = calc_fout_45;
  assign calc_dlv_elem_92 = calc_fout_46;
  assign calc_dlv_elem_94 = calc_fout_47;
  assign calc_dlv_elem_96 = calc_fout_48;
  assign calc_dlv_elem_98 = calc_fout_49;
  assign calc_dlv_elem_mask = accu_ctrl_pd[339:148];
  assign calc_dlv_en_fp = calc_dlv_elem_en[191:128];
  assign calc_dlv_en_int = calc_dlv_elem_en[127:0];
  assign calc_elem_100_w = calc_data_4[131:110];
  assign calc_elem_101_w = calc_data_5[131:110];
  assign calc_elem_102_w = calc_data_6[131:110];
  assign calc_elem_103_w = calc_data_7[131:110];
  assign calc_elem_104_w = calc_data_8[131:110];
  assign calc_elem_105_w = calc_data_9[131:110];
  assign calc_elem_106_w = calc_data_10[131:110];
  assign calc_elem_107_w = calc_data_11[131:110];
  assign calc_elem_108_w = calc_data_12[131:110];
  assign calc_elem_109_w = calc_data_13[131:110];
  assign calc_elem_110_w = calc_data_14[131:110];
  assign calc_elem_111_w = calc_data_15[131:110];
  assign calc_elem_112_w = calc_data_0[175:154];
  assign calc_elem_113_w = calc_data_1[175:154];
  assign calc_elem_114_w = calc_data_2[175:154];
  assign calc_elem_115_w = calc_data_3[175:154];
  assign calc_elem_116_w = calc_data_4[175:154];
  assign calc_elem_117_w = calc_data_5[175:154];
  assign calc_elem_118_w = calc_data_6[175:154];
  assign calc_elem_119_w = calc_data_7[175:154];
  assign calc_elem_120_w = calc_data_8[175:154];
  assign calc_elem_121_w = calc_data_9[175:154];
  assign calc_elem_122_w = calc_data_10[175:154];
  assign calc_elem_123_w = calc_data_11[175:154];
  assign calc_elem_124_w = calc_data_12[175:154];
  assign calc_elem_125_w = calc_data_13[175:154];
  assign calc_elem_126_w = calc_data_14[175:154];
  assign calc_elem_127_w = calc_data_15[175:154];
  assign calc_elem_64_w = calc_data_0[43:22];
  assign calc_elem_65_w = calc_data_1[43:22];
  assign calc_elem_66_w = calc_data_2[43:22];
  assign calc_elem_67_w = calc_data_3[43:22];
  assign calc_elem_68_w = calc_data_4[43:22];
  assign calc_elem_69_w = calc_data_5[43:22];
  assign calc_elem_70_w = calc_data_6[43:22];
  assign calc_elem_71_w = calc_data_7[43:22];
  assign calc_elem_72_w = calc_data_8[43:22];
  assign calc_elem_73_w = calc_data_9[43:22];
  assign calc_elem_74_w = calc_data_10[43:22];
  assign calc_elem_75_w = calc_data_11[43:22];
  assign calc_elem_76_w = calc_data_12[43:22];
  assign calc_elem_77_w = calc_data_13[43:22];
  assign calc_elem_78_w = calc_data_14[43:22];
  assign calc_elem_79_w = calc_data_15[43:22];
  assign calc_elem_80_w = calc_data_0[87:66];
  assign calc_elem_81_w = calc_data_1[87:66];
  assign calc_elem_82_w = calc_data_2[87:66];
  assign calc_elem_83_w = calc_data_3[87:66];
  assign calc_elem_84_w = calc_data_4[87:66];
  assign calc_elem_85_w = calc_data_5[87:66];
  assign calc_elem_86_w = calc_data_6[87:66];
  assign calc_elem_87_w = calc_data_7[87:66];
  assign calc_elem_88_w = calc_data_8[87:66];
  assign calc_elem_89_w = calc_data_9[87:66];
  assign calc_elem_90_w = calc_data_10[87:66];
  assign calc_elem_91_w = calc_data_11[87:66];
  assign calc_elem_92_w = calc_data_12[87:66];
  assign calc_elem_93_w = calc_data_13[87:66];
  assign calc_elem_94_w = calc_data_14[87:66];
  assign calc_elem_95_w = calc_data_15[87:66];
  assign calc_elem_96_w = calc_data_0[131:110];
  assign calc_elem_97_w = calc_data_1[131:110];
  assign calc_elem_98_w = calc_data_2[131:110];
  assign calc_elem_99_w = calc_data_3[131:110];
  assign calc_fout_0 = calc_dlv_elem_0;
  assign calc_fout_100 = calc_dlv_elem_73;
  assign calc_fout_101 = calc_dlv_elem_75;
  assign calc_fout_102 = calc_dlv_elem_77;
  assign calc_fout_103 = calc_dlv_elem_79;
  assign calc_fout_104 = calc_dlv_elem_81;
  assign calc_fout_105 = calc_dlv_elem_83;
  assign calc_fout_106 = calc_dlv_elem_85;
  assign calc_fout_107 = calc_dlv_elem_87;
  assign calc_fout_108 = calc_dlv_elem_89;
  assign calc_fout_109 = calc_dlv_elem_91;
  assign calc_fout_110 = calc_dlv_elem_93;
  assign calc_fout_111 = calc_dlv_elem_95;
  assign calc_fout_112 = calc_dlv_elem_97;
  assign calc_fout_113 = calc_dlv_elem_99;
  assign calc_fout_114 = calc_dlv_elem_101;
  assign calc_fout_115 = calc_dlv_elem_103;
  assign calc_fout_116 = calc_dlv_elem_105;
  assign calc_fout_117 = calc_dlv_elem_107;
  assign calc_fout_118 = calc_dlv_elem_109;
  assign calc_fout_119 = calc_dlv_elem_111;
  assign calc_fout_120 = calc_dlv_elem_113;
  assign calc_fout_121 = calc_dlv_elem_115;
  assign calc_fout_122 = calc_dlv_elem_117;
  assign calc_fout_123 = calc_dlv_elem_119;
  assign calc_fout_124 = calc_dlv_elem_121;
  assign calc_fout_125 = calc_dlv_elem_123;
  assign calc_fout_126 = calc_dlv_elem_125;
  assign calc_fout_127 = calc_dlv_elem_127;
  assign calc_fout_96 = calc_dlv_elem_65;
  assign calc_fout_97 = calc_dlv_elem_67;
  assign calc_fout_98 = calc_dlv_elem_69;
  assign calc_fout_99 = calc_dlv_elem_71;
  assign calc_layer_end = accu_ctrl_pd[19];
  assign calc_mode = accu_ctrl_pd[8:5];
  assign calc_op1_vld_fp = calc_elem_op1_vld[191:128];
  assign calc_op1_vld_int = calc_elem_op1_vld[127:0];
  assign calc_op_en_fp = calc_elem_en[191:128];
  assign calc_op_en_int = calc_elem_en[127:0];
  assign calc_pout_fp_0_sum_ext = calc_pout_fp_0_sum;
  assign calc_pout_fp_10_sum_ext = calc_pout_fp_10_sum;
  assign calc_pout_fp_11_sum_ext = calc_pout_fp_11_sum;
  assign calc_pout_fp_12_sum_ext = calc_pout_fp_12_sum;
  assign calc_pout_fp_13_sum_ext = calc_pout_fp_13_sum;
  assign calc_pout_fp_14_sum_ext = calc_pout_fp_14_sum;
  assign calc_pout_fp_15_sum_ext = calc_pout_fp_15_sum;
  assign calc_pout_fp_16_sum_ext = calc_pout_fp_16_sum;
  assign calc_pout_fp_17_sum_ext = calc_pout_fp_17_sum;
  assign calc_pout_fp_18_sum_ext = calc_pout_fp_18_sum;
  assign calc_pout_fp_19_sum_ext = calc_pout_fp_19_sum;
  assign calc_pout_fp_1_sum_ext = calc_pout_fp_1_sum;
  assign calc_pout_fp_20_sum_ext = calc_pout_fp_20_sum;
  assign calc_pout_fp_21_sum_ext = calc_pout_fp_21_sum;
  assign calc_pout_fp_22_sum_ext = calc_pout_fp_22_sum;
  assign calc_pout_fp_23_sum_ext = calc_pout_fp_23_sum;
  assign calc_pout_fp_24_sum_ext = calc_pout_fp_24_sum;
  assign calc_pout_fp_25_sum_ext = calc_pout_fp_25_sum;
  assign calc_pout_fp_26_sum_ext = calc_pout_fp_26_sum;
  assign calc_pout_fp_27_sum_ext = calc_pout_fp_27_sum;
  assign calc_pout_fp_28_sum_ext = calc_pout_fp_28_sum;
  assign calc_pout_fp_29_sum_ext = calc_pout_fp_29_sum;
  assign calc_pout_fp_2_sum_ext = calc_pout_fp_2_sum;
  assign calc_pout_fp_30_sum_ext = calc_pout_fp_30_sum;
  assign calc_pout_fp_31_sum_ext = calc_pout_fp_31_sum;
  assign calc_pout_fp_32_sum_ext = calc_pout_fp_32_sum;
  assign calc_pout_fp_33_sum_ext = calc_pout_fp_33_sum;
  assign calc_pout_fp_34_sum_ext = calc_pout_fp_34_sum;
  assign calc_pout_fp_35_sum_ext = calc_pout_fp_35_sum;
  assign calc_pout_fp_36_sum_ext = calc_pout_fp_36_sum;
  assign calc_pout_fp_37_sum_ext = calc_pout_fp_37_sum;
  assign calc_pout_fp_38_sum_ext = calc_pout_fp_38_sum;
  assign calc_pout_fp_39_sum_ext = calc_pout_fp_39_sum;
  assign calc_pout_fp_3_sum_ext = calc_pout_fp_3_sum;
  assign calc_pout_fp_40_sum_ext = calc_pout_fp_40_sum;
  assign calc_pout_fp_41_sum_ext = calc_pout_fp_41_sum;
  assign calc_pout_fp_42_sum_ext = calc_pout_fp_42_sum;
  assign calc_pout_fp_43_sum_ext = calc_pout_fp_43_sum;
  assign calc_pout_fp_44_sum_ext = calc_pout_fp_44_sum;
  assign calc_pout_fp_45_sum_ext = calc_pout_fp_45_sum;
  assign calc_pout_fp_46_sum_ext = calc_pout_fp_46_sum;
  assign calc_pout_fp_47_sum_ext = calc_pout_fp_47_sum;
  assign calc_pout_fp_48_sum_ext = calc_pout_fp_48_sum;
  assign calc_pout_fp_49_sum_ext = calc_pout_fp_49_sum;
  assign calc_pout_fp_4_sum_ext = calc_pout_fp_4_sum;
  assign calc_pout_fp_50_sum_ext = calc_pout_fp_50_sum;
  assign calc_pout_fp_51_sum_ext = calc_pout_fp_51_sum;
  assign calc_pout_fp_52_sum_ext = calc_pout_fp_52_sum;
  assign calc_pout_fp_53_sum_ext = calc_pout_fp_53_sum;
  assign calc_pout_fp_54_sum_ext = calc_pout_fp_54_sum;
  assign calc_pout_fp_55_sum_ext = calc_pout_fp_55_sum;
  assign calc_pout_fp_56_sum_ext = calc_pout_fp_56_sum;
  assign calc_pout_fp_57_sum_ext = calc_pout_fp_57_sum;
  assign calc_pout_fp_58_sum_ext = calc_pout_fp_58_sum;
  assign calc_pout_fp_59_sum_ext = calc_pout_fp_59_sum;
  assign calc_pout_fp_5_sum_ext = calc_pout_fp_5_sum;
  assign calc_pout_fp_60_sum_ext = calc_pout_fp_60_sum;
  assign calc_pout_fp_61_sum_ext = calc_pout_fp_61_sum;
  assign calc_pout_fp_62_sum_ext = calc_pout_fp_62_sum;
  assign calc_pout_fp_63_sum_ext = calc_pout_fp_63_sum;
  assign calc_pout_fp_6_sum_ext = calc_pout_fp_6_sum;
  assign calc_pout_fp_7_sum_ext = calc_pout_fp_7_sum;
  assign calc_pout_fp_8_sum_ext = calc_pout_fp_8_sum;
  assign calc_pout_fp_9_sum_ext = calc_pout_fp_9_sum;
  assign calc_ram_sel_0 = accu_ctrl_pd[35:20];
  assign calc_ram_sel_0_ext = { accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35], accu_ctrl_pd[35:34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34], accu_ctrl_pd[34:33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33], accu_ctrl_pd[33:32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32], accu_ctrl_pd[32:31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31], accu_ctrl_pd[31:30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30], accu_ctrl_pd[30:29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29], accu_ctrl_pd[29:28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28], accu_ctrl_pd[28:27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27], accu_ctrl_pd[27:26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26], accu_ctrl_pd[26:25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25], accu_ctrl_pd[25:24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24], accu_ctrl_pd[24:23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23], accu_ctrl_pd[23:22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22], accu_ctrl_pd[22:21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21], accu_ctrl_pd[21:20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20], accu_ctrl_pd[20] };
  assign calc_ram_sel_1 = accu_ctrl_pd[51:36];
  assign calc_ram_sel_1_ext = { accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51], accu_ctrl_pd[51:50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50], accu_ctrl_pd[50:49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49], accu_ctrl_pd[49:48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48], accu_ctrl_pd[48:47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47], accu_ctrl_pd[47:46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46], accu_ctrl_pd[46:45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45], accu_ctrl_pd[45:44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44], accu_ctrl_pd[44:43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43], accu_ctrl_pd[43:42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42], accu_ctrl_pd[42:41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41], accu_ctrl_pd[41:40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40], accu_ctrl_pd[40:39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39], accu_ctrl_pd[39:38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38], accu_ctrl_pd[38:37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37], accu_ctrl_pd[37:36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36], accu_ctrl_pd[36] };
  assign calc_ram_sel_2 = accu_ctrl_pd[67:52];
  assign calc_ram_sel_2_ext = { accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67], accu_ctrl_pd[67:66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66], accu_ctrl_pd[66:65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65], accu_ctrl_pd[65:64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64], accu_ctrl_pd[64:63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63], accu_ctrl_pd[63:62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62], accu_ctrl_pd[62:61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61], accu_ctrl_pd[61:60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60], accu_ctrl_pd[60:59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59], accu_ctrl_pd[59:58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58], accu_ctrl_pd[58:57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57], accu_ctrl_pd[57:56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56], accu_ctrl_pd[56:55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55], accu_ctrl_pd[55:54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54], accu_ctrl_pd[54:53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53], accu_ctrl_pd[53:52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52], accu_ctrl_pd[52] };
  assign calc_ram_sel_3 = accu_ctrl_pd[83:68];
  assign calc_ram_sel_3_ext = { accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83], accu_ctrl_pd[83:82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82], accu_ctrl_pd[82:81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81], accu_ctrl_pd[81:80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80], accu_ctrl_pd[80:79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79], accu_ctrl_pd[79:78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78], accu_ctrl_pd[78:77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77], accu_ctrl_pd[77:76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76], accu_ctrl_pd[76:75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75], accu_ctrl_pd[75:74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74], accu_ctrl_pd[74:73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73], accu_ctrl_pd[73:72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72], accu_ctrl_pd[72:71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71], accu_ctrl_pd[71:70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70], accu_ctrl_pd[70:69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69], accu_ctrl_pd[69:68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68], accu_ctrl_pd[68] };
  assign calc_ram_sel_4 = accu_ctrl_pd[99:84];
  assign calc_ram_sel_4_ext = { accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99], accu_ctrl_pd[99:98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98], accu_ctrl_pd[98:97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97], accu_ctrl_pd[97:96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96], accu_ctrl_pd[96:95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95], accu_ctrl_pd[95:94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94], accu_ctrl_pd[94:93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93], accu_ctrl_pd[93:92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92], accu_ctrl_pd[92:91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91], accu_ctrl_pd[91:90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90], accu_ctrl_pd[90:89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89], accu_ctrl_pd[89:88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88], accu_ctrl_pd[88:87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87], accu_ctrl_pd[87:86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86], accu_ctrl_pd[86:85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85], accu_ctrl_pd[85:84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84], accu_ctrl_pd[84] };
  assign calc_ram_sel_5 = accu_ctrl_pd[115:100];
  assign calc_ram_sel_5_ext = { accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115], accu_ctrl_pd[115:114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114], accu_ctrl_pd[114:113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113], accu_ctrl_pd[113:112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112], accu_ctrl_pd[112:111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111], accu_ctrl_pd[111:110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110], accu_ctrl_pd[110:109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109], accu_ctrl_pd[109:108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108], accu_ctrl_pd[108:107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107], accu_ctrl_pd[107:106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106], accu_ctrl_pd[106:105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105], accu_ctrl_pd[105:104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104], accu_ctrl_pd[104:103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103], accu_ctrl_pd[103:102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102], accu_ctrl_pd[102:101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101], accu_ctrl_pd[101:100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100], accu_ctrl_pd[100] };
  assign calc_ram_sel_6 = accu_ctrl_pd[131:116];
  assign calc_ram_sel_6_ext = { accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131], accu_ctrl_pd[131:130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130], accu_ctrl_pd[130:129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129], accu_ctrl_pd[129:128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128], accu_ctrl_pd[128:127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127], accu_ctrl_pd[127:126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126], accu_ctrl_pd[126:125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125], accu_ctrl_pd[125:124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124], accu_ctrl_pd[124:123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123], accu_ctrl_pd[123:122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122], accu_ctrl_pd[122:121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121], accu_ctrl_pd[121:120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120], accu_ctrl_pd[120:119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119], accu_ctrl_pd[119:118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118], accu_ctrl_pd[118:117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117], accu_ctrl_pd[117:116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116], accu_ctrl_pd[116] };
  assign calc_ram_sel_7 = accu_ctrl_pd[147:132];
  assign calc_ram_sel_7_ext = { accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147], accu_ctrl_pd[147:146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146], accu_ctrl_pd[146:145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145], accu_ctrl_pd[145:144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144], accu_ctrl_pd[144:143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143], accu_ctrl_pd[143:142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142], accu_ctrl_pd[142:141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141], accu_ctrl_pd[141:140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140], accu_ctrl_pd[140:139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139], accu_ctrl_pd[139:138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138], accu_ctrl_pd[138:137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137], accu_ctrl_pd[137:136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136], accu_ctrl_pd[136:135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135], accu_ctrl_pd[135:134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134], accu_ctrl_pd[134:133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133], accu_ctrl_pd[133:132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132], accu_ctrl_pd[132] };
  assign calc_rd_mask = accu_ctrl_pd[16:9];
  assign calc_stripe_end = accu_ctrl_pd[17];
  assign calc_valid_w = calc_valid_fw_3;
  assign cfg_truncate_0 = cfg_truncate[4:0];
  assign cfg_truncate_1 = cfg_truncate[9:5];
  assign cfg_truncate_10 = cfg_truncate[54:50];
  assign cfg_truncate_100 = cfg_truncate[504:500];
  assign cfg_truncate_101 = cfg_truncate[509:505];
  assign cfg_truncate_102 = cfg_truncate[514:510];
  assign cfg_truncate_103 = cfg_truncate[519:515];
  assign cfg_truncate_104 = cfg_truncate[524:520];
  assign cfg_truncate_105 = cfg_truncate[529:525];
  assign cfg_truncate_106 = cfg_truncate[534:530];
  assign cfg_truncate_107 = cfg_truncate[539:535];
  assign cfg_truncate_108 = cfg_truncate[544:540];
  assign cfg_truncate_109 = cfg_truncate[549:545];
  assign cfg_truncate_11 = cfg_truncate[59:55];
  assign cfg_truncate_110 = cfg_truncate[554:550];
  assign cfg_truncate_111 = cfg_truncate[559:555];
  assign cfg_truncate_112 = cfg_truncate[564:560];
  assign cfg_truncate_113 = cfg_truncate[569:565];
  assign cfg_truncate_114 = cfg_truncate[574:570];
  assign cfg_truncate_115 = cfg_truncate[579:575];
  assign cfg_truncate_116 = cfg_truncate[584:580];
  assign cfg_truncate_117 = cfg_truncate[589:585];
  assign cfg_truncate_118 = cfg_truncate[594:590];
  assign cfg_truncate_119 = cfg_truncate[599:595];
  assign cfg_truncate_12 = cfg_truncate[64:60];
  assign cfg_truncate_120 = cfg_truncate[604:600];
  assign cfg_truncate_121 = cfg_truncate[609:605];
  assign cfg_truncate_122 = cfg_truncate[614:610];
  assign cfg_truncate_123 = cfg_truncate[619:615];
  assign cfg_truncate_124 = cfg_truncate[624:620];
  assign cfg_truncate_125 = cfg_truncate[629:625];
  assign cfg_truncate_126 = cfg_truncate[634:630];
  assign cfg_truncate_127 = cfg_truncate[639:635];
  assign cfg_truncate_13 = cfg_truncate[69:65];
  assign cfg_truncate_14 = cfg_truncate[74:70];
  assign cfg_truncate_15 = cfg_truncate[79:75];
  assign cfg_truncate_16 = cfg_truncate[84:80];
  assign cfg_truncate_17 = cfg_truncate[89:85];
  assign cfg_truncate_18 = cfg_truncate[94:90];
  assign cfg_truncate_19 = cfg_truncate[99:95];
  assign cfg_truncate_2 = cfg_truncate[14:10];
  assign cfg_truncate_20 = cfg_truncate[104:100];
  assign cfg_truncate_21 = cfg_truncate[109:105];
  assign cfg_truncate_22 = cfg_truncate[114:110];
  assign cfg_truncate_23 = cfg_truncate[119:115];
  assign cfg_truncate_24 = cfg_truncate[124:120];
  assign cfg_truncate_25 = cfg_truncate[129:125];
  assign cfg_truncate_26 = cfg_truncate[134:130];
  assign cfg_truncate_27 = cfg_truncate[139:135];
  assign cfg_truncate_28 = cfg_truncate[144:140];
  assign cfg_truncate_29 = cfg_truncate[149:145];
  assign cfg_truncate_3 = cfg_truncate[19:15];
  assign cfg_truncate_30 = cfg_truncate[154:150];
  assign cfg_truncate_31 = cfg_truncate[159:155];
  assign cfg_truncate_32 = cfg_truncate[164:160];
  assign cfg_truncate_33 = cfg_truncate[169:165];
  assign cfg_truncate_34 = cfg_truncate[174:170];
  assign cfg_truncate_35 = cfg_truncate[179:175];
  assign cfg_truncate_36 = cfg_truncate[184:180];
  assign cfg_truncate_37 = cfg_truncate[189:185];
  assign cfg_truncate_38 = cfg_truncate[194:190];
  assign cfg_truncate_39 = cfg_truncate[199:195];
  assign cfg_truncate_4 = cfg_truncate[24:20];
  assign cfg_truncate_40 = cfg_truncate[204:200];
  assign cfg_truncate_41 = cfg_truncate[209:205];
  assign cfg_truncate_42 = cfg_truncate[214:210];
  assign cfg_truncate_43 = cfg_truncate[219:215];
  assign cfg_truncate_44 = cfg_truncate[224:220];
  assign cfg_truncate_45 = cfg_truncate[229:225];
  assign cfg_truncate_46 = cfg_truncate[234:230];
  assign cfg_truncate_47 = cfg_truncate[239:235];
  assign cfg_truncate_48 = cfg_truncate[244:240];
  assign cfg_truncate_49 = cfg_truncate[249:245];
  assign cfg_truncate_5 = cfg_truncate[29:25];
  assign cfg_truncate_50 = cfg_truncate[254:250];
  assign cfg_truncate_51 = cfg_truncate[259:255];
  assign cfg_truncate_52 = cfg_truncate[264:260];
  assign cfg_truncate_53 = cfg_truncate[269:265];
  assign cfg_truncate_54 = cfg_truncate[274:270];
  assign cfg_truncate_55 = cfg_truncate[279:275];
  assign cfg_truncate_56 = cfg_truncate[284:280];
  assign cfg_truncate_57 = cfg_truncate[289:285];
  assign cfg_truncate_58 = cfg_truncate[294:290];
  assign cfg_truncate_59 = cfg_truncate[299:295];
  assign cfg_truncate_6 = cfg_truncate[34:30];
  assign cfg_truncate_60 = cfg_truncate[304:300];
  assign cfg_truncate_61 = cfg_truncate[309:305];
  assign cfg_truncate_62 = cfg_truncate[314:310];
  assign cfg_truncate_63 = cfg_truncate[319:315];
  assign cfg_truncate_64 = cfg_truncate[324:320];
  assign cfg_truncate_65 = cfg_truncate[329:325];
  assign cfg_truncate_66 = cfg_truncate[334:330];
  assign cfg_truncate_67 = cfg_truncate[339:335];
  assign cfg_truncate_68 = cfg_truncate[344:340];
  assign cfg_truncate_69 = cfg_truncate[349:345];
  assign cfg_truncate_7 = cfg_truncate[39:35];
  assign cfg_truncate_70 = cfg_truncate[354:350];
  assign cfg_truncate_71 = cfg_truncate[359:355];
  assign cfg_truncate_72 = cfg_truncate[364:360];
  assign cfg_truncate_73 = cfg_truncate[369:365];
  assign cfg_truncate_74 = cfg_truncate[374:370];
  assign cfg_truncate_75 = cfg_truncate[379:375];
  assign cfg_truncate_76 = cfg_truncate[384:380];
  assign cfg_truncate_77 = cfg_truncate[389:385];
  assign cfg_truncate_78 = cfg_truncate[394:390];
  assign cfg_truncate_79 = cfg_truncate[399:395];
  assign cfg_truncate_8 = cfg_truncate[44:40];
  assign cfg_truncate_80 = cfg_truncate[404:400];
  assign cfg_truncate_81 = cfg_truncate[409:405];
  assign cfg_truncate_82 = cfg_truncate[414:410];
  assign cfg_truncate_83 = cfg_truncate[419:415];
  assign cfg_truncate_84 = cfg_truncate[424:420];
  assign cfg_truncate_85 = cfg_truncate[429:425];
  assign cfg_truncate_86 = cfg_truncate[434:430];
  assign cfg_truncate_87 = cfg_truncate[439:435];
  assign cfg_truncate_88 = cfg_truncate[444:440];
  assign cfg_truncate_89 = cfg_truncate[449:445];
  assign cfg_truncate_9 = cfg_truncate[49:45];
  assign cfg_truncate_90 = cfg_truncate[454:450];
  assign cfg_truncate_91 = cfg_truncate[459:455];
  assign cfg_truncate_92 = cfg_truncate[464:460];
  assign cfg_truncate_93 = cfg_truncate[469:465];
  assign cfg_truncate_94 = cfg_truncate[474:470];
  assign cfg_truncate_95 = cfg_truncate[479:475];
  assign cfg_truncate_96 = cfg_truncate[484:480];
  assign cfg_truncate_97 = cfg_truncate[489:485];
  assign cfg_truncate_98 = cfg_truncate[494:490];
  assign cfg_truncate_99 = cfg_truncate[499:495];
  assign dlv_data_0_w = { calc_dlv_elem_15, calc_dlv_elem_14, calc_dlv_elem_13, calc_dlv_elem_12, calc_dlv_elem_11, calc_dlv_elem_10, calc_dlv_elem_9, calc_dlv_elem_8, calc_dlv_elem_7, calc_dlv_elem_6, calc_dlv_elem_5, calc_dlv_elem_4, calc_dlv_elem_3, calc_dlv_elem_2, calc_dlv_elem_1, calc_dlv_elem_0 };
  assign dlv_data_1_w = { calc_dlv_elem_31, calc_dlv_elem_30, calc_dlv_elem_29, calc_dlv_elem_28, calc_dlv_elem_27, calc_dlv_elem_26, calc_dlv_elem_25, calc_dlv_elem_24, calc_dlv_elem_23, calc_dlv_elem_22, calc_dlv_elem_21, calc_dlv_elem_20, calc_dlv_elem_19, calc_dlv_elem_18, calc_dlv_elem_17, calc_dlv_elem_16 };
  assign dlv_data_2_w = { calc_dlv_elem_47, calc_dlv_elem_46, calc_dlv_elem_45, calc_dlv_elem_44, calc_dlv_elem_43, calc_dlv_elem_42, calc_dlv_elem_41, calc_dlv_elem_40, calc_dlv_elem_39, calc_dlv_elem_38, calc_dlv_elem_37, calc_dlv_elem_36, calc_dlv_elem_35, calc_dlv_elem_34, calc_dlv_elem_33, calc_dlv_elem_32 };
  assign dlv_data_3_w = { calc_dlv_elem_63, calc_dlv_elem_62, calc_dlv_elem_61, calc_dlv_elem_60, calc_dlv_elem_59, calc_dlv_elem_58, calc_dlv_elem_57, calc_dlv_elem_56, calc_dlv_elem_55, calc_dlv_elem_54, calc_dlv_elem_53, calc_dlv_elem_52, calc_dlv_elem_51, calc_dlv_elem_50, calc_dlv_elem_49, calc_dlv_elem_48 };
  assign dlv_data_4_w = { calc_dlv_elem_79, calc_fout_39, calc_dlv_elem_77, calc_fout_38, calc_dlv_elem_75, calc_fout_37, calc_dlv_elem_73, calc_fout_36, calc_dlv_elem_71, calc_fout_35, calc_dlv_elem_69, calc_fout_34, calc_dlv_elem_67, calc_fout_33, calc_dlv_elem_65, calc_fout_32 };
  assign dlv_data_5_w = { calc_dlv_elem_95, calc_fout_47, calc_dlv_elem_93, calc_fout_46, calc_dlv_elem_91, calc_fout_45, calc_dlv_elem_89, calc_fout_44, calc_dlv_elem_87, calc_fout_43, calc_dlv_elem_85, calc_fout_42, calc_dlv_elem_83, calc_fout_41, calc_dlv_elem_81, calc_fout_40 };
  assign dlv_data_6_w = { calc_dlv_elem_111, calc_fout_55, calc_dlv_elem_109, calc_fout_54, calc_dlv_elem_107, calc_fout_53, calc_dlv_elem_105, calc_fout_52, calc_dlv_elem_103, calc_fout_51, calc_dlv_elem_101, calc_fout_50, calc_dlv_elem_99, calc_fout_49, calc_dlv_elem_97, calc_fout_48 };
  assign dlv_data_7_w = { calc_dlv_elem_127, calc_fout_63, calc_dlv_elem_125, calc_fout_62, calc_dlv_elem_123, calc_fout_61, calc_dlv_elem_121, calc_fout_60, calc_dlv_elem_119, calc_fout_59, calc_dlv_elem_117, calc_fout_58, calc_dlv_elem_115, calc_fout_57, calc_dlv_elem_113, calc_fout_56 };
  assign dlv_pd = { dlv_layer_end, dlv_stripe_end };
  assign dlv_sat_bit = calc_fout_int_sat;
  assign dlv_valid = dlv_sat_vld_d1;
  assign dp2reg_sat_count = sat_count;
endmodule
