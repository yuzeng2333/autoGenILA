module one_round(clk, key, state_in, state_out);
  input [0:0] clk ;
  input [127:0] key ;
  input [127:0] state_in ;
  output [127:0] state_out ;
// moduleRegs
// regWithFunc
endmodule
