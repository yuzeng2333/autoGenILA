module MixColsModule(io_in_0_0, io_in_0_1, io_in_0_2, io_in_0_3, io_in_1_0, io_in_1_1, io_in_1_2, io_in_1_3, io_in_2_0, io_in_2_1, io_in_2_2, io_in_2_3, io_in_3_0, io_in_3_1, io_in_3_2, io_in_3_3, io_out_0_0, io_out_0_1, io_out_0_2, io_out_0_3, io_out_1_0, io_out_1_1, io_out_1_2, io_out_1_3, io_out_2_0, io_out_2_1, io_out_2_2, io_out_2_3, io_out_3_0, io_out_3_1, io_out_3_2, io_out_3_3);
  (* src = "crypto_accelerator.v:428" *)
  wire [8:0] _GEN_0;
  (* src = "crypto_accelerator.v:438" *)
  wire [8:0] _GEN_1;
  (* src = "crypto_accelerator.v:532" *)
  wire [8:0] _GEN_10;
  (* src = "crypto_accelerator.v:542" *)
  wire [8:0] _GEN_11;
  (* src = "crypto_accelerator.v:554" *)
  wire [8:0] _GEN_12;
  (* src = "crypto_accelerator.v:564" *)
  wire [8:0] _GEN_13;
  (* src = "crypto_accelerator.v:574" *)
  wire [8:0] _GEN_14;
  (* src = "crypto_accelerator.v:584" *)
  wire [8:0] _GEN_15;
  (* src = "crypto_accelerator.v:448" *)
  wire [8:0] _GEN_2;
  (* src = "crypto_accelerator.v:458" *)
  wire [8:0] _GEN_3;
  (* src = "crypto_accelerator.v:470" *)
  wire [8:0] _GEN_4;
  (* src = "crypto_accelerator.v:480" *)
  wire [8:0] _GEN_5;
  (* src = "crypto_accelerator.v:490" *)
  wire [8:0] _GEN_6;
  (* src = "crypto_accelerator.v:500" *)
  wire [8:0] _GEN_7;
  (* src = "crypto_accelerator.v:512" *)
  wire [8:0] _GEN_8;
  (* src = "crypto_accelerator.v:522" *)
  wire [8:0] _GEN_9;
  (* src = "crypto_accelerator.v:418" *)
  wire [7:0] _T;
  (* src = "crypto_accelerator.v:419" *)
  wire [7:0] _T_1;
  (* src = "crypto_accelerator.v:515" *)
  wire [7:0] _T_100;
  (* src = "crypto_accelerator.v:516" *)
  wire [7:0] _T_101;
  (* src = "crypto_accelerator.v:517" *)
  wire _T_102;
  (* src = "crypto_accelerator.v:518" *)
  wire [8:0] _T_103;
  wire [7:0] _T_104;
  wire [7:0] _T_105;
  (* src = "crypto_accelerator.v:521" *)
  wire [8:0] _T_107;
  (* src = "crypto_accelerator.v:523" *)
  wire [8:0] _T_108;
  (* src = "crypto_accelerator.v:524" *)
  wire [7:0] _T_109;
  wire [7:0] _T_11;
  (* src = "crypto_accelerator.v:525" *)
  wire [7:0] _T_110;
  (* src = "crypto_accelerator.v:526" *)
  wire [7:0] _T_111;
  (* src = "crypto_accelerator.v:527" *)
  wire _T_112;
  (* src = "crypto_accelerator.v:528" *)
  wire [8:0] _T_113;
  wire [7:0] _T_114;
  wire [7:0] _T_115;
  (* src = "crypto_accelerator.v:531" *)
  wire [8:0] _T_117;
  (* src = "crypto_accelerator.v:533" *)
  wire [8:0] _T_118;
  (* src = "crypto_accelerator.v:534" *)
  wire [7:0] _T_119;
  (* src = "crypto_accelerator.v:429" *)
  wire [8:0] _T_12;
  (* src = "crypto_accelerator.v:535" *)
  wire [7:0] _T_120;
  (* src = "crypto_accelerator.v:536" *)
  wire [7:0] _T_121;
  (* src = "crypto_accelerator.v:537" *)
  wire _T_122;
  (* src = "crypto_accelerator.v:538" *)
  wire [8:0] _T_123;
  wire [7:0] _T_124;
  wire [7:0] _T_125;
  (* src = "crypto_accelerator.v:541" *)
  wire [8:0] _T_127;
  (* src = "crypto_accelerator.v:543" *)
  wire [8:0] _T_128;
  (* src = "crypto_accelerator.v:544" *)
  wire [7:0] _T_129;
  (* src = "crypto_accelerator.v:430" *)
  wire [7:0] _T_13;
  (* src = "crypto_accelerator.v:545" *)
  wire [7:0] _T_130;
  (* src = "crypto_accelerator.v:546" *)
  wire [7:0] _T_131;
  (* src = "crypto_accelerator.v:547" *)
  wire [7:0] _T_132;
  (* src = "crypto_accelerator.v:548" *)
  wire [7:0] _T_134;
  (* src = "crypto_accelerator.v:549" *)
  wire _T_135;
  (* src = "crypto_accelerator.v:550" *)
  wire [8:0] _T_136;
  wire [7:0] _T_137;
  wire [7:0] _T_138;
  (* src = "crypto_accelerator.v:431" *)
  wire [7:0] _T_14;
  (* src = "crypto_accelerator.v:553" *)
  wire [8:0] _T_140;
  (* src = "crypto_accelerator.v:555" *)
  wire [8:0] _T_141;
  (* src = "crypto_accelerator.v:556" *)
  wire [7:0] _T_142;
  (* src = "crypto_accelerator.v:557" *)
  wire [7:0] _T_143;
  (* src = "crypto_accelerator.v:558" *)
  wire [7:0] _T_144;
  (* src = "crypto_accelerator.v:559" *)
  wire _T_145;
  (* src = "crypto_accelerator.v:560" *)
  wire [8:0] _T_146;
  wire [7:0] _T_147;
  wire [7:0] _T_148;
  (* src = "crypto_accelerator.v:432" *)
  wire [7:0] _T_15;
  (* src = "crypto_accelerator.v:563" *)
  wire [8:0] _T_150;
  (* src = "crypto_accelerator.v:565" *)
  wire [8:0] _T_151;
  (* src = "crypto_accelerator.v:566" *)
  wire [7:0] _T_152;
  (* src = "crypto_accelerator.v:567" *)
  wire [7:0] _T_153;
  (* src = "crypto_accelerator.v:568" *)
  wire [7:0] _T_154;
  (* src = "crypto_accelerator.v:569" *)
  wire _T_155;
  (* src = "crypto_accelerator.v:570" *)
  wire [8:0] _T_156;
  wire [7:0] _T_157;
  wire [7:0] _T_158;
  (* src = "crypto_accelerator.v:433" *)
  wire _T_16;
  (* src = "crypto_accelerator.v:573" *)
  wire [8:0] _T_160;
  (* src = "crypto_accelerator.v:575" *)
  wire [8:0] _T_161;
  (* src = "crypto_accelerator.v:576" *)
  wire [7:0] _T_162;
  (* src = "crypto_accelerator.v:577" *)
  wire [7:0] _T_163;
  (* src = "crypto_accelerator.v:578" *)
  wire [7:0] _T_164;
  (* src = "crypto_accelerator.v:579" *)
  wire _T_165;
  (* src = "crypto_accelerator.v:580" *)
  wire [8:0] _T_166;
  wire [7:0] _T_167;
  (* src = "crypto_accelerator.v:582" *)
  wire [8:0] _T_168;
  (* src = "crypto_accelerator.v:434" *)
  wire [8:0] _T_17;
  (* src = "crypto_accelerator.v:583" *)
  wire [8:0] _T_170;
  (* src = "crypto_accelerator.v:585" *)
  wire [8:0] _T_171;
  wire [7:0] _T_18;
  (* src = "crypto_accelerator.v:436" *)
  wire [8:0] _T_19;
  (* src = "crypto_accelerator.v:420" *)
  wire [7:0] _T_2;
  (* src = "crypto_accelerator.v:437" *)
  wire [8:0] _T_21;
  (* src = "crypto_accelerator.v:439" *)
  wire [8:0] _T_22;
  (* src = "crypto_accelerator.v:440" *)
  wire [7:0] _T_23;
  (* src = "crypto_accelerator.v:441" *)
  wire [7:0] _T_24;
  (* src = "crypto_accelerator.v:442" *)
  wire [7:0] _T_25;
  (* src = "crypto_accelerator.v:443" *)
  wire _T_26;
  (* src = "crypto_accelerator.v:444" *)
  wire [8:0] _T_27;
  wire [7:0] _T_28;
  wire [7:0] _T_29;
  (* src = "crypto_accelerator.v:421" *)
  wire [7:0] _T_3;
  (* src = "crypto_accelerator.v:447" *)
  wire [8:0] _T_31;
  (* src = "crypto_accelerator.v:449" *)
  wire [8:0] _T_32;
  (* src = "crypto_accelerator.v:450" *)
  wire [7:0] _T_33;
  (* src = "crypto_accelerator.v:451" *)
  wire [7:0] _T_34;
  (* src = "crypto_accelerator.v:452" *)
  wire [7:0] _T_35;
  (* src = "crypto_accelerator.v:453" *)
  wire _T_36;
  (* src = "crypto_accelerator.v:454" *)
  wire [8:0] _T_37;
  wire [7:0] _T_38;
  wire [7:0] _T_39;
  (* src = "crypto_accelerator.v:457" *)
  wire [8:0] _T_41;
  (* src = "crypto_accelerator.v:459" *)
  wire [8:0] _T_42;
  (* src = "crypto_accelerator.v:460" *)
  wire [7:0] _T_43;
  (* src = "crypto_accelerator.v:461" *)
  wire [7:0] _T_44;
  (* src = "crypto_accelerator.v:462" *)
  wire [7:0] _T_45;
  (* src = "crypto_accelerator.v:463" *)
  wire [7:0] _T_46;
  (* src = "crypto_accelerator.v:464" *)
  wire [7:0] _T_48;
  (* src = "crypto_accelerator.v:465" *)
  wire _T_49;
  (* src = "crypto_accelerator.v:422" *)
  wire [7:0] _T_5;
  (* src = "crypto_accelerator.v:466" *)
  wire [8:0] _T_50;
  wire [7:0] _T_51;
  wire [7:0] _T_52;
  (* src = "crypto_accelerator.v:469" *)
  wire [8:0] _T_54;
  (* src = "crypto_accelerator.v:471" *)
  wire [8:0] _T_55;
  (* src = "crypto_accelerator.v:472" *)
  wire [7:0] _T_56;
  (* src = "crypto_accelerator.v:473" *)
  wire [7:0] _T_57;
  (* src = "crypto_accelerator.v:474" *)
  wire [7:0] _T_58;
  (* src = "crypto_accelerator.v:475" *)
  wire _T_59;
  (* src = "crypto_accelerator.v:423" *)
  wire _T_6;
  (* src = "crypto_accelerator.v:476" *)
  wire [8:0] _T_60;
  wire [7:0] _T_61;
  wire [7:0] _T_62;
  (* src = "crypto_accelerator.v:479" *)
  wire [8:0] _T_64;
  (* src = "crypto_accelerator.v:481" *)
  wire [8:0] _T_65;
  (* src = "crypto_accelerator.v:482" *)
  wire [7:0] _T_66;
  (* src = "crypto_accelerator.v:483" *)
  wire [7:0] _T_67;
  (* src = "crypto_accelerator.v:484" *)
  wire [7:0] _T_68;
  (* src = "crypto_accelerator.v:485" *)
  wire _T_69;
  (* src = "crypto_accelerator.v:424" *)
  wire [8:0] _T_7;
  (* src = "crypto_accelerator.v:486" *)
  wire [8:0] _T_70;
  wire [7:0] _T_71;
  wire [7:0] _T_72;
  (* src = "crypto_accelerator.v:489" *)
  wire [8:0] _T_74;
  (* src = "crypto_accelerator.v:491" *)
  wire [8:0] _T_75;
  (* src = "crypto_accelerator.v:492" *)
  wire [7:0] _T_76;
  (* src = "crypto_accelerator.v:493" *)
  wire [7:0] _T_77;
  (* src = "crypto_accelerator.v:494" *)
  wire [7:0] _T_78;
  (* src = "crypto_accelerator.v:495" *)
  wire _T_79;
  wire [7:0] _T_8;
  (* src = "crypto_accelerator.v:496" *)
  wire [8:0] _T_80;
  wire [7:0] _T_81;
  wire [7:0] _T_82;
  (* src = "crypto_accelerator.v:499" *)
  wire [8:0] _T_84;
  (* src = "crypto_accelerator.v:501" *)
  wire [8:0] _T_85;
  (* src = "crypto_accelerator.v:502" *)
  wire [7:0] _T_86;
  (* src = "crypto_accelerator.v:503" *)
  wire [7:0] _T_87;
  (* src = "crypto_accelerator.v:504" *)
  wire [7:0] _T_88;
  (* src = "crypto_accelerator.v:505" *)
  wire [7:0] _T_89;
  (* src = "crypto_accelerator.v:426" *)
  wire [8:0] _T_9;
  (* src = "crypto_accelerator.v:506" *)
  wire [7:0] _T_91;
  (* src = "crypto_accelerator.v:507" *)
  wire _T_92;
  (* src = "crypto_accelerator.v:508" *)
  wire [8:0] _T_93;
  wire [7:0] _T_94;
  wire [7:0] _T_95;
  (* src = "crypto_accelerator.v:511" *)
  wire [8:0] _T_97;
  (* src = "crypto_accelerator.v:513" *)
  wire [8:0] _T_98;
  (* src = "crypto_accelerator.v:514" *)
  wire [7:0] _T_99;
  (* src = "crypto_accelerator.v:385" *)
  input [7:0] io_in_0_0;
  (* src = "crypto_accelerator.v:386" *)
  input [7:0] io_in_0_1;
  (* src = "crypto_accelerator.v:387" *)
  input [7:0] io_in_0_2;
  (* src = "crypto_accelerator.v:388" *)
  input [7:0] io_in_0_3;
  (* src = "crypto_accelerator.v:389" *)
  input [7:0] io_in_1_0;
  (* src = "crypto_accelerator.v:390" *)
  input [7:0] io_in_1_1;
  (* src = "crypto_accelerator.v:391" *)
  input [7:0] io_in_1_2;
  (* src = "crypto_accelerator.v:392" *)
  input [7:0] io_in_1_3;
  (* src = "crypto_accelerator.v:393" *)
  input [7:0] io_in_2_0;
  (* src = "crypto_accelerator.v:394" *)
  input [7:0] io_in_2_1;
  (* src = "crypto_accelerator.v:395" *)
  input [7:0] io_in_2_2;
  (* src = "crypto_accelerator.v:396" *)
  input [7:0] io_in_2_3;
  (* src = "crypto_accelerator.v:397" *)
  input [7:0] io_in_3_0;
  (* src = "crypto_accelerator.v:398" *)
  input [7:0] io_in_3_1;
  (* src = "crypto_accelerator.v:399" *)
  input [7:0] io_in_3_2;
  (* src = "crypto_accelerator.v:400" *)
  input [7:0] io_in_3_3;
  (* src = "crypto_accelerator.v:401" *)
  output [7:0] io_out_0_0;
  (* src = "crypto_accelerator.v:402" *)
  output [7:0] io_out_0_1;
  (* src = "crypto_accelerator.v:403" *)
  output [7:0] io_out_0_2;
  (* src = "crypto_accelerator.v:404" *)
  output [7:0] io_out_0_3;
  (* src = "crypto_accelerator.v:405" *)
  output [7:0] io_out_1_0;
  (* src = "crypto_accelerator.v:406" *)
  output [7:0] io_out_1_1;
  (* src = "crypto_accelerator.v:407" *)
  output [7:0] io_out_1_2;
  (* src = "crypto_accelerator.v:408" *)
  output [7:0] io_out_1_3;
  (* src = "crypto_accelerator.v:409" *)
  output [7:0] io_out_2_0;
  (* src = "crypto_accelerator.v:410" *)
  output [7:0] io_out_2_1;
  (* src = "crypto_accelerator.v:411" *)
  output [7:0] io_out_2_2;
  (* src = "crypto_accelerator.v:412" *)
  output [7:0] io_out_2_3;
  (* src = "crypto_accelerator.v:413" *)
  output [7:0] io_out_3_0;
  (* src = "crypto_accelerator.v:414" *)
  output [7:0] io_out_3_1;
  (* src = "crypto_accelerator.v:415" *)
  output [7:0] io_out_3_2;
  (* src = "crypto_accelerator.v:416" *)
  output [7:0] io_out_3_3;
  assign _T_5 = _T & (* src = "crypto_accelerator.v:422" *) 8'b10000000;
  assign _T_9[7:0] = _T_8 & (* src = "crypto_accelerator.v:426" *) 8'b11111111;
  assign _T_15 = _T_14 & (* src = "crypto_accelerator.v:432" *) 8'b10000000;
  assign _T_19[7:0] = _T_18 & (* src = "crypto_accelerator.v:436" *) 8'b11111111;
  assign _T_25 = _T_24 & (* src = "crypto_accelerator.v:442" *) 8'b10000000;
  assign _T_29 = _T_28 & (* src = "crypto_accelerator.v:446" *) 8'b11111111;
  assign _T_35 = _T_34 & (* src = "crypto_accelerator.v:452" *) 8'b10000000;
  assign _T_39 = _T_38 & (* src = "crypto_accelerator.v:456" *) 8'b11111111;
  assign _T_48 = _T_43 & (* src = "crypto_accelerator.v:464" *) 8'b10000000;
  assign _T_52 = _T_51 & (* src = "crypto_accelerator.v:468" *) 8'b11111111;
  assign _T_58 = _T_57 & (* src = "crypto_accelerator.v:474" *) 8'b10000000;
  assign _T_62 = _T_61 & (* src = "crypto_accelerator.v:478" *) 8'b11111111;
  assign _T_68 = _T_67 & (* src = "crypto_accelerator.v:484" *) 8'b10000000;
  assign _T_72 = _T_71 & (* src = "crypto_accelerator.v:488" *) 8'b11111111;
  assign _T_78 = _T_77 & (* src = "crypto_accelerator.v:494" *) 8'b10000000;
  assign _T_82 = _T_81 & (* src = "crypto_accelerator.v:498" *) 8'b11111111;
  assign _T_91 = _T_86 & (* src = "crypto_accelerator.v:506" *) 8'b10000000;
  assign _T_95 = _T_94 & (* src = "crypto_accelerator.v:510" *) 8'b11111111;
  assign _T_101 = _T_100 & (* src = "crypto_accelerator.v:516" *) 8'b10000000;
  assign _T_105 = _T_104 & (* src = "crypto_accelerator.v:520" *) 8'b11111111;
  assign _T_111 = _T_110 & (* src = "crypto_accelerator.v:526" *) 8'b10000000;
  assign _T_115 = _T_114 & (* src = "crypto_accelerator.v:530" *) 8'b11111111;
  assign _T_121 = _T_120 & (* src = "crypto_accelerator.v:536" *) 8'b10000000;
  assign _T_125 = _T_124 & (* src = "crypto_accelerator.v:540" *) 8'b11111111;
  assign _T_134 = _T_129 & (* src = "crypto_accelerator.v:548" *) 8'b10000000;
  assign _T_138 = _T_137 & (* src = "crypto_accelerator.v:552" *) 8'b11111111;
  assign _T_144 = _T_143 & (* src = "crypto_accelerator.v:558" *) 8'b10000000;
  assign _T_148 = _T_147 & (* src = "crypto_accelerator.v:562" *) 8'b11111111;
  assign _T_154 = _T_153 & (* src = "crypto_accelerator.v:568" *) 8'b10000000;
  assign _T_158 = _T_157 & (* src = "crypto_accelerator.v:572" *) 8'b11111111;
  assign _T_164 = _T_163 & (* src = "crypto_accelerator.v:578" *) 8'b10000000;
  assign _T_168[7:0] = _T_167 & (* src = "crypto_accelerator.v:582" *) 8'b11111111;
  assign _T_6 = | (* src = "crypto_accelerator.v:423" *) _T_5;
  assign _T_16 = | (* src = "crypto_accelerator.v:433" *) _T_15;
  assign _T_26 = | (* src = "crypto_accelerator.v:443" *) _T_25;
  assign _T_36 = | (* src = "crypto_accelerator.v:453" *) _T_35;
  assign _T_49 = | (* src = "crypto_accelerator.v:465" *) _T_48;
  assign _T_59 = | (* src = "crypto_accelerator.v:475" *) _T_58;
  assign _T_69 = | (* src = "crypto_accelerator.v:485" *) _T_68;
  assign _T_79 = | (* src = "crypto_accelerator.v:495" *) _T_78;
  assign _T_92 = | (* src = "crypto_accelerator.v:507" *) _T_91;
  assign _T_102 = | (* src = "crypto_accelerator.v:517" *) _T_101;
  assign _T_112 = | (* src = "crypto_accelerator.v:527" *) _T_111;
  assign _T_122 = | (* src = "crypto_accelerator.v:537" *) _T_121;
  assign _T_135 = | (* src = "crypto_accelerator.v:549" *) _T_134;
  assign _T_145 = | (* src = "crypto_accelerator.v:559" *) _T_144;
  assign _T_155 = | (* src = "crypto_accelerator.v:569" *) _T_154;
  assign _T_165 = | (* src = "crypto_accelerator.v:579" *) _T_164;
  assign _T_11 = _T_6 ? (* src = "crypto_accelerator.v:427" *) _T_9[7:0] : { _T[6:0], 1'b0 };
  assign _T_21[7:0] = _T_16 ? (* src = "crypto_accelerator.v:437" *) _T_19[7:0] : { _T_14[6:0], 1'b0 };
  assign _T_31[7:0] = _T_26 ? (* src = "crypto_accelerator.v:447" *) _T_29 : { _T_24[6:0], 1'b0 };
  assign _T_41[7:0] = _T_36 ? (* src = "crypto_accelerator.v:457" *) _T_39 : { _T_34[6:0], 1'b0 };
  assign _T_54[7:0] = _T_49 ? (* src = "crypto_accelerator.v:469" *) _T_52 : { _T_43[6:0], 1'b0 };
  assign _T_64[7:0] = _T_59 ? (* src = "crypto_accelerator.v:479" *) _T_62 : { _T_57[6:0], 1'b0 };
  assign _T_74[7:0] = _T_69 ? (* src = "crypto_accelerator.v:489" *) _T_72 : { _T_67[6:0], 1'b0 };
  assign _T_84[7:0] = _T_79 ? (* src = "crypto_accelerator.v:499" *) _T_82 : { _T_77[6:0], 1'b0 };
  assign _T_97[7:0] = _T_92 ? (* src = "crypto_accelerator.v:511" *) _T_95 : { _T_86[6:0], 1'b0 };
  assign _T_107[7:0] = _T_102 ? (* src = "crypto_accelerator.v:521" *) _T_105 : { _T_100[6:0], 1'b0 };
  assign _T_117[7:0] = _T_112 ? (* src = "crypto_accelerator.v:531" *) _T_115 : { _T_110[6:0], 1'b0 };
  assign _T_127[7:0] = _T_122 ? (* src = "crypto_accelerator.v:541" *) _T_125 : { _T_120[6:0], 1'b0 };
  assign _T_140[7:0] = _T_135 ? (* src = "crypto_accelerator.v:553" *) _T_138 : { _T_129[6:0], 1'b0 };
  assign _T_150[7:0] = _T_145 ? (* src = "crypto_accelerator.v:563" *) _T_148 : { _T_143[6:0], 1'b0 };
  assign _T_160[7:0] = _T_155 ? (* src = "crypto_accelerator.v:573" *) _T_158 : { _T_153[6:0], 1'b0 };
  assign _T_170[7:0] = _T_165 ? (* src = "crypto_accelerator.v:583" *) _T_168[7:0] : { _T_163[6:0], 1'b0 };
  assign _T = io_in_0_0 ^ (* src = "crypto_accelerator.v:418" *) io_in_0_1;
  assign _T_1 = _T ^ (* src = "crypto_accelerator.v:419" *) io_in_0_2;
  assign _T_2 = _T_1 ^ (* src = "crypto_accelerator.v:420" *) io_in_0_3;
  assign _T_3 = io_in_0_0 ^ (* src = "crypto_accelerator.v:421" *) _T_2;
  assign _T_8 = { _T[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:425" *) 5'b11011;
  assign io_out_0_0 = _T_3 ^ (* src = "crypto_accelerator.v:429" *) _T_11;
  assign _T_13 = io_in_0_1 ^ (* src = "crypto_accelerator.v:430" *) _T_2;
  assign _T_14 = io_in_0_1 ^ (* src = "crypto_accelerator.v:431" *) io_in_0_2;
  assign _T_18 = { _T_14[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:435" *) 5'b11011;
  assign io_out_0_1 = _T_13 ^ (* src = "crypto_accelerator.v:439" *) _T_21[7:0];
  assign _T_23 = io_in_0_2 ^ (* src = "crypto_accelerator.v:440" *) _T_2;
  assign _T_24 = io_in_0_2 ^ (* src = "crypto_accelerator.v:441" *) io_in_0_3;
  assign _T_28 = { _T_24[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:445" *) 5'b11011;
  assign io_out_0_2 = _T_23 ^ (* src = "crypto_accelerator.v:449" *) _T_31[7:0];
  assign _T_33 = io_in_0_3 ^ (* src = "crypto_accelerator.v:450" *) _T_2;
  assign _T_34 = io_in_0_3 ^ (* src = "crypto_accelerator.v:451" *) io_in_0_0;
  assign _T_38 = { _T_34[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:455" *) 5'b11011;
  assign io_out_0_3 = _T_33 ^ (* src = "crypto_accelerator.v:459" *) _T_41[7:0];
  assign _T_43 = io_in_1_0 ^ (* src = "crypto_accelerator.v:460" *) io_in_1_1;
  assign _T_44 = _T_43 ^ (* src = "crypto_accelerator.v:461" *) io_in_1_2;
  assign _T_45 = _T_44 ^ (* src = "crypto_accelerator.v:462" *) io_in_1_3;
  assign _T_46 = io_in_1_0 ^ (* src = "crypto_accelerator.v:463" *) _T_45;
  assign _T_51 = { _T_43[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:467" *) 5'b11011;
  assign io_out_1_0 = _T_46 ^ (* src = "crypto_accelerator.v:471" *) _T_54[7:0];
  assign _T_56 = io_in_1_1 ^ (* src = "crypto_accelerator.v:472" *) _T_45;
  assign _T_57 = io_in_1_1 ^ (* src = "crypto_accelerator.v:473" *) io_in_1_2;
  assign _T_61 = { _T_57[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:477" *) 5'b11011;
  assign io_out_1_1 = _T_56 ^ (* src = "crypto_accelerator.v:481" *) _T_64[7:0];
  assign _T_66 = io_in_1_2 ^ (* src = "crypto_accelerator.v:482" *) _T_45;
  assign _T_67 = io_in_1_2 ^ (* src = "crypto_accelerator.v:483" *) io_in_1_3;
  assign _T_71 = { _T_67[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:487" *) 5'b11011;
  assign io_out_1_2 = _T_66 ^ (* src = "crypto_accelerator.v:491" *) _T_74[7:0];
  assign _T_76 = io_in_1_3 ^ (* src = "crypto_accelerator.v:492" *) _T_45;
  assign _T_77 = io_in_1_3 ^ (* src = "crypto_accelerator.v:493" *) io_in_1_0;
  assign _T_81 = { _T_77[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:497" *) 5'b11011;
  assign io_out_1_3 = _T_76 ^ (* src = "crypto_accelerator.v:501" *) _T_84[7:0];
  assign _T_86 = io_in_2_0 ^ (* src = "crypto_accelerator.v:502" *) io_in_2_1;
  assign _T_87 = _T_86 ^ (* src = "crypto_accelerator.v:503" *) io_in_2_2;
  assign _T_88 = _T_87 ^ (* src = "crypto_accelerator.v:504" *) io_in_2_3;
  assign _T_89 = io_in_2_0 ^ (* src = "crypto_accelerator.v:505" *) _T_88;
  assign _T_94 = { _T_86[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:509" *) 5'b11011;
  assign io_out_2_0 = _T_89 ^ (* src = "crypto_accelerator.v:513" *) _T_97[7:0];
  assign _T_99 = io_in_2_1 ^ (* src = "crypto_accelerator.v:514" *) _T_88;
  assign _T_100 = io_in_2_1 ^ (* src = "crypto_accelerator.v:515" *) io_in_2_2;
  assign _T_104 = { _T_100[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:519" *) 5'b11011;
  assign io_out_2_1 = _T_99 ^ (* src = "crypto_accelerator.v:523" *) _T_107[7:0];
  assign _T_109 = io_in_2_2 ^ (* src = "crypto_accelerator.v:524" *) _T_88;
  assign _T_110 = io_in_2_2 ^ (* src = "crypto_accelerator.v:525" *) io_in_2_3;
  assign _T_114 = { _T_110[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:529" *) 5'b11011;
  assign io_out_2_2 = _T_109 ^ (* src = "crypto_accelerator.v:533" *) _T_117[7:0];
  assign _T_119 = io_in_2_3 ^ (* src = "crypto_accelerator.v:534" *) _T_88;
  assign _T_120 = io_in_2_3 ^ (* src = "crypto_accelerator.v:535" *) io_in_2_0;
  assign _T_124 = { _T_120[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:539" *) 5'b11011;
  assign io_out_2_3 = _T_119 ^ (* src = "crypto_accelerator.v:543" *) _T_127[7:0];
  assign _T_129 = io_in_3_0 ^ (* src = "crypto_accelerator.v:544" *) io_in_3_1;
  assign _T_130 = _T_129 ^ (* src = "crypto_accelerator.v:545" *) io_in_3_2;
  assign _T_131 = _T_130 ^ (* src = "crypto_accelerator.v:546" *) io_in_3_3;
  assign _T_132 = io_in_3_0 ^ (* src = "crypto_accelerator.v:547" *) _T_131;
  assign _T_137 = { _T_129[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:551" *) 5'b11011;
  assign io_out_3_0 = _T_132 ^ (* src = "crypto_accelerator.v:555" *) _T_140[7:0];
  assign _T_142 = io_in_3_1 ^ (* src = "crypto_accelerator.v:556" *) _T_131;
  assign _T_143 = io_in_3_1 ^ (* src = "crypto_accelerator.v:557" *) io_in_3_2;
  assign _T_147 = { _T_143[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:561" *) 5'b11011;
  assign io_out_3_1 = _T_142 ^ (* src = "crypto_accelerator.v:565" *) _T_150[7:0];
  assign _T_152 = io_in_3_2 ^ (* src = "crypto_accelerator.v:566" *) _T_131;
  assign _T_153 = io_in_3_2 ^ (* src = "crypto_accelerator.v:567" *) io_in_3_3;
  assign _T_157 = { _T_153[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:571" *) 5'b11011;
  assign io_out_3_2 = _T_152 ^ (* src = "crypto_accelerator.v:575" *) _T_160[7:0];
  assign _T_162 = io_in_3_3 ^ (* src = "crypto_accelerator.v:576" *) _T_131;
  assign _T_163 = io_in_3_3 ^ (* src = "crypto_accelerator.v:577" *) io_in_3_0;
  assign _T_167 = { _T_163[6:0], 1'b0 } ^ (* src = "crypto_accelerator.v:581" *) 5'b11011;
  assign io_out_3_3 = _T_162 ^ (* src = "crypto_accelerator.v:585" *) _T_170[7:0];
  assign _GEN_0 = { 1'b0, _T_3 };
  assign _GEN_1 = { 1'b0, _T_13 };
  assign _GEN_10 = { 1'b0, _T_109 };
  assign _GEN_11 = { 1'b0, _T_119 };
  assign _GEN_12 = { 1'b0, _T_132 };
  assign _GEN_13 = { 1'b0, _T_142 };
  assign _GEN_14 = { 1'b0, _T_152 };
  assign _GEN_15 = { 1'b0, _T_162 };
  assign _GEN_2 = { 1'b0, _T_23 };
  assign _GEN_3 = { 1'b0, _T_33 };
  assign _GEN_4 = { 1'b0, _T_46 };
  assign _GEN_5 = { 1'b0, _T_56 };
  assign _GEN_6 = { 1'b0, _T_66 };
  assign _GEN_7 = { 1'b0, _T_76 };
  assign _GEN_8 = { 1'b0, _T_89 };
  assign _GEN_9 = { 1'b0, _T_99 };
  assign _T_103 = { _T_100, 1'b0 };
  assign _T_107[8] = 1'bx;
  assign _T_108[7:0] = io_out_2_1;
  assign _T_113 = { _T_110, 1'b0 };
  assign _T_117[8] = 1'bx;
  assign _T_118[7:0] = io_out_2_2;
  assign _T_12[7:0] = io_out_0_0;
  assign _T_123 = { _T_120, 1'b0 };
  assign _T_127[8] = 1'bx;
  assign _T_128[7:0] = io_out_2_3;
  assign _T_136 = { _T_129, 1'b0 };
  assign _T_140[8] = 1'bx;
  assign _T_141[7:0] = io_out_3_0;
  assign _T_146 = { _T_143, 1'b0 };
  assign _T_150[8] = 1'bx;
  assign _T_151[7:0] = io_out_3_1;
  assign _T_156 = { _T_153, 1'b0 };
  assign _T_160[8] = 1'bx;
  assign _T_161[7:0] = io_out_3_2;
  assign _T_166 = { _T_163, 1'b0 };
  assign _T_17 = { _T_14, 1'b0 };
  assign _T_170[8] = 1'bx;
  assign _T_171[7:0] = io_out_3_3;
  assign _T_21[8] = 1'bx;
  assign _T_22[7:0] = io_out_0_1;
  assign _T_27 = { _T_24, 1'b0 };
  assign _T_31[8] = 1'bx;
  assign _T_32[7:0] = io_out_0_2;
  assign _T_37 = { _T_34, 1'b0 };
  assign _T_41[8] = 1'bx;
  assign _T_42[7:0] = io_out_0_3;
  assign _T_50 = { _T_43, 1'b0 };
  assign _T_54[8] = 1'bx;
  assign _T_55[7:0] = io_out_1_0;
  assign _T_60 = { _T_57, 1'b0 };
  assign _T_64[8] = 1'bx;
  assign _T_65[7:0] = io_out_1_1;
  assign _T_7 = { _T, 1'b0 };
  assign _T_70 = { _T_67, 1'b0 };
  assign _T_74[8] = 1'bx;
  assign _T_75[7:0] = io_out_1_2;
  assign _T_80 = { _T_77, 1'b0 };
  assign _T_84[8] = 1'bx;
  assign _T_85[7:0] = io_out_1_3;
  assign _T_93 = { _T_86, 1'b0 };
  assign _T_97[8] = 1'bx;
  assign _T_98[7:0] = io_out_2_0;
endmodule
