module FP17_ADD_chn_a_rsci_unreg(in_0, outsig);
  (* src = "./vmod/vlibs/HLS_fp17_add.v:299" *)
  input in_0;
  (* src = "./vmod/vlibs/HLS_fp17_add.v:300" *)
  output outsig;
  assign outsig = in_0;
endmodule
